//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n591, new_n592, new_n593, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n633, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n464), .A2(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(KEYINPUT67), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n462), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n465), .A2(new_n466), .B1(G137), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT66), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n468), .A2(new_n475), .A3(new_n469), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(new_n476), .A3(G125), .ZN(new_n477));
  INV_X1    g052(.A(G113), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(new_n462), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  XNOR2_X1  g057(.A(new_n470), .B(KEYINPUT68), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n462), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n487), .A2(new_n489), .B1(new_n491), .B2(G124), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n473), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g074(.A(new_n499), .B(KEYINPUT70), .Z(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n470), .B2(G138), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n501), .A2(new_n496), .A3(G138), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n474), .A2(new_n476), .A3(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n474), .A2(new_n476), .A3(KEYINPUT71), .A4(new_n503), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n500), .A2(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT73), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT72), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n515), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G88), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n511), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G50), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n526), .A2(new_n528), .A3(KEYINPUT74), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT74), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n518), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(G166));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n521), .A2(new_n522), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(new_n515), .ZN(new_n539));
  INV_X1    g114(.A(G89), .ZN(new_n540));
  OAI221_X1 g115(.A(new_n536), .B1(new_n524), .B2(new_n537), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G51), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n527), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT75), .B1(new_n523), .B2(new_n511), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n541), .A2(new_n546), .ZN(G168));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n544), .B2(new_n545), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n539), .A2(new_n550), .B1(new_n517), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(G171));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n544), .B2(new_n545), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n524), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n525), .A2(G81), .B1(G651), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(new_n563));
  XOR2_X1   g138(.A(new_n563), .B(KEYINPUT76), .Z(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n511), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n521), .A2(new_n569), .A3(new_n522), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT77), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NOR3_X1   g150(.A1(new_n523), .A2(new_n570), .A3(new_n511), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n574), .B1(new_n578), .B2(new_n573), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n517), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(KEYINPUT80), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(KEYINPUT80), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n521), .A2(G91), .A3(new_n515), .A4(new_n522), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT79), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(KEYINPUT79), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n582), .A2(new_n583), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n579), .A2(new_n587), .ZN(G299));
  INV_X1    g163(.A(G171), .ZN(G301));
  INV_X1    g164(.A(G168), .ZN(G286));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n531), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g167(.A(KEYINPUT81), .B(new_n518), .C1(new_n529), .C2(new_n530), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n592), .A2(new_n593), .ZN(G303));
  NAND2_X1  g169(.A1(new_n527), .A2(G49), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n525), .A2(G87), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G288));
  AOI22_X1  g173(.A1(G48), .A2(new_n527), .B1(new_n525), .B2(G86), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n515), .A2(KEYINPUT82), .A3(G61), .ZN(new_n600));
  INV_X1    g175(.A(G73), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n601), .A2(new_n511), .A3(KEYINPUT83), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT83), .B1(new_n601), .B2(new_n511), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT82), .B1(new_n515), .B2(G61), .ZN(new_n605));
  OAI21_X1  g180(.A(G651), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n599), .A2(new_n606), .ZN(G305));
  NAND2_X1  g182(.A1(new_n544), .A2(new_n545), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n608), .A2(G47), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n539), .A2(new_n610), .B1(new_n517), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(new_n608), .A2(G54), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n539), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT84), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n517), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(new_n621), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n615), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n626), .B2(G171), .ZN(G284));
  OAI21_X1  g203(.A(new_n627), .B1(new_n626), .B2(G171), .ZN(G321));
  NAND2_X1  g204(.A1(G299), .A2(new_n626), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n626), .B2(G168), .ZN(G297));
  OAI21_X1  g206(.A(new_n630), .B1(new_n626), .B2(G168), .ZN(G280));
  INV_X1    g207(.A(new_n625), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT85), .B(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(G860), .B2(new_n634), .ZN(G148));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g214(.A1(new_n474), .A2(new_n476), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(new_n463), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT13), .B(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n496), .A2(G111), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(KEYINPUT87), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n646), .B2(KEYINPUT87), .ZN(new_n649));
  AOI22_X1  g224(.A1(new_n647), .A2(new_n649), .B1(new_n491), .B2(G123), .ZN(new_n650));
  INV_X1    g225(.A(G135), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n650), .B1(new_n483), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT88), .B(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n645), .A2(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(G2427), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT90), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT89), .B(G2438), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n657), .B(new_n658), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(new_n661), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n665), .A3(KEYINPUT14), .ZN(new_n666));
  XOR2_X1   g241(.A(G2443), .B(G2446), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2451), .B(G2454), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT91), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1341), .B(G1348), .Z(new_n673));
  OAI21_X1  g248(.A(G14), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT92), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT92), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n672), .A2(new_n677), .A3(new_n673), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n674), .B1(new_n676), .B2(new_n678), .ZN(G401));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT93), .B(KEYINPUT17), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2067), .B(G2678), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2084), .B(G2090), .Z(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT94), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n685), .B1(new_n684), .B2(new_n680), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n682), .B2(new_n684), .ZN(new_n689));
  INV_X1    g264(.A(new_n680), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n690), .A2(new_n683), .A3(new_n685), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT18), .Z(new_n692));
  NAND3_X1  g267(.A1(new_n687), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G2096), .B(G2100), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G227));
  XNOR2_X1  g270(.A(G1971), .B(G1976), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT19), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1956), .B(G2474), .Z(new_n699));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT20), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n699), .A2(new_n700), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n698), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n698), .B2(new_n704), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT95), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(G1991), .B(G1996), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT96), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1981), .B(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(G229));
  NAND3_X1  g290(.A1(new_n496), .A2(G103), .A3(G2104), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT25), .Z(new_n717));
  INV_X1    g292(.A(G139), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n483), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n640), .A2(G127), .ZN(new_n720));
  NAND2_X1  g295(.A1(G115), .A2(G2104), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n496), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT99), .Z(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n725), .B2(G33), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT100), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(G2072), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(G2072), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT30), .B(G28), .ZN(new_n731));
  OR2_X1    g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  NAND2_X1  g307(.A1(KEYINPUT31), .A2(G11), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n731), .A2(new_n725), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n652), .B2(new_n725), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n484), .A2(G141), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n463), .A2(G105), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT26), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n737), .B(new_n739), .C1(new_n491), .C2(G129), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(new_n725), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n725), .B2(G32), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n735), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G34), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(KEYINPUT24), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(KEYINPUT24), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n725), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G160), .B2(new_n725), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n746), .B(new_n753), .C1(new_n744), .C2(new_n745), .ZN(new_n754));
  INV_X1    g329(.A(G16), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G21), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G168), .B2(new_n755), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT101), .B(G1966), .Z(new_n758));
  XOR2_X1   g333(.A(new_n757), .B(new_n758), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n725), .A2(G27), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G164), .B2(new_n725), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2078), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n755), .A2(G5), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G171), .B2(new_n755), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1961), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n754), .A2(new_n759), .A3(new_n762), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n729), .A2(new_n730), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT102), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G19), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n562), .B2(G16), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(G1341), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(G1341), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n725), .A2(G35), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G162), .B2(new_n725), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT29), .B(G2090), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n725), .A2(G26), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT28), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n491), .A2(G128), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n496), .A2(G116), .ZN(new_n782));
  OAI21_X1  g357(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n783));
  INV_X1    g358(.A(G140), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n781), .B1(new_n782), .B2(new_n783), .C1(new_n483), .C2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n780), .B1(new_n785), .B2(G29), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2067), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n773), .A2(new_n774), .A3(new_n778), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT103), .B(KEYINPUT23), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n755), .A2(G20), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G299), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1956), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G4), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n633), .B2(G16), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G1348), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI22_X1  g374(.A1(new_n796), .A2(G1348), .B1(new_n793), .B2(new_n792), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n788), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n769), .A2(new_n770), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n755), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n755), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1971), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G23), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT98), .Z(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G288), .B2(new_n755), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT33), .B(G1976), .Z(new_n809));
  XOR2_X1   g384(.A(new_n808), .B(new_n809), .Z(new_n810));
  MUX2_X1   g385(.A(G6), .B(G305), .S(G16), .Z(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT32), .B(G1981), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n805), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT34), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n755), .A2(G24), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n613), .B2(new_n755), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(G1986), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n725), .A2(G25), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n484), .A2(G131), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n823));
  INV_X1    g398(.A(G107), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(G2105), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n491), .B2(G119), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n821), .B1(new_n828), .B2(new_n725), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT35), .B(G1991), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT97), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n829), .B(new_n831), .Z(new_n832));
  NOR2_X1   g407(.A1(new_n819), .A2(G1986), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n820), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n816), .A2(new_n817), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT36), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n835), .A2(KEYINPUT36), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n802), .B1(new_n836), .B2(new_n837), .ZN(G311));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n836), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n839), .A2(new_n770), .A3(new_n769), .A4(new_n801), .ZN(G150));
  NAND2_X1  g415(.A1(new_n633), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  INV_X1    g417(.A(G55), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n544), .B2(new_n545), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(G80), .A2(G543), .ZN(new_n846));
  INV_X1    g421(.A(G67), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n524), .B2(new_n847), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n525), .A2(G93), .B1(G651), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n556), .A2(new_n845), .A3(new_n560), .A4(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n560), .ZN(new_n851));
  INV_X1    g426(.A(new_n849), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n555), .A2(new_n851), .B1(new_n844), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n842), .B(new_n854), .Z(new_n855));
  OR2_X1    g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT104), .B(G860), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n845), .B2(new_n849), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(G145));
  NAND2_X1  g437(.A1(new_n506), .A2(new_n507), .ZN(new_n863));
  INV_X1    g438(.A(new_n502), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n499), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT106), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n865), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT107), .B1(new_n508), .B2(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n785), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n741), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(new_n723), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n724), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n491), .A2(G130), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n496), .A2(G118), .ZN(new_n881));
  OAI21_X1  g456(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n484), .B2(G142), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n827), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n643), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n877), .A2(new_n878), .A3(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n493), .B(new_n652), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT105), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n481), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(G37), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n886), .B1(new_n877), .B2(new_n878), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n896), .A2(KEYINPUT108), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n889), .B(new_n893), .C1(new_n896), .C2(KEYINPUT108), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g475(.A1(G290), .A2(G166), .ZN(new_n901));
  XOR2_X1   g476(.A(G305), .B(G288), .Z(new_n902));
  NOR2_X1   g477(.A1(new_n613), .A2(new_n531), .ZN(new_n903));
  OR3_X1    g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT42), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n636), .B(new_n854), .ZN(new_n908));
  INV_X1    g483(.A(G299), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n625), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n633), .A2(G299), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(new_n633), .B2(G299), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(KEYINPUT109), .A3(new_n625), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n916), .A3(new_n911), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n633), .B2(G299), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n917), .A2(new_n918), .B1(new_n910), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n913), .B1(new_n920), .B2(new_n908), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT110), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n907), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n924));
  INV_X1    g499(.A(new_n921), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n907), .A2(new_n925), .A3(new_n924), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n626), .B1(new_n844), .B2(new_n852), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(G295));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n929), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n917), .A2(new_n918), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n919), .A2(new_n910), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n936));
  NAND2_X1  g511(.A1(G168), .A2(G171), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n541), .A2(new_n546), .B1(new_n549), .B2(new_n552), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n854), .A3(KEYINPUT111), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n854), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n937), .A2(new_n850), .A3(new_n853), .A4(new_n938), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n935), .A2(new_n936), .A3(new_n940), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n943), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n912), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(new_n940), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT112), .B1(new_n920), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n906), .ZN(new_n952));
  AOI21_X1  g527(.A(G37), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n945), .A2(new_n950), .A3(new_n906), .A4(new_n948), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n932), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n944), .A2(new_n940), .B1(new_n911), .B2(new_n910), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n915), .A2(new_n916), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n958), .A2(new_n919), .B1(new_n918), .B2(new_n912), .ZN(new_n959));
  OAI22_X1  g534(.A1(new_n956), .A2(new_n957), .B1(new_n959), .B2(new_n947), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n956), .A2(new_n957), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n952), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G37), .ZN(new_n963));
  AND4_X1   g538(.A1(new_n932), .A2(new_n962), .A3(new_n963), .A4(new_n954), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n955), .A2(new_n964), .A3(KEYINPUT44), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n963), .A3(new_n954), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n953), .A2(new_n932), .A3(new_n954), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n965), .A2(new_n970), .ZN(G397));
  XOR2_X1   g546(.A(new_n785), .B(G2067), .Z(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(G1996), .B2(new_n741), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n874), .A2(G1384), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n471), .A2(new_n480), .A3(G40), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n974), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(G1996), .A3(new_n741), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n827), .B(new_n831), .Z(new_n984));
  NAND2_X1  g559(.A1(new_n976), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n613), .B(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n976), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT120), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n865), .A2(new_n870), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n993), .B(new_n994), .C1(new_n508), .C2(new_n869), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT117), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n994), .B1(new_n500), .B2(new_n508), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n975), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n798), .ZN(new_n1002));
  INV_X1    g577(.A(new_n975), .ZN(new_n1003));
  AOI21_X1  g578(.A(G1384), .B1(new_n865), .B2(new_n870), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(G2067), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n990), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1348), .B1(new_n998), .B2(new_n1000), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1009), .A2(KEYINPUT120), .A3(new_n1006), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n499), .B(KEYINPUT70), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n865), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1003), .B1(new_n1013), .B2(KEYINPUT45), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n994), .A2(KEYINPUT45), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n872), .A2(new_n873), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT115), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n872), .A2(new_n873), .A3(new_n1018), .A4(new_n1015), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1014), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT56), .B(G2072), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n975), .B1(new_n1013), .B2(new_n993), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n993), .B2(new_n1004), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1020), .A2(new_n1021), .B1(new_n793), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT57), .B1(new_n587), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G299), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n579), .B(new_n587), .C1(new_n1025), .C2(KEYINPUT57), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1011), .A2(new_n633), .A3(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1024), .A2(KEYINPUT121), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1028), .B(new_n1027), .C1(new_n1024), .C2(KEYINPUT121), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT60), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1003), .B1(new_n1013), .B2(new_n993), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n997), .B2(new_n995), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n990), .B(new_n1007), .C1(new_n1037), .C2(G1348), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT120), .B1(new_n1009), .B2(new_n1006), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1035), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT123), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT60), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT123), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n625), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1040), .A2(KEYINPUT123), .A3(new_n633), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1041), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1011), .A2(new_n1035), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1996), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT58), .B(G1341), .Z(new_n1050));
  AOI22_X1  g625(.A1(new_n1020), .A2(new_n1049), .B1(new_n1005), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n561), .ZN(new_n1052));
  NAND2_X1  g627(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT61), .B(new_n1030), .C1(new_n1033), .C2(new_n1032), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1030), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1054), .A2(new_n1055), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1034), .B1(new_n1048), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n592), .A2(G8), .A3(new_n593), .ZN(new_n1062));
  NAND2_X1  g637(.A1(KEYINPUT118), .A2(KEYINPUT55), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n592), .A2(G8), .A3(new_n593), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1023), .A2(G2090), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1020), .A2(new_n1071), .ZN(new_n1072));
  AOI211_X1 g647(.A(KEYINPUT116), .B(new_n1014), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1971), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1070), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G8), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1069), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1072), .A2(new_n1073), .A3(G1971), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1001), .A2(G2090), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1068), .B(G8), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1005), .A2(G8), .ZN(new_n1082));
  XNOR2_X1  g657(.A(G305), .B(G1981), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT49), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1084), .B2(new_n1083), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1082), .ZN(new_n1087));
  INV_X1    g662(.A(G1976), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT52), .B1(G288), .B2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1087), .B(new_n1089), .C1(new_n1088), .C2(G288), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G288), .A2(new_n1088), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT52), .B1(new_n1082), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1086), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n998), .A2(new_n752), .A3(new_n1000), .ZN(new_n1095));
  OAI211_X1 g670(.A(KEYINPUT45), .B(new_n994), .C1(new_n500), .C2(new_n508), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n1003), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1004), .A2(KEYINPUT45), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n758), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1095), .A2(G168), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G8), .ZN(new_n1101));
  AOI21_X1  g676(.A(G168), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT51), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(new_n1104), .A3(G8), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  AND4_X1   g681(.A1(new_n1078), .A2(new_n1081), .A3(new_n1094), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n975), .A2(new_n1110), .A3(G2078), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1109), .B(new_n1111), .C1(KEYINPUT45), .C2(new_n974), .ZN(new_n1112));
  INV_X1    g687(.A(G1961), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1001), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G2078), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1117), .B2(new_n1110), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1118), .A2(G301), .ZN(new_n1119));
  OR4_X1    g694(.A1(new_n1110), .A2(new_n1097), .A3(new_n1098), .A4(G2078), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1114), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1117), .B2(new_n1110), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(G301), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1108), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1108), .B1(new_n1122), .B2(G301), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n1126));
  OAI21_X1  g701(.A(G171), .B1(new_n1118), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g702(.A(KEYINPUT124), .B(new_n1115), .C1(new_n1117), .C2(new_n1110), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1107), .A2(new_n1124), .A3(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1061), .A2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g706(.A(new_n1077), .B(G286), .C1(new_n1095), .C2(new_n1099), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1078), .A2(new_n1081), .A3(new_n1094), .A4(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(G8), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1069), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1132), .A2(KEYINPUT63), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1137), .A2(new_n1081), .A3(new_n1094), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G288), .A2(G1976), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1086), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(G305), .A2(G1981), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1087), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1081), .B2(new_n1093), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1106), .A2(KEYINPUT62), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1103), .A2(new_n1147), .A3(new_n1105), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1146), .A2(new_n1123), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1072), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1073), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1075), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1070), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1068), .B1(new_n1154), .B2(G8), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1081), .A2(new_n1094), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1145), .B1(new_n1149), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1140), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n989), .B1(new_n1131), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n976), .A2(new_n987), .A3(new_n613), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT126), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT48), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1163), .A2(new_n985), .A3(new_n983), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n972), .A2(new_n742), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n976), .A2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT125), .Z(new_n1167));
  NAND2_X1  g742(.A1(new_n976), .A2(new_n1049), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT46), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT47), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n828), .A2(new_n831), .ZN(new_n1172));
  OAI22_X1  g747(.A1(new_n982), .A2(new_n1172), .B1(G2067), .B2(new_n785), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1164), .B(new_n1171), .C1(new_n976), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1160), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1177));
  NOR2_X1   g751(.A1(G227), .A2(new_n460), .ZN(new_n1178));
  INV_X1    g752(.A(new_n1178), .ZN(new_n1179));
  OR3_X1    g753(.A1(G401), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g754(.A(new_n1177), .B1(G401), .B2(new_n1179), .ZN(new_n1181));
  AOI21_X1  g755(.A(G229), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g756(.A(new_n1182), .B(new_n899), .C1(new_n955), .C2(new_n964), .ZN(G225));
  INV_X1    g757(.A(G225), .ZN(G308));
endmodule


