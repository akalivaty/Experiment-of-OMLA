

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725;

  XNOR2_X1 U371 ( .A(n385), .B(KEYINPUT70), .ZN(n467) );
  INV_X1 U372 ( .A(KEYINPUT64), .ZN(n411) );
  NAND2_X1 U373 ( .A1(n383), .A2(n525), .ZN(n396) );
  XNOR2_X1 U374 ( .A(n393), .B(n531), .ZN(n379) );
  NOR2_X1 U375 ( .A1(n591), .A2(n692), .ZN(n592) );
  NOR2_X1 U376 ( .A1(n583), .A2(n692), .ZN(n585) );
  AND2_X2 U377 ( .A1(n693), .A2(n571), .ZN(n638) );
  XNOR2_X2 U378 ( .A(n429), .B(n428), .ZN(n542) );
  XNOR2_X2 U379 ( .A(n440), .B(G469), .ZN(n489) );
  AND2_X1 U380 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U381 ( .A1(n549), .A2(n548), .ZN(n552) );
  AND2_X1 U382 ( .A1(n524), .A2(n675), .ZN(n525) );
  INV_X1 U383 ( .A(KEYINPUT0), .ZN(n395) );
  XNOR2_X1 U384 ( .A(n562), .B(KEYINPUT84), .ZN(n568) );
  NAND2_X1 U385 ( .A1(n561), .A2(n560), .ZN(n562) );
  AND2_X1 U386 ( .A1(n379), .A2(n538), .ZN(n561) );
  AND2_X1 U387 ( .A1(n389), .A2(n386), .ZN(n510) );
  XNOR2_X1 U388 ( .A(n480), .B(KEYINPUT40), .ZN(n723) );
  AND2_X1 U389 ( .A1(n511), .A2(n629), .ZN(n480) );
  XNOR2_X1 U390 ( .A(n552), .B(n551), .ZN(n681) );
  OR2_X1 U391 ( .A1(n627), .A2(n490), .ZN(n491) );
  OR2_X1 U392 ( .A1(n580), .A2(G902), .ZN(n440) );
  XNOR2_X1 U393 ( .A(n411), .B(G953), .ZN(n417) );
  INV_X2 U394 ( .A(G101), .ZN(n370) );
  INV_X2 U395 ( .A(KEYINPUT74), .ZN(n368) );
  BUF_X1 U396 ( .A(n597), .Z(n350) );
  INV_X1 U397 ( .A(n644), .ZN(n351) );
  XNOR2_X1 U398 ( .A(n558), .B(n557), .ZN(n597) );
  XNOR2_X1 U399 ( .A(n489), .B(KEYINPUT1), .ZN(n512) );
  BUF_X1 U400 ( .A(n379), .Z(n352) );
  BUF_X1 U401 ( .A(n586), .Z(n353) );
  AND2_X2 U402 ( .A1(n541), .A2(n647), .ZN(n619) );
  XNOR2_X2 U403 ( .A(n570), .B(n569), .ZN(n693) );
  NOR2_X2 U404 ( .A1(n568), .A2(n567), .ZN(n570) );
  XNOR2_X2 U405 ( .A(n392), .B(n356), .ZN(n518) );
  INV_X1 U406 ( .A(G131), .ZN(n385) );
  XNOR2_X1 U407 ( .A(n711), .B(G146), .ZN(n439) );
  XNOR2_X1 U408 ( .A(n446), .B(n361), .ZN(n702) );
  XNOR2_X1 U409 ( .A(n445), .B(n444), .ZN(n361) );
  XNOR2_X1 U410 ( .A(G119), .B(G137), .ZN(n420) );
  XNOR2_X1 U411 ( .A(n419), .B(n418), .ZN(n459) );
  INV_X1 U412 ( .A(KEYINPUT8), .ZN(n418) );
  XNOR2_X1 U413 ( .A(n702), .B(n358), .ZN(n586) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n362), .B(n450), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n364), .B(n363), .ZN(n360) );
  INV_X1 U417 ( .A(KEYINPUT34), .ZN(n555) );
  XNOR2_X1 U418 ( .A(n427), .B(KEYINPUT25), .ZN(n428) );
  NOR2_X1 U419 ( .A1(n689), .A2(G902), .ZN(n429) );
  XNOR2_X1 U420 ( .A(KEYINPUT3), .B(G116), .ZN(n401) );
  NAND2_X1 U421 ( .A1(n388), .A2(n502), .ZN(n387) );
  INV_X1 U422 ( .A(n625), .ZN(n388) );
  XNOR2_X1 U423 ( .A(n462), .B(n384), .ZN(n711) );
  XNOR2_X1 U424 ( .A(n467), .B(n398), .ZN(n384) );
  XNOR2_X1 U425 ( .A(KEYINPUT4), .B(G137), .ZN(n398) );
  INV_X1 U426 ( .A(G953), .ZN(n521) );
  XNOR2_X1 U427 ( .A(n382), .B(G125), .ZN(n447) );
  INV_X1 U428 ( .A(G146), .ZN(n382) );
  XNOR2_X1 U429 ( .A(G143), .B(G128), .ZN(n448) );
  XNOR2_X1 U430 ( .A(G113), .B(G143), .ZN(n468) );
  XNOR2_X1 U431 ( .A(G122), .B(G104), .ZN(n469) );
  XNOR2_X1 U432 ( .A(n447), .B(n380), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n381), .B(KEYINPUT76), .ZN(n380) );
  INV_X1 U434 ( .A(KEYINPUT18), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n448), .B(n449), .ZN(n362) );
  XNOR2_X1 U436 ( .A(KEYINPUT4), .B(KEYINPUT87), .ZN(n449) );
  INV_X1 U437 ( .A(KEYINPUT30), .ZN(n390) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n643) );
  INV_X1 U439 ( .A(KEYINPUT69), .ZN(n376) );
  NAND2_X1 U440 ( .A1(n542), .A2(n378), .ZN(n377) );
  OR2_X1 U441 ( .A1(n607), .A2(G902), .ZN(n408) );
  XNOR2_X1 U442 ( .A(n448), .B(G134), .ZN(n462) );
  XNOR2_X1 U443 ( .A(n453), .B(n357), .ZN(n511) );
  NAND2_X1 U444 ( .A1(n518), .A2(n662), .ZN(n499) );
  AND2_X1 U445 ( .A1(n526), .A2(n378), .ZN(n527) );
  INV_X1 U446 ( .A(n542), .ZN(n647) );
  XNOR2_X1 U447 ( .A(n372), .B(n373), .ZN(n371) );
  XNOR2_X1 U448 ( .A(n375), .B(n555), .ZN(n374) );
  NOR2_X1 U449 ( .A1(n536), .A2(n553), .ZN(n354) );
  INV_X1 U450 ( .A(n648), .ZN(n378) );
  XOR2_X1 U451 ( .A(G110), .B(G128), .Z(n355) );
  AND2_X1 U452 ( .A1(G210), .A2(n451), .ZN(n356) );
  XOR2_X1 U453 ( .A(n452), .B(KEYINPUT73), .Z(n357) );
  XNOR2_X1 U454 ( .A(n371), .B(n709), .ZN(n689) );
  OR2_X1 U455 ( .A1(n713), .A2(G952), .ZN(n610) );
  NAND2_X1 U456 ( .A1(n713), .A2(G224), .ZN(n364) );
  XNOR2_X2 U457 ( .A(n365), .B(n402), .ZN(n446) );
  XNOR2_X2 U458 ( .A(n367), .B(n432), .ZN(n445) );
  XNOR2_X2 U459 ( .A(n369), .B(n399), .ZN(n365) );
  NOR2_X1 U460 ( .A1(n638), .A2(KEYINPUT2), .ZN(n366) );
  NOR2_X4 U461 ( .A1(n366), .A2(n578), .ZN(n688) );
  XNOR2_X2 U462 ( .A(n368), .B(G110), .ZN(n367) );
  XNOR2_X2 U463 ( .A(n370), .B(G113), .ZN(n369) );
  NAND2_X1 U464 ( .A1(n459), .A2(G221), .ZN(n373) );
  XNOR2_X1 U465 ( .A(n422), .B(n421), .ZN(n372) );
  NAND2_X1 U466 ( .A1(n374), .A2(n556), .ZN(n558) );
  NAND2_X1 U467 ( .A1(n681), .A2(n554), .ZN(n375) );
  INV_X1 U468 ( .A(n643), .ZN(n532) );
  XNOR2_X1 U469 ( .A(n352), .B(n721), .ZN(G3) );
  NAND2_X1 U470 ( .A1(n500), .A2(n383), .ZN(n626) );
  XNOR2_X2 U471 ( .A(n499), .B(KEYINPUT19), .ZN(n383) );
  NOR2_X1 U472 ( .A1(n634), .A2(n387), .ZN(n386) );
  XNOR2_X1 U473 ( .A(n488), .B(KEYINPUT46), .ZN(n389) );
  INV_X1 U474 ( .A(n651), .ZN(n483) );
  XNOR2_X1 U475 ( .A(n391), .B(n390), .ZN(n416) );
  NAND2_X1 U476 ( .A1(n651), .A2(n662), .ZN(n391) );
  XNOR2_X2 U477 ( .A(n408), .B(G472), .ZN(n651) );
  NAND2_X1 U478 ( .A1(n586), .A2(n576), .ZN(n392) );
  NAND2_X1 U479 ( .A1(n394), .A2(n542), .ZN(n393) );
  XNOR2_X1 U480 ( .A(n530), .B(KEYINPUT83), .ZN(n394) );
  INV_X1 U481 ( .A(n528), .ZN(n553) );
  XNOR2_X2 U482 ( .A(n396), .B(n395), .ZN(n528) );
  NOR2_X2 U483 ( .A1(n545), .A2(n351), .ZN(n539) );
  XNOR2_X1 U484 ( .A(KEYINPUT120), .B(n593), .ZN(n397) );
  AND2_X1 U485 ( .A1(n597), .A2(n563), .ZN(n564) );
  XNOR2_X2 U486 ( .A(KEYINPUT91), .B(G119), .ZN(n399) );
  INV_X1 U487 ( .A(KEYINPUT71), .ZN(n400) );
  XNOR2_X1 U488 ( .A(n401), .B(n400), .ZN(n402) );
  NOR2_X1 U489 ( .A1(G953), .A2(G237), .ZN(n473) );
  NAND2_X1 U490 ( .A1(n473), .A2(G210), .ZN(n403) );
  XNOR2_X1 U491 ( .A(n403), .B(KEYINPUT5), .ZN(n405) );
  XNOR2_X1 U492 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n404) );
  XNOR2_X1 U493 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U494 ( .A(n446), .B(n406), .ZN(n407) );
  XNOR2_X1 U495 ( .A(n439), .B(n407), .ZN(n607) );
  OR2_X1 U496 ( .A1(G237), .A2(G902), .ZN(n451) );
  NAND2_X1 U497 ( .A1(n451), .A2(G214), .ZN(n409) );
  XOR2_X1 U498 ( .A(KEYINPUT92), .B(n409), .Z(n513) );
  NAND2_X1 U499 ( .A1(G234), .A2(G237), .ZN(n410) );
  XNOR2_X1 U500 ( .A(n410), .B(KEYINPUT14), .ZN(n675) );
  BUF_X2 U501 ( .A(n417), .Z(n713) );
  NOR2_X1 U502 ( .A1(n713), .A2(G900), .ZN(n412) );
  NAND2_X1 U503 ( .A1(G902), .A2(n412), .ZN(n413) );
  NAND2_X1 U504 ( .A1(G952), .A2(n521), .ZN(n522) );
  NAND2_X1 U505 ( .A1(n413), .A2(n522), .ZN(n414) );
  NAND2_X1 U506 ( .A1(n675), .A2(n414), .ZN(n415) );
  XOR2_X1 U507 ( .A(KEYINPUT78), .B(n415), .Z(n481) );
  AND2_X1 U508 ( .A1(n416), .A2(n481), .ZN(n442) );
  NAND2_X1 U509 ( .A1(n417), .A2(G234), .ZN(n419) );
  XNOR2_X1 U510 ( .A(n355), .B(n420), .ZN(n422) );
  XOR2_X1 U511 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n421) );
  XNOR2_X1 U512 ( .A(G140), .B(KEYINPUT10), .ZN(n424) );
  INV_X1 U513 ( .A(n447), .ZN(n423) );
  XNOR2_X1 U514 ( .A(n424), .B(n423), .ZN(n709) );
  XNOR2_X1 U515 ( .A(KEYINPUT90), .B(KEYINPUT15), .ZN(n425) );
  XNOR2_X1 U516 ( .A(n425), .B(G902), .ZN(n576) );
  NAND2_X1 U517 ( .A1(n576), .A2(G234), .ZN(n426) );
  XNOR2_X1 U518 ( .A(KEYINPUT20), .B(n426), .ZN(n430) );
  NAND2_X1 U519 ( .A1(n430), .A2(G217), .ZN(n427) );
  NAND2_X1 U520 ( .A1(n430), .A2(G221), .ZN(n431) );
  XNOR2_X1 U521 ( .A(n431), .B(KEYINPUT21), .ZN(n648) );
  XNOR2_X2 U522 ( .A(G104), .B(G107), .ZN(n432) );
  XOR2_X1 U523 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n434) );
  XNOR2_X1 U524 ( .A(G101), .B(G140), .ZN(n433) );
  XNOR2_X1 U525 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U526 ( .A(n445), .B(n435), .Z(n437) );
  NAND2_X1 U527 ( .A1(G227), .A2(n713), .ZN(n436) );
  XNOR2_X1 U528 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U529 ( .A(n439), .B(n438), .ZN(n580) );
  INV_X1 U530 ( .A(n489), .ZN(n441) );
  NOR2_X1 U531 ( .A1(n643), .A2(n441), .ZN(n535) );
  NAND2_X1 U532 ( .A1(n442), .A2(n535), .ZN(n443) );
  XNOR2_X1 U533 ( .A(n443), .B(KEYINPUT75), .ZN(n503) );
  XOR2_X1 U534 ( .A(KEYINPUT16), .B(G122), .Z(n444) );
  XOR2_X1 U535 ( .A(KEYINPUT77), .B(KEYINPUT17), .Z(n450) );
  INV_X1 U536 ( .A(n518), .ZN(n509) );
  XNOR2_X1 U537 ( .A(KEYINPUT38), .B(n509), .ZN(n663) );
  NAND2_X1 U538 ( .A1(n503), .A2(n663), .ZN(n453) );
  XNOR2_X1 U539 ( .A(KEYINPUT82), .B(KEYINPUT39), .ZN(n452) );
  XNOR2_X1 U540 ( .A(G116), .B(G122), .ZN(n454) );
  XNOR2_X1 U541 ( .A(n454), .B(KEYINPUT7), .ZN(n458) );
  XOR2_X1 U542 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n456) );
  XNOR2_X1 U543 ( .A(G107), .B(KEYINPUT100), .ZN(n455) );
  XNOR2_X1 U544 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U545 ( .A(n458), .B(n457), .Z(n461) );
  NAND2_X1 U546 ( .A1(G217), .A2(n459), .ZN(n460) );
  XNOR2_X1 U547 ( .A(n461), .B(n460), .ZN(n463) );
  XNOR2_X1 U548 ( .A(n463), .B(n462), .ZN(n593) );
  INV_X1 U549 ( .A(G902), .ZN(n464) );
  NAND2_X1 U550 ( .A1(n593), .A2(n464), .ZN(n466) );
  INV_X1 U551 ( .A(G478), .ZN(n465) );
  XNOR2_X1 U552 ( .A(n466), .B(n465), .ZN(n504) );
  XNOR2_X1 U553 ( .A(n468), .B(n467), .ZN(n472) );
  XOR2_X1 U554 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n470) );
  XNOR2_X1 U555 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U556 ( .A(n472), .B(n471), .Z(n475) );
  NAND2_X1 U557 ( .A1(G214), .A2(n473), .ZN(n474) );
  XNOR2_X1 U558 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U559 ( .A(n476), .B(n709), .ZN(n600) );
  NOR2_X1 U560 ( .A1(n600), .A2(G902), .ZN(n479) );
  XOR2_X1 U561 ( .A(G475), .B(KEYINPUT98), .Z(n477) );
  XNOR2_X1 U562 ( .A(KEYINPUT13), .B(n477), .ZN(n478) );
  XNOR2_X1 U563 ( .A(n479), .B(n478), .ZN(n505) );
  XNOR2_X1 U564 ( .A(n505), .B(KEYINPUT99), .ZN(n496) );
  NAND2_X1 U565 ( .A1(n504), .A2(n496), .ZN(n627) );
  INV_X1 U566 ( .A(n627), .ZN(n629) );
  NOR2_X1 U567 ( .A1(n648), .A2(n542), .ZN(n482) );
  NAND2_X1 U568 ( .A1(n482), .A2(n481), .ZN(n490) );
  NOR2_X1 U569 ( .A1(n490), .A2(n483), .ZN(n484) );
  XNOR2_X1 U570 ( .A(n484), .B(KEYINPUT28), .ZN(n485) );
  NAND2_X1 U571 ( .A1(n485), .A2(n489), .ZN(n498) );
  INV_X1 U572 ( .A(n513), .ZN(n662) );
  NAND2_X1 U573 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U574 ( .A1(n505), .A2(n504), .ZN(n665) );
  NOR2_X1 U575 ( .A1(n666), .A2(n665), .ZN(n486) );
  XNOR2_X1 U576 ( .A(KEYINPUT41), .B(n486), .ZN(n679) );
  NOR2_X1 U577 ( .A1(n498), .A2(n679), .ZN(n487) );
  XNOR2_X1 U578 ( .A(n487), .B(KEYINPUT42), .ZN(n724) );
  NOR2_X1 U579 ( .A1(n723), .A2(n724), .ZN(n488) );
  INV_X1 U580 ( .A(n512), .ZN(n644) );
  XNOR2_X1 U581 ( .A(n651), .B(KEYINPUT6), .ZN(n548) );
  OR2_X1 U582 ( .A1(n548), .A2(n491), .ZN(n492) );
  XNOR2_X1 U583 ( .A(n492), .B(KEYINPUT107), .ZN(n515) );
  INV_X1 U584 ( .A(n515), .ZN(n493) );
  NOR2_X1 U585 ( .A1(n493), .A2(n499), .ZN(n494) );
  XOR2_X1 U586 ( .A(KEYINPUT36), .B(n494), .Z(n495) );
  NOR2_X1 U587 ( .A1(n644), .A2(n495), .ZN(n634) );
  NOR2_X1 U588 ( .A1(n496), .A2(n504), .ZN(n497) );
  XNOR2_X1 U589 ( .A(n497), .B(KEYINPUT102), .ZN(n632) );
  NOR2_X1 U590 ( .A1(n632), .A2(n629), .ZN(n667) );
  INV_X1 U591 ( .A(n498), .ZN(n500) );
  NOR2_X1 U592 ( .A1(n667), .A2(n626), .ZN(n501) );
  XNOR2_X1 U593 ( .A(n501), .B(KEYINPUT47), .ZN(n502) );
  OR2_X1 U594 ( .A1(n505), .A2(n504), .ZN(n507) );
  INV_X1 U595 ( .A(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U596 ( .A(n507), .B(n506), .ZN(n556) );
  NAND2_X1 U597 ( .A1(n503), .A2(n556), .ZN(n508) );
  NOR2_X1 U598 ( .A1(n509), .A2(n508), .ZN(n625) );
  XNOR2_X1 U599 ( .A(n510), .B(KEYINPUT48), .ZN(n708) );
  NAND2_X1 U600 ( .A1(n511), .A2(n632), .ZN(n636) );
  INV_X1 U601 ( .A(n636), .ZN(n520) );
  XOR2_X1 U602 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n517) );
  NOR2_X1 U603 ( .A1(n513), .A2(n351), .ZN(n514) );
  NAND2_X1 U604 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U605 ( .A(n517), .B(n516), .ZN(n519) );
  NOR2_X1 U606 ( .A1(n519), .A2(n518), .ZN(n637) );
  NOR2_X1 U607 ( .A1(n520), .A2(n637), .ZN(n707) );
  AND2_X1 U608 ( .A1(n708), .A2(n707), .ZN(n571) );
  NOR2_X1 U609 ( .A1(G898), .A2(n521), .ZN(n701) );
  NAND2_X1 U610 ( .A1(n701), .A2(G902), .ZN(n523) );
  NAND2_X1 U611 ( .A1(n523), .A2(n522), .ZN(n524) );
  INV_X1 U612 ( .A(n665), .ZN(n526) );
  NAND2_X1 U613 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U614 ( .A(n529), .B(KEYINPUT22), .ZN(n545) );
  NAND2_X1 U615 ( .A1(n539), .A2(n548), .ZN(n530) );
  INV_X1 U616 ( .A(KEYINPUT103), .ZN(n531) );
  NAND2_X1 U617 ( .A1(n532), .A2(n512), .ZN(n549) );
  OR2_X1 U618 ( .A1(n549), .A2(n483), .ZN(n656) );
  NOR2_X1 U619 ( .A1(n656), .A2(n553), .ZN(n534) );
  XNOR2_X1 U620 ( .A(KEYINPUT31), .B(KEYINPUT97), .ZN(n533) );
  XNOR2_X1 U621 ( .A(n534), .B(n533), .ZN(n631) );
  NAND2_X1 U622 ( .A1(n535), .A2(n483), .ZN(n536) );
  NOR2_X1 U623 ( .A1(n631), .A2(n354), .ZN(n537) );
  OR2_X1 U624 ( .A1(n537), .A2(n667), .ZN(n538) );
  NAND2_X1 U625 ( .A1(n539), .A2(n483), .ZN(n540) );
  XNOR2_X1 U626 ( .A(n540), .B(KEYINPUT65), .ZN(n541) );
  NOR2_X1 U627 ( .A1(n644), .A2(n542), .ZN(n543) );
  XOR2_X1 U628 ( .A(KEYINPUT104), .B(n543), .Z(n544) );
  NOR2_X1 U629 ( .A1(n545), .A2(n544), .ZN(n546) );
  AND2_X1 U630 ( .A1(n546), .A2(n548), .ZN(n547) );
  XNOR2_X1 U631 ( .A(n547), .B(KEYINPUT32), .ZN(n722) );
  NOR2_X2 U632 ( .A1(n619), .A2(n722), .ZN(n565) );
  XNOR2_X1 U633 ( .A(KEYINPUT105), .B(KEYINPUT33), .ZN(n550) );
  XNOR2_X1 U634 ( .A(n550), .B(KEYINPUT72), .ZN(n551) );
  INV_X1 U635 ( .A(n553), .ZN(n554) );
  INV_X1 U636 ( .A(KEYINPUT35), .ZN(n557) );
  NAND2_X1 U637 ( .A1(n565), .A2(n597), .ZN(n559) );
  NAND2_X1 U638 ( .A1(n559), .A2(KEYINPUT44), .ZN(n560) );
  INV_X1 U639 ( .A(KEYINPUT44), .ZN(n563) );
  XNOR2_X1 U640 ( .A(n564), .B(KEYINPUT68), .ZN(n566) );
  XNOR2_X1 U641 ( .A(KEYINPUT81), .B(KEYINPUT45), .ZN(n569) );
  NAND2_X1 U642 ( .A1(n636), .A2(KEYINPUT2), .ZN(n572) );
  XOR2_X1 U643 ( .A(n572), .B(KEYINPUT79), .Z(n573) );
  NOR2_X1 U644 ( .A1(n573), .A2(n637), .ZN(n574) );
  AND2_X1 U645 ( .A1(n708), .A2(n574), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n693), .A2(n575), .ZN(n641) );
  INV_X1 U647 ( .A(n576), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n641), .A2(n577), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n688), .A2(G469), .ZN(n582) );
  XOR2_X1 U650 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n579) );
  XNOR2_X1 U651 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U652 ( .A(n582), .B(n581), .ZN(n583) );
  INV_X1 U653 ( .A(n610), .ZN(n692) );
  INV_X1 U654 ( .A(KEYINPUT119), .ZN(n584) );
  XNOR2_X1 U655 ( .A(n585), .B(n584), .ZN(G54) );
  NAND2_X1 U656 ( .A1(n688), .A2(G210), .ZN(n590) );
  XNOR2_X1 U657 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n588) );
  XNOR2_X1 U658 ( .A(n353), .B(KEYINPUT86), .ZN(n587) );
  XNOR2_X1 U659 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U660 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U661 ( .A(n592), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U662 ( .A1(n688), .A2(G478), .ZN(n594) );
  XNOR2_X1 U663 ( .A(n594), .B(n397), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n595), .A2(n610), .ZN(n596) );
  XNOR2_X1 U665 ( .A(n596), .B(KEYINPUT121), .ZN(G63) );
  XNOR2_X1 U666 ( .A(n350), .B(G122), .ZN(G24) );
  NAND2_X1 U667 ( .A1(n688), .A2(G475), .ZN(n602) );
  XNOR2_X1 U668 ( .A(KEYINPUT66), .B(KEYINPUT88), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT59), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n600), .B(n599), .ZN(n601) );
  XNOR2_X1 U671 ( .A(n602), .B(n601), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n603), .A2(n610), .ZN(n605) );
  XNOR2_X1 U673 ( .A(KEYINPUT67), .B(KEYINPUT60), .ZN(n604) );
  XNOR2_X1 U674 ( .A(n605), .B(n604), .ZN(G60) );
  NAND2_X1 U675 ( .A1(n688), .A2(G472), .ZN(n609) );
  XNOR2_X1 U676 ( .A(KEYINPUT109), .B(KEYINPUT62), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U678 ( .A(n609), .B(n608), .ZN(n611) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(n614) );
  XNOR2_X1 U680 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n612) );
  XNOR2_X1 U681 ( .A(n612), .B(KEYINPUT85), .ZN(n613) );
  XNOR2_X1 U682 ( .A(n614), .B(n613), .ZN(G57) );
  NAND2_X1 U683 ( .A1(n354), .A2(n629), .ZN(n615) );
  XNOR2_X1 U684 ( .A(n615), .B(G104), .ZN(G6) );
  XOR2_X1 U685 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n617) );
  NAND2_X1 U686 ( .A1(n354), .A2(n632), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U688 ( .A(G107), .B(n618), .ZN(G9) );
  XOR2_X1 U689 ( .A(G110), .B(n619), .Z(G12) );
  INV_X1 U690 ( .A(n632), .ZN(n620) );
  NOR2_X1 U691 ( .A1(n626), .A2(n620), .ZN(n624) );
  XOR2_X1 U692 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n622) );
  XNOR2_X1 U693 ( .A(G128), .B(KEYINPUT112), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n624), .B(n623), .ZN(G30) );
  XOR2_X1 U696 ( .A(G143), .B(n625), .Z(G45) );
  NOR2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U698 ( .A(G146), .B(n628), .Z(G48) );
  NAND2_X1 U699 ( .A1(n631), .A2(n629), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(G113), .ZN(G15) );
  NAND2_X1 U701 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n633), .B(G116), .ZN(G18) );
  XNOR2_X1 U703 ( .A(G125), .B(n634), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n635), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U705 ( .A(G134), .B(n636), .ZN(G36) );
  XOR2_X1 U706 ( .A(G140), .B(n637), .Z(G42) );
  INV_X1 U707 ( .A(n638), .ZN(n640) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n639) );
  NAND2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n642) );
  AND2_X1 U710 ( .A1(n642), .A2(n641), .ZN(n685) );
  XNOR2_X1 U711 ( .A(KEYINPUT51), .B(KEYINPUT116), .ZN(n659) );
  XOR2_X1 U712 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n646) );
  NAND2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n646), .B(n645), .ZN(n655) );
  XOR2_X1 U715 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n650) );
  NAND2_X1 U716 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U717 ( .A(n650), .B(n649), .ZN(n652) );
  NOR2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U719 ( .A(n653), .B(KEYINPUT114), .ZN(n654) );
  NAND2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U721 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U722 ( .A(n659), .B(n658), .ZN(n660) );
  NOR2_X1 U723 ( .A1(n679), .A2(n660), .ZN(n661) );
  XOR2_X1 U724 ( .A(KEYINPUT117), .B(n661), .Z(n673) );
  INV_X1 U725 ( .A(n681), .ZN(n671) );
  NOR2_X1 U726 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U727 ( .A1(n665), .A2(n664), .ZN(n669) );
  NOR2_X1 U728 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U729 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U730 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U731 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U732 ( .A(KEYINPUT52), .B(n674), .ZN(n677) );
  NAND2_X1 U733 ( .A1(G952), .A2(n675), .ZN(n676) );
  NOR2_X1 U734 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U735 ( .A1(G953), .A2(n678), .ZN(n683) );
  INV_X1 U736 ( .A(n679), .ZN(n680) );
  NAND2_X1 U737 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U738 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U739 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U740 ( .A(n686), .B(KEYINPUT53), .ZN(n687) );
  XNOR2_X1 U741 ( .A(n687), .B(KEYINPUT118), .ZN(G75) );
  NAND2_X1 U742 ( .A1(n688), .A2(G217), .ZN(n690) );
  XNOR2_X1 U743 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U744 ( .A1(n692), .A2(n691), .ZN(G66) );
  INV_X1 U745 ( .A(n693), .ZN(n694) );
  NOR2_X1 U746 ( .A1(n694), .A2(G953), .ZN(n700) );
  NAND2_X1 U747 ( .A1(G224), .A2(G953), .ZN(n695) );
  XNOR2_X1 U748 ( .A(n695), .B(KEYINPUT122), .ZN(n696) );
  XNOR2_X1 U749 ( .A(KEYINPUT61), .B(n696), .ZN(n697) );
  NAND2_X1 U750 ( .A1(n697), .A2(G898), .ZN(n698) );
  XNOR2_X1 U751 ( .A(n698), .B(KEYINPUT123), .ZN(n699) );
  NOR2_X1 U752 ( .A1(n700), .A2(n699), .ZN(n706) );
  XNOR2_X1 U753 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n704) );
  NOR2_X1 U754 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U755 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U756 ( .A(n706), .B(n705), .ZN(G69) );
  NAND2_X1 U757 ( .A1(n708), .A2(n707), .ZN(n712) );
  XNOR2_X1 U758 ( .A(n709), .B(KEYINPUT93), .ZN(n710) );
  XOR2_X1 U759 ( .A(n711), .B(n710), .Z(n716) );
  XNOR2_X1 U760 ( .A(n712), .B(n716), .ZN(n714) );
  NAND2_X1 U761 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U762 ( .A(n715), .B(KEYINPUT126), .ZN(n720) );
  XNOR2_X1 U763 ( .A(G227), .B(n716), .ZN(n717) );
  NAND2_X1 U764 ( .A1(n717), .A2(G900), .ZN(n718) );
  NAND2_X1 U765 ( .A1(G953), .A2(n718), .ZN(n719) );
  NAND2_X1 U766 ( .A1(n720), .A2(n719), .ZN(G72) );
  XNOR2_X1 U767 ( .A(G101), .B(KEYINPUT110), .ZN(n721) );
  XOR2_X1 U768 ( .A(G119), .B(n722), .Z(G21) );
  XOR2_X1 U769 ( .A(n723), .B(G131), .Z(G33) );
  XNOR2_X1 U770 ( .A(G137), .B(KEYINPUT127), .ZN(n725) );
  XNOR2_X1 U771 ( .A(n725), .B(n724), .ZN(G39) );
endmodule

