//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT15), .ZN(new_n204));
  NOR2_X1   g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G29gat), .A2(G36gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n205), .B1(KEYINPUT14), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  NOR3_X1   g007(.A1(new_n208), .A2(G29gat), .A3(G36gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n204), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n206), .A2(KEYINPUT14), .ZN(new_n211));
  OR2_X1    g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n205), .A2(KEYINPUT14), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(KEYINPUT15), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n203), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n207), .A2(new_n204), .A3(new_n209), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(new_n202), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT17), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G15gat), .ZN(new_n220));
  INV_X1    g019(.A(G22gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G15gat), .A2(G22gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT16), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n224), .A2(G1gat), .A3(G8gat), .ZN(new_n225));
  INV_X1    g024(.A(G8gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n227));
  AND2_X1   g026(.A1(G15gat), .A2(G22gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G15gat), .A2(G22gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G1gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n226), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n228), .A2(new_n229), .ZN(new_n233));
  OAI22_X1  g032(.A1(new_n225), .A2(new_n232), .B1(KEYINPUT88), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(G8gat), .B1(new_n224), .B2(G1gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n233), .A2(KEYINPUT88), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n230), .A2(new_n231), .A3(new_n226), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT15), .B1(new_n213), .B2(new_n214), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n202), .B1(new_n217), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n215), .A2(new_n203), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n219), .A2(new_n239), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT89), .ZN(new_n246));
  INV_X1    g045(.A(new_n239), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n216), .A2(new_n218), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT89), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n219), .A2(new_n239), .A3(new_n244), .A4(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n246), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT90), .ZN(new_n253));
  NAND2_X1  g052(.A1(G229gat), .A2(G233gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT18), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n246), .A2(new_n254), .A3(new_n249), .A4(new_n251), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(KEYINPUT90), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(KEYINPUT18), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n255), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n252), .A2(KEYINPUT92), .A3(KEYINPUT18), .A4(new_n254), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT92), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT18), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n263), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n247), .A2(new_n248), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n267), .A2(KEYINPUT93), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(KEYINPUT93), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n249), .A3(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n254), .B(KEYINPUT13), .Z(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n261), .A2(new_n266), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n274));
  XNOR2_X1  g073(.A(G113gat), .B(G141gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G169gat), .B(G197gat), .Z(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT12), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n261), .A2(new_n266), .A3(new_n279), .A4(new_n272), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n285));
  XNOR2_X1  g084(.A(G71gat), .B(G99gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G15gat), .B(G43gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  XNOR2_X1  g088(.A(G113gat), .B(G120gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(KEYINPUT1), .ZN(new_n291));
  INV_X1    g090(.A(G127gat), .ZN(new_n292));
  INV_X1    g091(.A(G134gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G127gat), .A2(G134gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n290), .A2(new_n300), .B1(new_n294), .B2(new_n295), .ZN(new_n301));
  INV_X1    g100(.A(G120gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G113gat), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT1), .B1(new_n303), .B2(KEYINPUT72), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n299), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(G113gat), .ZN(new_n306));
  INV_X1    g105(.A(G113gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G120gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n308), .A3(new_n300), .ZN(new_n309));
  AND4_X1   g108(.A1(new_n299), .A2(new_n304), .A3(new_n296), .A4(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n298), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(KEYINPUT23), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(KEYINPUT23), .B2(new_n312), .ZN(new_n315));
  NAND3_X1  g114(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT24), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT67), .B(G190gat), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n316), .B(new_n319), .C1(new_n320), .C2(G183gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n315), .A2(KEYINPUT25), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G169gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT65), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT65), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G169gat), .ZN(new_n326));
  AOI21_X1  g125(.A(G176gat), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n314), .B1(new_n327), .B2(KEYINPUT23), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT64), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n319), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT64), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n330), .A2(new_n316), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT25), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT66), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n339));
  AOI211_X1 g138(.A(new_n339), .B(KEYINPUT25), .C1(new_n328), .C2(new_n335), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n322), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n343), .B(new_n322), .C1(new_n338), .C2(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n312), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(KEYINPUT26), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT26), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n313), .B1(new_n312), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n317), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT71), .ZN(new_n351));
  XOR2_X1   g150(.A(KEYINPUT27), .B(G183gat), .Z(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT69), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT69), .ZN(new_n354));
  INV_X1    g153(.A(G183gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(KEYINPUT27), .ZN(new_n356));
  INV_X1    g155(.A(new_n320), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT70), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n353), .A2(KEYINPUT70), .A3(new_n356), .A4(new_n357), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT28), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  OR3_X1    g162(.A1(new_n352), .A2(new_n362), .A3(new_n320), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n351), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n311), .B1(new_n345), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n304), .A2(new_n296), .A3(new_n309), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT73), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n301), .A2(new_n299), .A3(new_n304), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n297), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI211_X1 g170(.A(new_n371), .B(new_n365), .C1(new_n342), .C2(new_n344), .ZN(new_n372));
  INV_X1    g171(.A(G227gat), .ZN(new_n373));
  INV_X1    g172(.A(G233gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n367), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n289), .B1(new_n377), .B2(KEYINPUT33), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n324), .A2(new_n326), .ZN(new_n379));
  INV_X1    g178(.A(G176gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(KEYINPUT23), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n314), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n316), .B1(new_n333), .B2(KEYINPUT64), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n317), .A2(KEYINPUT64), .A3(new_n318), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n384), .A2(new_n385), .A3(new_n331), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n337), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n339), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n336), .A2(KEYINPUT66), .A3(new_n337), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n343), .B1(new_n390), .B2(new_n322), .ZN(new_n391));
  INV_X1    g190(.A(new_n344), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n366), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n371), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n365), .B1(new_n342), .B2(new_n344), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n311), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n375), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT34), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n397), .A2(KEYINPUT32), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n397), .B2(KEYINPUT32), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n375), .B1(new_n394), .B2(new_n396), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n401), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT32), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT34), .B1(new_n377), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n397), .A2(KEYINPUT32), .A3(new_n398), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n378), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n401), .B1(new_n399), .B2(new_n400), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n405), .A2(new_n406), .A3(new_n403), .ZN(new_n410));
  INV_X1    g209(.A(new_n378), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G57gat), .ZN(new_n415));
  INV_X1    g214(.A(G85gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT78), .ZN(new_n419));
  INV_X1    g218(.A(G141gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G148gat), .ZN(new_n421));
  INV_X1    g220(.A(G148gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G141gat), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n419), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G155gat), .B(G162gat), .ZN(new_n425));
  INV_X1    g224(.A(G155gat), .ZN(new_n426));
  INV_X1    g225(.A(G162gat), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT2), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n424), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n425), .B1(new_n424), .B2(new_n428), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT3), .B1(new_n429), .B2(new_n430), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n311), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT5), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n371), .B2(new_n431), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n369), .A2(new_n370), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n442), .A2(new_n431), .A3(new_n440), .A4(new_n298), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(KEYINPUT80), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n443), .B2(KEYINPUT80), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n441), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n447), .ZN(new_n449));
  INV_X1    g248(.A(new_n441), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n445), .ZN(new_n451));
  AOI211_X1 g250(.A(new_n436), .B(new_n439), .C1(new_n448), .C2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n431), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n311), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n371), .A2(new_n431), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n437), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n438), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n443), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n437), .B(new_n435), .C1(new_n459), .C2(new_n441), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n458), .A2(new_n460), .A3(KEYINPUT79), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT79), .B1(new_n458), .B2(new_n460), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n418), .B1(new_n452), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n458), .A2(new_n460), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT79), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n458), .A2(new_n460), .A3(KEYINPUT79), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n448), .A2(new_n451), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n435), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n469), .B(new_n417), .C1(new_n471), .C2(new_n439), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n464), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(KEYINPUT6), .B(new_n418), .C1(new_n452), .C2(new_n463), .ZN(new_n475));
  XNOR2_X1  g274(.A(G8gat), .B(G36gat), .ZN(new_n476));
  INV_X1    g275(.A(G64gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G92gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n481));
  INV_X1    g280(.A(G211gat), .ZN(new_n482));
  INV_X1    g281(.A(G218gat), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G197gat), .B(G204gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XOR2_X1   g285(.A(G211gat), .B(G218gat), .Z(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n487), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n489), .A3(new_n485), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT77), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(G226gat), .A2(G233gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n366), .A2(new_n341), .A3(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(KEYINPUT29), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n493), .B(new_n495), .C1(new_n395), .C2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n345), .A2(new_n366), .A3(new_n494), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n366), .A2(new_n341), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n496), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n491), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n480), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n480), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n395), .A2(new_n494), .B1(new_n501), .B2(new_n496), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n498), .B(new_n505), .C1(new_n506), .C2(new_n491), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(KEYINPUT30), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n503), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n505), .A4(new_n498), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n474), .A2(new_n475), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(G228gat), .A2(G233gat), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT29), .B1(new_n488), .B2(new_n490), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n453), .B1(new_n514), .B2(KEYINPUT3), .ZN(new_n515));
  INV_X1    g314(.A(new_n433), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(KEYINPUT29), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n513), .B(new_n515), .C1(new_n492), .C2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n491), .B1(new_n516), .B2(KEYINPUT29), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n513), .B1(new_n519), .B2(new_n515), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT83), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI211_X1 g321(.A(KEYINPUT83), .B(new_n513), .C1(new_n519), .C2(new_n515), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n221), .B(new_n518), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT84), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(G22gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n528));
  INV_X1    g327(.A(G50gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(G78gat), .B(G106gat), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  AND4_X1   g331(.A1(new_n524), .A2(new_n525), .A3(new_n527), .A4(new_n532), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n525), .A2(new_n532), .B1(new_n527), .B2(new_n524), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n408), .A2(new_n412), .A3(new_n512), .A4(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT35), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n409), .A2(new_n411), .A3(new_n410), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n411), .B1(new_n409), .B2(new_n410), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n408), .A2(KEYINPUT36), .A3(new_n412), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n508), .A2(new_n511), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n454), .A2(new_n455), .A3(new_n437), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n436), .B1(new_n448), .B2(new_n451), .ZN(new_n547));
  OAI211_X1 g346(.A(KEYINPUT39), .B(new_n546), .C1(new_n547), .C2(new_n437), .ZN(new_n548));
  XOR2_X1   g347(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n549));
  NAND3_X1  g348(.A1(new_n471), .A2(new_n457), .A3(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n548), .A2(new_n550), .A3(KEYINPUT40), .A4(new_n417), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n551), .A2(new_n464), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n550), .A3(new_n417), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT40), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n545), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n498), .B1(new_n506), .B2(new_n491), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT86), .B1(new_n557), .B2(KEYINPUT37), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT86), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n509), .A2(new_n559), .A3(new_n560), .A4(new_n498), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(KEYINPUT37), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n558), .A2(new_n561), .A3(new_n562), .A4(new_n480), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT38), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n507), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n561), .A3(new_n480), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT38), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n495), .B1(new_n395), .B2(new_n497), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n491), .A2(new_n506), .B1(new_n568), .B2(new_n492), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n569), .B2(new_n560), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n475), .B(new_n474), .C1(new_n566), .C2(new_n570), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n556), .B(new_n535), .C1(new_n565), .C2(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n512), .A2(new_n535), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n543), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n284), .B1(new_n537), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT105), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT102), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT8), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n416), .A2(new_n479), .ZN(new_n585));
  NAND4_X1  g384(.A1(KEYINPUT97), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n582), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G99gat), .B(G106gat), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g388(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n416), .B2(new_n479), .ZN(new_n590));
  XNOR2_X1  g389(.A(G99gat), .B(G106gat), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n590), .A2(new_n591), .A3(new_n582), .A4(new_n586), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n589), .A2(KEYINPUT98), .A3(new_n592), .ZN(new_n593));
  OR3_X1    g392(.A1(new_n587), .A2(KEYINPUT98), .A3(new_n588), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT99), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT9), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(G71gat), .A2(G78gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(KEYINPUT94), .A2(new_n602), .B1(new_n603), .B2(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n477), .A2(G57gat), .ZN(new_n605));
  INV_X1    g404(.A(G57gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(G64gat), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT94), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n605), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n606), .A2(G64gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n477), .A2(G57gat), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT9), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n603), .A2(new_n600), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n604), .A2(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n615), .A2(KEYINPUT10), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n579), .B1(new_n599), .B2(new_n616), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT99), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT99), .B1(new_n593), .B2(new_n594), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n579), .B(new_n616), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n615), .B1(new_n593), .B2(new_n594), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n589), .A2(new_n592), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n625), .A2(new_n615), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n623), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT101), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n629), .B(new_n623), .C1(new_n624), .C2(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n578), .B1(new_n622), .B2(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n624), .A2(new_n626), .A3(new_n576), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n576), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n622), .B2(new_n631), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n633), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n615), .A2(KEYINPUT21), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n239), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G183gat), .B(G211gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n426), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G127gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n652), .B(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n615), .A2(KEYINPUT21), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n652), .A2(new_n655), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n652), .A2(new_n655), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(G232gat), .A2(G233gat), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(KEYINPUT41), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G162gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n597), .A2(new_n219), .A3(new_n598), .A4(new_n244), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n670), .A2(new_n671), .B1(KEYINPUT41), .B2(new_n666), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n599), .A2(new_n248), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n618), .A2(new_n619), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n674), .A2(KEYINPUT100), .A3(new_n219), .A4(new_n244), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(G134gat), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n672), .A2(new_n675), .A3(new_n293), .A4(new_n673), .ZN(new_n678));
  XNOR2_X1  g477(.A(G190gat), .B(G218gat), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n680), .B1(new_n677), .B2(new_n678), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n669), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n683), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(new_n668), .A3(new_n681), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n665), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n575), .A2(new_n646), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n474), .A2(new_n475), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(new_n231), .ZN(G1324gat));
  NOR2_X1   g491(.A1(new_n689), .A2(new_n544), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n227), .A2(new_n226), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n698), .A2(new_n700), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT42), .B1(new_n693), .B2(new_n226), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT106), .B1(new_n703), .B2(new_n698), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n701), .B1(new_n702), .B2(new_n704), .ZN(G1325gat));
  NOR3_X1   g504(.A1(new_n689), .A2(new_n220), .A3(new_n543), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n537), .A2(new_n574), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n707), .A2(new_n283), .A3(new_n688), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n539), .A2(new_n540), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n646), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n706), .B1(new_n710), .B2(new_n220), .ZN(G1326gat));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713));
  INV_X1    g512(.A(new_n535), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n708), .A2(new_n713), .A3(new_n646), .A4(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT107), .B1(new_n689), .B2(new_n535), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n715), .A2(new_n716), .A3(new_n712), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(G22gat), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n719), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n221), .B1(new_n721), .B2(new_n717), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(G1327gat));
  NAND3_X1  g522(.A1(new_n665), .A2(new_n646), .A3(new_n687), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT108), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n724), .A2(KEYINPUT108), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n707), .A2(new_n283), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n727), .A2(G29gat), .A3(new_n690), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT45), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n665), .B(KEYINPUT109), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n645), .B(KEYINPUT110), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n707), .B2(new_n687), .ZN(new_n735));
  INV_X1    g534(.A(new_n687), .ZN(new_n736));
  AOI211_X1 g535(.A(KEYINPUT44), .B(new_n736), .C1(new_n537), .C2(new_n574), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n283), .B(new_n733), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n690), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n729), .A2(new_n739), .ZN(G1328gat));
  NOR3_X1   g539(.A1(new_n727), .A2(G36gat), .A3(new_n544), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G36gat), .B1(new_n738), .B2(new_n544), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n742), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(G1329gat));
  OAI21_X1  g545(.A(G43gat), .B1(new_n738), .B2(new_n543), .ZN(new_n747));
  INV_X1    g546(.A(new_n709), .ZN(new_n748));
  OR3_X1    g547(.A1(new_n727), .A2(G43gat), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n747), .A2(KEYINPUT47), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1330gat));
  OAI21_X1  g553(.A(G50gat), .B1(new_n738), .B2(new_n535), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n575), .A2(KEYINPUT112), .A3(new_n725), .A4(new_n726), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(new_n529), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n535), .B1(new_n727), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g560(.A1(KEYINPUT111), .A2(KEYINPUT48), .ZN(new_n762));
  NAND2_X1  g561(.A1(KEYINPUT111), .A2(KEYINPUT48), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  AND4_X1   g563(.A1(KEYINPUT113), .A2(new_n759), .A3(new_n529), .A4(new_n756), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT113), .B1(new_n757), .B2(new_n759), .ZN(new_n766));
  OAI211_X1 g565(.A(KEYINPUT48), .B(new_n755), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(G1331gat));
  INV_X1    g567(.A(new_n732), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n537), .B2(new_n574), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n665), .A2(new_n687), .A3(new_n283), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n690), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(new_n606), .ZN(G1332gat));
  INV_X1    g573(.A(new_n772), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n545), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT49), .B(G64gat), .Z(new_n777));
  OR2_X1    g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT114), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n782), .A3(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1333gat));
  INV_X1    g583(.A(new_n543), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n775), .A2(G71gat), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n772), .A2(new_n748), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(G71gat), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g588(.A1(new_n772), .A2(new_n535), .ZN(new_n790));
  XOR2_X1   g589(.A(KEYINPUT115), .B(G78gat), .Z(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1335gat));
  INV_X1    g591(.A(new_n665), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n283), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n707), .A2(new_n687), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n707), .A2(KEYINPUT51), .A3(new_n687), .A4(new_n794), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(KEYINPUT117), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n798), .A2(KEYINPUT117), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n690), .A2(new_n646), .A3(G85gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n794), .A2(new_n645), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT116), .Z(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n707), .A2(new_n687), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT44), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n707), .A2(new_n734), .A3(new_n687), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n690), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n802), .B1(new_n811), .B2(new_n416), .ZN(G1336gat));
  NOR3_X1   g611(.A1(new_n769), .A2(G92gat), .A3(new_n544), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n799), .A2(new_n800), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n545), .B(new_n804), .C1(new_n735), .C2(new_n737), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(new_n817), .B2(G92gat), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n799), .A2(new_n800), .A3(KEYINPUT118), .A4(new_n813), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n817), .A2(G92gat), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n797), .A2(new_n798), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n813), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT52), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n820), .A2(new_n824), .ZN(G1337gat));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n785), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G99gat), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n748), .A2(G99gat), .A3(new_n646), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n799), .A2(new_n800), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(G1338gat));
  NAND2_X1  g629(.A1(new_n809), .A2(new_n714), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(G106gat), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n769), .A2(G106gat), .A3(new_n535), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n799), .A2(new_n800), .A3(new_n835), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n831), .A2(G106gat), .B1(new_n822), .B2(new_n835), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n834), .A2(new_n836), .B1(new_n837), .B2(new_n833), .ZN(G1339gat));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT102), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n631), .A2(new_n578), .A3(new_n841), .A4(new_n620), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n843), .B2(new_n642), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n639), .B1(new_n632), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n628), .A2(new_n630), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n841), .A2(new_n620), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n576), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n849), .A2(KEYINPUT119), .A3(KEYINPUT54), .A4(new_n842), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n844), .A2(new_n846), .A3(KEYINPUT55), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n644), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT120), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n844), .A2(new_n846), .A3(new_n850), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n281), .A2(new_n282), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n851), .A2(new_n857), .A3(new_n644), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n853), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  OAI22_X1  g658(.A1(new_n270), .A2(new_n271), .B1(new_n254), .B2(new_n252), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n278), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n282), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n645), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n687), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n854), .A2(new_n855), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n862), .B1(new_n684), .B2(new_n686), .ZN(new_n867));
  AND4_X1   g666(.A1(new_n866), .A2(new_n867), .A3(new_n853), .A4(new_n858), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n730), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n771), .A2(new_n646), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n709), .A2(new_n535), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n869), .A2(KEYINPUT121), .A3(new_n870), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n545), .A2(new_n690), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n873), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n284), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(new_n307), .ZN(G1340gat));
  OAI21_X1  g679(.A(G120gat), .B1(new_n878), .B2(new_n769), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n645), .A2(new_n302), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n878), .B2(new_n882), .ZN(G1341gat));
  OR3_X1    g682(.A1(new_n878), .A2(new_n292), .A3(new_n730), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n292), .B1(new_n878), .B2(new_n665), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT122), .ZN(G1342gat));
  NOR3_X1   g686(.A1(new_n878), .A2(G134gat), .A3(new_n736), .ZN(new_n888));
  XOR2_X1   g687(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n889));
  OR2_X1    g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G134gat), .B1(new_n878), .B2(new_n736), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G1343gat));
  NAND2_X1  g692(.A1(new_n873), .A2(new_n876), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n543), .A2(new_n877), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n894), .A2(new_n535), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n284), .A2(G141gat), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n896), .A2(new_n897), .B1(KEYINPUT124), .B2(KEYINPUT58), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n873), .A2(new_n899), .A3(new_n714), .A4(new_n876), .ZN(new_n900));
  INV_X1    g699(.A(new_n852), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n856), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n687), .B1(new_n902), .B2(new_n864), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n868), .A2(new_n903), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n904), .A2(new_n665), .B1(new_n646), .B2(new_n771), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT57), .B1(new_n905), .B2(new_n535), .ZN(new_n906));
  INV_X1    g705(.A(new_n895), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n900), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G141gat), .B1(new_n908), .B2(new_n284), .ZN(new_n909));
  OR2_X1    g708(.A1(KEYINPUT124), .A2(KEYINPUT58), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n898), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n898), .B2(new_n909), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(G1344gat));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n422), .A3(new_n645), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(new_n908), .B2(new_n646), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(new_n422), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n873), .A2(KEYINPUT57), .A3(new_n714), .A4(new_n876), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n899), .B1(new_n905), .B2(new_n535), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n645), .A3(new_n907), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n915), .B1(new_n921), .B2(G148gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n914), .B1(new_n917), .B2(new_n922), .ZN(G1345gat));
  OAI21_X1  g722(.A(G155gat), .B1(new_n908), .B2(new_n730), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n896), .A2(new_n426), .A3(new_n793), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT125), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1346gat));
  OAI21_X1  g729(.A(G162gat), .B1(new_n908), .B2(new_n736), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n896), .A2(new_n427), .A3(new_n687), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1347gat));
  NOR3_X1   g732(.A1(new_n874), .A2(new_n810), .A3(new_n544), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n873), .A2(new_n876), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n283), .ZN(new_n936));
  MUX2_X1   g735(.A(new_n379), .B(G169gat), .S(new_n936), .Z(G1348gat));
  AOI21_X1  g736(.A(G176gat), .B1(new_n935), .B2(new_n645), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n769), .A2(new_n380), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n935), .B2(new_n939), .ZN(G1349gat));
  NAND4_X1  g739(.A1(new_n873), .A2(new_n731), .A3(new_n876), .A4(new_n934), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G183gat), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n665), .A2(new_n352), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n873), .A2(new_n876), .A3(new_n934), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n942), .A2(new_n947), .A3(new_n944), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n946), .A2(new_n948), .A3(KEYINPUT127), .A4(KEYINPUT60), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n942), .A2(new_n947), .A3(new_n944), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n947), .B1(new_n942), .B2(new_n944), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT60), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954));
  INV_X1    g753(.A(new_n945), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n952), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n949), .B1(new_n953), .B2(new_n956), .ZN(G1350gat));
  NAND2_X1  g756(.A1(new_n935), .A2(new_n687), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G190gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n958), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n961), .B(new_n962), .C1(new_n320), .C2(new_n958), .ZN(G1351gat));
  NOR2_X1   g762(.A1(new_n810), .A2(new_n544), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n543), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n965), .B1(new_n918), .B2(new_n919), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(G197gat), .B1(new_n967), .B2(new_n284), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n894), .A2(new_n535), .A3(new_n965), .ZN(new_n969));
  INV_X1    g768(.A(G197gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(new_n970), .A3(new_n283), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n971), .ZN(G1352gat));
  INV_X1    g771(.A(G204gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n969), .A2(new_n973), .A3(new_n645), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n975));
  OAI21_X1  g774(.A(G204gat), .B1(new_n967), .B2(new_n769), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(G1353gat));
  NAND3_X1  g777(.A1(new_n969), .A2(new_n482), .A3(new_n793), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n966), .A2(new_n793), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n980), .B2(G211gat), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT63), .ZN(new_n982));
  AOI211_X1 g781(.A(new_n982), .B(new_n482), .C1(new_n966), .C2(new_n793), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n979), .B1(new_n981), .B2(new_n983), .ZN(G1354gat));
  AOI21_X1  g783(.A(G218gat), .B1(new_n969), .B2(new_n687), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n736), .A2(new_n483), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(new_n966), .B2(new_n986), .ZN(G1355gat));
endmodule


