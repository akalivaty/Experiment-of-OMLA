//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT86), .ZN(new_n206));
  INV_X1    g005(.A(G22gat), .ZN(new_n207));
  NOR3_X1   g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n208), .B1(new_n207), .B2(new_n205), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT73), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(G197gat), .B(G204gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT22), .ZN(new_n214));
  INV_X1    g013(.A(G211gat), .ZN(new_n215));
  INV_X1    g014(.A(G218gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n212), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT73), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n213), .A2(new_n217), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT74), .B1(new_n222), .B2(new_n219), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n222), .A2(new_n219), .A3(KEYINPUT74), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT3), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G141gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT77), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT77), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G141gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n232), .A3(G148gat), .ZN(new_n233));
  INV_X1    g032(.A(G148gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G141gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(G155gat), .A2(G162gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT2), .ZN(new_n238));
  NOR2_X1   g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n229), .A2(G148gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n238), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n237), .A2(new_n239), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n236), .A2(new_n241), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(G228gat), .B(G233gat), .C1(new_n228), .C2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT84), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n250), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n237), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n239), .A2(new_n238), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n233), .A2(new_n235), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G155gat), .B(G162gat), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(new_n238), .B2(new_n243), .ZN(new_n257));
  NOR4_X1   g056(.A1(new_n255), .A2(new_n257), .A3(KEYINPUT78), .A4(KEYINPUT3), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n227), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n226), .B1(new_n259), .B2(KEYINPUT83), .ZN(new_n260));
  XNOR2_X1  g059(.A(G141gat), .B(G148gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n245), .B1(new_n261), .B2(KEYINPUT2), .ZN(new_n262));
  INV_X1    g061(.A(new_n235), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT77), .B(G141gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(G148gat), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n251), .B(new_n262), .C1(new_n265), .C2(new_n240), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT78), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n236), .A2(new_n241), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n268), .A2(new_n250), .A3(new_n251), .A4(new_n262), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT29), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT83), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n249), .B1(new_n260), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n225), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n274), .A2(new_n223), .B1(new_n220), .B2(new_n218), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(new_n270), .B2(new_n271), .ZN(new_n276));
  AOI211_X1 g075(.A(KEYINPUT83), .B(KEYINPUT29), .C1(new_n267), .C2(new_n269), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n276), .A2(KEYINPUT84), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n248), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT85), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT84), .B1(new_n276), .B2(new_n277), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n259), .A2(KEYINPUT83), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n283), .A2(new_n249), .A3(new_n275), .A4(new_n272), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT85), .A3(new_n248), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n274), .A2(new_n223), .B1(new_n219), .B2(new_n222), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n288), .A2(KEYINPUT29), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n246), .B1(new_n289), .B2(new_n251), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n270), .A2(new_n226), .ZN(new_n291));
  INV_X1    g090(.A(G228gat), .ZN(new_n292));
  INV_X1    g091(.A(G233gat), .ZN(new_n293));
  OAI22_X1  g092(.A1(new_n290), .A2(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n210), .B1(new_n287), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT85), .B1(new_n285), .B2(new_n248), .ZN(new_n296));
  AOI211_X1 g095(.A(new_n280), .B(new_n247), .C1(new_n282), .C2(new_n284), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n294), .B(new_n210), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR3_X1   g103(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT27), .B(G183gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(KEYINPUT68), .ZN(new_n309));
  INV_X1    g108(.A(G183gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT27), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT68), .ZN(new_n312));
  INV_X1    g111(.A(G190gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n307), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n308), .A2(KEYINPUT28), .A3(new_n313), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n306), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT65), .B(KEYINPUT25), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT24), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(G183gat), .A3(G190gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G183gat), .B(G190gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n322), .B2(new_n320), .ZN(new_n323));
  INV_X1    g122(.A(G169gat), .ZN(new_n324));
  INV_X1    g123(.A(G176gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT23), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(G169gat), .B2(G176gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n328), .A3(new_n303), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n319), .B1(new_n323), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n301), .A2(KEYINPUT24), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n310), .A2(G190gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n313), .A2(G183gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n331), .B1(new_n334), .B2(KEYINPUT24), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT67), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n303), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n326), .A2(new_n337), .A3(new_n328), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT25), .B1(new_n303), .B2(new_n336), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n330), .A2(KEYINPUT66), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT66), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n342), .B(new_n319), .C1(new_n323), .C2(new_n329), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n317), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G113gat), .B(G120gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n346), .B1(new_n347), .B2(KEYINPUT1), .ZN(new_n348));
  INV_X1    g147(.A(G120gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G113gat), .ZN(new_n350));
  INV_X1    g149(.A(G113gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G120gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  INV_X1    g153(.A(G134gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G127gat), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n348), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n357), .B1(new_n348), .B2(new_n356), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n306), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT27), .B(G183gat), .Z(new_n363));
  INV_X1    g162(.A(KEYINPUT68), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(G190gat), .B1(new_n311), .B2(KEYINPUT68), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT28), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n316), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n362), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n340), .A2(new_n335), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n326), .A2(new_n328), .A3(new_n303), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n318), .B1(new_n335), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n372), .B2(new_n342), .ZN(new_n373));
  INV_X1    g172(.A(new_n343), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n369), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n360), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT71), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT34), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n361), .A2(new_n377), .B1(G227gat), .B2(G233gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT34), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT71), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n379), .B(KEYINPUT64), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n378), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G71gat), .B(G99gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT70), .ZN(new_n392));
  INV_X1    g191(.A(G15gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(G43gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n361), .A2(new_n377), .A3(new_n387), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(KEYINPUT32), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n396), .B(KEYINPUT32), .C1(new_n397), .C2(new_n395), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n390), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n386), .A2(new_n389), .A3(new_n401), .A4(new_n400), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n300), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  NAND2_X1  g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(new_n344), .B2(KEYINPUT29), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT75), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n344), .A2(new_n412), .A3(new_n410), .ZN(new_n413));
  INV_X1    g212(.A(new_n410), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT75), .B1(new_n375), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n411), .B(new_n226), .C1(new_n413), .C2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n375), .B2(new_n227), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n330), .A2(KEYINPUT66), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(new_n343), .A3(new_n370), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n410), .B1(new_n419), .B2(new_n369), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n275), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n409), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n416), .A2(new_n421), .A3(new_n409), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n423), .B2(KEYINPUT30), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n416), .A2(new_n421), .A3(new_n409), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(KEYINPUT76), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT76), .B1(new_n425), .B2(new_n426), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT87), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n424), .B(new_n432), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT3), .B1(new_n255), .B2(new_n257), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n347), .A2(KEYINPUT1), .A3(G134gat), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n345), .B1(new_n353), .B2(new_n354), .ZN(new_n437));
  OAI21_X1  g236(.A(G127gat), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n348), .A2(new_n356), .A3(new_n357), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n267), .A2(new_n269), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G225gat), .A2(G233gat), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n262), .B1(new_n265), .B2(new_n240), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n438), .B2(new_n439), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n446), .B(new_n246), .C1(new_n358), .C2(new_n359), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n442), .B(new_n443), .C1(new_n447), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT79), .ZN(new_n451));
  INV_X1    g250(.A(new_n443), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n358), .A2(new_n246), .A3(new_n359), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(new_n445), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT5), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(KEYINPUT79), .A3(new_n455), .ZN(new_n458));
  XOR2_X1   g257(.A(G1gat), .B(G29gat), .Z(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G57gat), .B(G85gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n457), .A2(KEYINPUT6), .A3(new_n458), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n450), .A2(KEYINPUT79), .A3(new_n455), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n455), .B1(new_n450), .B2(KEYINPUT79), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n470), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n464), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT6), .B1(new_n470), .B2(new_n464), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n467), .A2(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(KEYINPUT35), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n406), .A2(new_n434), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT90), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n406), .A2(new_n434), .A3(new_n475), .A4(KEYINPUT90), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n474), .A2(new_n430), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n287), .A2(new_n294), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n209), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n298), .ZN(new_n483));
  INV_X1    g282(.A(new_n405), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n480), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n478), .A2(new_n479), .A3(new_n486), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n403), .A2(new_n404), .B1(KEYINPUT72), .B2(KEYINPUT36), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(new_n405), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n457), .A2(new_n458), .A3(new_n464), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n447), .A2(new_n449), .ZN(new_n493));
  INV_X1    g292(.A(new_n442), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n452), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OR3_X1    g294(.A1(new_n453), .A2(new_n445), .A3(new_n452), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(KEYINPUT39), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(new_n463), .C1(KEYINPUT39), .C2(new_n495), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n492), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT88), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(KEYINPUT88), .A3(new_n499), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n431), .A2(new_n505), .A3(new_n433), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n471), .A2(new_n467), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n409), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n416), .A2(new_n421), .ZN(new_n510));
  INV_X1    g309(.A(new_n409), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n508), .B1(new_n416), .B2(new_n421), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT38), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n473), .A2(new_n492), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n507), .A2(new_n514), .A3(new_n516), .A4(new_n425), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n411), .B1(new_n410), .B2(new_n344), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n508), .B1(new_n518), .B2(new_n226), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n411), .B(new_n275), .C1(new_n413), .C2(new_n415), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT38), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n521), .B(new_n522), .C1(new_n422), .C2(new_n509), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT38), .ZN(new_n524));
  INV_X1    g323(.A(new_n520), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n375), .A2(new_n227), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n420), .B1(new_n526), .B2(new_n410), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT37), .B1(new_n527), .B2(new_n275), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n524), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT89), .B1(new_n512), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n483), .B1(new_n517), .B2(new_n531), .ZN(new_n532));
  OAI221_X1 g331(.A(new_n491), .B1(new_n480), .B2(new_n483), .C1(new_n506), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n487), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT14), .ZN(new_n535));
  INV_X1    g334(.A(G36gat), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n535), .A2(new_n536), .A3(G29gat), .ZN(new_n537));
  INV_X1    g336(.A(G29gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(KEYINPUT91), .ZN(new_n543));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n543), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT92), .B(KEYINPUT15), .ZN(new_n547));
  OR3_X1    g346(.A1(new_n542), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G99gat), .B(G106gat), .Z(new_n551));
  INV_X1    g350(.A(KEYINPUT96), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT7), .ZN(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  INV_X1    g355(.A(G85gat), .ZN(new_n557));
  INV_X1    g356(.A(G92gat), .ZN(new_n558));
  AOI22_X1  g357(.A1(KEYINPUT8), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n553), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n551), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(KEYINPUT96), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(KEYINPUT96), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n563), .A2(new_n555), .A3(new_n553), .A4(new_n559), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n550), .A2(new_n565), .B1(KEYINPUT41), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n549), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n546), .A2(KEYINPUT17), .A3(new_n548), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n568), .B1(new_n573), .B2(new_n565), .ZN(new_n574));
  XOR2_X1   g373(.A(G190gat), .B(G218gat), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n567), .A2(KEYINPUT41), .ZN(new_n577));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n575), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n580), .B(new_n568), .C1(new_n573), .C2(new_n565), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n576), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n579), .B1(new_n576), .B2(new_n581), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(G57gat), .A2(G64gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G57gat), .A2(G64gat), .ZN(new_n586));
  AND2_X1   g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(KEYINPUT9), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n589));
  NOR2_X1   g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n587), .A2(new_n590), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n357), .ZN(new_n599));
  XNOR2_X1  g398(.A(G15gat), .B(G22gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT93), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT16), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n601), .B1(new_n602), .B2(G1gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n601), .A2(new_n602), .A3(G1gat), .ZN(new_n605));
  OAI221_X1 g404(.A(KEYINPUT94), .B1(G1gat), .B2(new_n600), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G8gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(KEYINPUT21), .B2(new_n595), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n599), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n612));
  INV_X1    g411(.A(G155gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n611), .A2(new_n617), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n584), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n571), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT17), .B1(new_n546), .B2(new_n548), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n608), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n550), .A2(new_n609), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT18), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n623), .A2(KEYINPUT18), .A3(new_n624), .A4(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n549), .A2(new_n608), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n624), .B(KEYINPUT13), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G197gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT11), .B(G169gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n628), .A2(new_n629), .A3(new_n639), .A4(new_n633), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n565), .A2(new_n595), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n562), .A2(new_n593), .A3(new_n564), .A4(new_n594), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n565), .A2(new_n595), .A3(KEYINPUT10), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n644), .A2(new_n646), .ZN(new_n652));
  INV_X1    g451(.A(new_n650), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n651), .A2(new_n654), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n620), .A2(new_n643), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n534), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n468), .A2(new_n469), .A3(new_n463), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT81), .B1(new_n666), .B2(KEYINPUT6), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n465), .A2(new_n466), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n516), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g470(.A1(new_n665), .A2(new_n434), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  AOI21_X1  g472(.A(KEYINPUT42), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT97), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(KEYINPUT42), .A3(new_n673), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n675), .B(new_n676), .C1(new_n607), .C2(new_n672), .ZN(G1325gat));
  OAI21_X1  g476(.A(G15gat), .B1(new_n665), .B2(new_n491), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n484), .A2(new_n393), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n665), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n483), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n534), .A2(new_n584), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n618), .A2(new_n619), .ZN(new_n685));
  INV_X1    g484(.A(new_n643), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n685), .A2(new_n686), .A3(new_n662), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR4_X1   g487(.A1(new_n684), .A2(G29gat), .A3(new_n669), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT45), .Z(new_n690));
  OAI21_X1  g489(.A(new_n491), .B1(new_n506), .B2(new_n532), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT98), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n480), .B2(new_n483), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n510), .A2(new_n511), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n416), .A2(KEYINPUT30), .A3(new_n421), .A4(new_n409), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT76), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(new_n423), .B2(KEYINPUT30), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n698), .B2(new_n427), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n669), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(new_n300), .A3(KEYINPUT98), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT99), .B1(new_n691), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n490), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n488), .B1(new_n484), .B2(new_n704), .ZN(new_n705));
  AND4_X1   g504(.A1(new_n507), .A2(new_n514), .A3(new_n516), .A4(new_n425), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n523), .A2(new_n530), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n300), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n431), .A2(new_n505), .A3(new_n433), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n700), .A2(new_n300), .A3(KEYINPUT98), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT98), .B1(new_n700), .B2(new_n300), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT99), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n710), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n476), .A2(new_n477), .B1(KEYINPUT35), .B2(new_n485), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n703), .A2(new_n715), .B1(new_n479), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n584), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(KEYINPUT44), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT100), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n691), .A2(new_n702), .A3(KEYINPUT99), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n714), .B1(new_n710), .B2(new_n713), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n487), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT100), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n725), .A3(new_n719), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n684), .A2(KEYINPUT44), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n721), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n687), .ZN(new_n729));
  OAI21_X1  g528(.A(G29gat), .B1(new_n729), .B2(new_n669), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n690), .A2(new_n730), .ZN(G1328gat));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(new_n534), .B2(new_n584), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n720), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(new_n725), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n688), .B1(new_n735), .B2(new_n721), .ZN(new_n736));
  INV_X1    g535(.A(new_n434), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n536), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n434), .A2(G36gat), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n534), .A2(new_n584), .A3(new_n687), .A4(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n742), .A2(new_n743), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT103), .B1(new_n738), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G36gat), .B1(new_n729), .B2(new_n434), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n751), .A2(new_n752), .A3(new_n746), .A4(new_n748), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(G1329gat));
  NAND2_X1  g553(.A1(new_n705), .A2(G43gat), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n684), .A2(new_n405), .A3(new_n688), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n729), .A2(new_n755), .B1(G43gat), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g557(.A1(new_n728), .A2(new_n300), .A3(new_n687), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT104), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT104), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n728), .A2(new_n761), .A3(new_n300), .A4(new_n687), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(G50gat), .A3(new_n762), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n684), .A2(G50gat), .A3(new_n483), .A4(new_n688), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n759), .A2(G50gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(new_n768), .B2(new_n764), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1331gat));
  NAND3_X1  g569(.A1(new_n620), .A2(new_n686), .A3(new_n662), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT105), .Z(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n717), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n474), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT106), .B(G57gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1332gat));
  AOI21_X1  g575(.A(new_n434), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT107), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n779), .B(new_n780), .Z(G1333gat));
  NAND2_X1  g580(.A1(new_n773), .A2(new_n705), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n405), .A2(G71gat), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n782), .A2(G71gat), .B1(new_n773), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g584(.A1(new_n773), .A2(new_n300), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g586(.A1(new_n685), .A2(new_n643), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n584), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n717), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT51), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n717), .B2(new_n789), .ZN(new_n795));
  INV_X1    g594(.A(new_n789), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n724), .A2(KEYINPUT108), .A3(KEYINPUT51), .A4(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n793), .A2(KEYINPUT109), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT108), .B1(new_n790), .B2(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n795), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n803), .A2(new_n557), .A3(new_n474), .A4(new_n662), .ZN(new_n804));
  INV_X1    g603(.A(new_n788), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n663), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n728), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G85gat), .B1(new_n807), .B2(new_n669), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n808), .ZN(G1336gat));
  INV_X1    g608(.A(new_n806), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n735), .B2(new_n721), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n558), .B1(new_n811), .B2(new_n737), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n434), .A2(G92gat), .A3(new_n663), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n791), .B2(new_n795), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT52), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n800), .A2(new_n801), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n814), .ZN(new_n819));
  OAI21_X1  g618(.A(G92gat), .B1(new_n807), .B2(new_n434), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  OAI211_X1 g620(.A(KEYINPUT110), .B(new_n813), .C1(new_n800), .C2(new_n801), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n816), .A2(new_n823), .ZN(G1337gat));
  NOR3_X1   g623(.A1(new_n405), .A2(G99gat), .A3(new_n663), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n803), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n807), .A2(KEYINPUT111), .A3(new_n491), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT111), .B1(new_n807), .B2(new_n491), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(G99gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n826), .B1(new_n827), .B2(new_n829), .ZN(G1338gat));
  NOR3_X1   g629(.A1(new_n483), .A2(G106gat), .A3(new_n663), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT112), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n791), .B2(new_n795), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n811), .A2(new_n300), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(G106gat), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  INV_X1    g635(.A(G106gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n811), .B2(new_n300), .ZN(new_n838));
  INV_X1    g637(.A(new_n831), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n818), .B2(new_n839), .ZN(new_n840));
  OAI22_X1  g639(.A1(new_n835), .A2(new_n836), .B1(new_n838), .B2(new_n840), .ZN(G1339gat));
  NAND3_X1  g640(.A1(new_n620), .A2(new_n686), .A3(new_n663), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n647), .A2(new_n648), .A3(new_n653), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT113), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n647), .A2(new_n845), .A3(new_n648), .A4(new_n653), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n844), .A2(new_n651), .A3(KEYINPUT54), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n653), .B1(new_n647), .B2(new_n648), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n658), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(KEYINPUT55), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n661), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT55), .B1(new_n847), .B2(new_n850), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n609), .B1(new_n570), .B2(new_n571), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n549), .A2(new_n608), .ZN(new_n856));
  OAI211_X1 g655(.A(G229gat), .B(G233gat), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n632), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n625), .A2(new_n630), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT114), .B1(new_n860), .B2(new_n638), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n862));
  INV_X1    g661(.A(new_n638), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n862), .B(new_n863), .C1(new_n857), .C2(new_n859), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AND4_X1   g664(.A1(new_n642), .A2(new_n584), .A3(new_n854), .A4(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n865), .A2(KEYINPUT115), .A3(new_n642), .A4(new_n662), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n624), .B1(new_n623), .B2(new_n625), .ZN(new_n868));
  INV_X1    g667(.A(new_n859), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n638), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n862), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n860), .A2(KEYINPUT114), .A3(new_n638), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n871), .A2(new_n872), .A3(new_n642), .A4(new_n662), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n643), .A2(new_n854), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n867), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n866), .B1(new_n877), .B2(new_n718), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n842), .B1(new_n878), .B2(new_n685), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n737), .A2(new_n669), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n406), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G113gat), .B1(new_n881), .B2(new_n686), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT116), .Z(new_n883));
  AND2_X1   g682(.A1(new_n879), .A2(new_n474), .ZN(new_n884));
  INV_X1    g683(.A(new_n406), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n737), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n351), .A3(new_n643), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n883), .A2(new_n889), .ZN(G1340gat));
  NOR3_X1   g689(.A1(new_n881), .A2(new_n349), .A3(new_n663), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n662), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n349), .ZN(G1341gat));
  XNOR2_X1  g692(.A(KEYINPUT69), .B(G127gat), .ZN(new_n894));
  INV_X1    g693(.A(new_n685), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n881), .B2(new_n895), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n895), .A2(new_n894), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n887), .B2(new_n897), .ZN(G1342gat));
  NAND3_X1  g697(.A1(new_n888), .A2(new_n355), .A3(new_n584), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT56), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT117), .ZN(new_n901));
  OAI21_X1  g700(.A(G134gat), .B1(new_n881), .B2(new_n718), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n901), .B(new_n902), .C1(KEYINPUT56), .C2(new_n899), .ZN(G1343gat));
  NAND2_X1  g702(.A1(new_n880), .A2(new_n491), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n852), .B2(new_n853), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n847), .A2(new_n850), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT55), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n911), .A2(KEYINPUT119), .A3(new_n661), .A4(new_n851), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n908), .A2(new_n643), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n873), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(KEYINPUT120), .A3(new_n873), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n916), .A2(new_n718), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n895), .B1(new_n918), .B2(new_n866), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n483), .B1(new_n919), .B2(new_n842), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n906), .B1(new_n920), .B2(KEYINPUT57), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n584), .B1(new_n914), .B2(new_n915), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n866), .B1(new_n922), .B2(new_n917), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n842), .B1(new_n923), .B2(new_n685), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n924), .A2(new_n906), .A3(KEYINPUT57), .A4(new_n300), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n879), .A2(new_n300), .ZN(new_n926));
  XOR2_X1   g725(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n643), .B(new_n905), .C1(new_n921), .C2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n264), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND4_X1   g731(.A1(new_n300), .A2(new_n884), .A3(new_n434), .A4(new_n491), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n229), .A3(new_n643), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT58), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT58), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n932), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1344gat));
  NAND3_X1  g738(.A1(new_n933), .A2(new_n234), .A3(new_n662), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n905), .A2(new_n662), .ZN(new_n942));
  INV_X1    g741(.A(new_n927), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n879), .A2(new_n300), .A3(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n924), .A2(new_n300), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT57), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n942), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n234), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n944), .B(KEYINPUT122), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n920), .A2(KEYINPUT57), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT123), .B1(new_n955), .B2(new_n942), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n941), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n941), .A2(G148gat), .ZN(new_n958));
  INV_X1    g757(.A(new_n921), .ZN(new_n959));
  INV_X1    g758(.A(new_n929), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n904), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n958), .B1(new_n961), .B2(new_n662), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n940), .B1(new_n957), .B2(new_n962), .ZN(G1345gat));
  NAND3_X1  g762(.A1(new_n933), .A2(new_n613), .A3(new_n685), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n961), .A2(new_n685), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n613), .ZN(G1346gat));
  INV_X1    g765(.A(G162gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n933), .A2(new_n967), .A3(new_n584), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n584), .B(new_n905), .C1(new_n921), .C2(new_n929), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT124), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(G162gat), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n969), .A2(KEYINPUT124), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1347gat));
  AND4_X1   g772(.A1(new_n669), .A2(new_n879), .A3(new_n737), .A4(new_n406), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n643), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n662), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g777(.A1(new_n974), .A2(new_n685), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n980));
  AOI22_X1  g779(.A1(new_n979), .A2(G183gat), .B1(new_n980), .B2(KEYINPUT60), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n981), .B1(new_n363), .B2(new_n979), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n980), .A2(KEYINPUT60), .ZN(new_n983));
  XOR2_X1   g782(.A(new_n982), .B(new_n983), .Z(G1350gat));
  AOI21_X1  g783(.A(new_n313), .B1(new_n974), .B2(new_n584), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n985), .A2(KEYINPUT126), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(KEYINPUT126), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n986), .A2(KEYINPUT61), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n974), .A2(new_n313), .A3(new_n584), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n988), .B(new_n989), .C1(KEYINPUT61), .C2(new_n986), .ZN(G1351gat));
  NOR3_X1   g789(.A1(new_n705), .A2(new_n474), .A3(new_n434), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n879), .A2(new_n300), .A3(new_n991), .ZN(new_n992));
  XOR2_X1   g791(.A(new_n992), .B(KEYINPUT127), .Z(new_n993));
  AOI21_X1  g792(.A(G197gat), .B1(new_n993), .B2(new_n643), .ZN(new_n994));
  INV_X1    g793(.A(new_n955), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(new_n991), .ZN(new_n996));
  INV_X1    g795(.A(new_n996), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n643), .A2(G197gat), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(G1352gat));
  OAI21_X1  g798(.A(G204gat), .B1(new_n996), .B2(new_n663), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n992), .A2(G204gat), .A3(new_n663), .ZN(new_n1001));
  XNOR2_X1  g800(.A(new_n1001), .B(KEYINPUT62), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1000), .A2(new_n1002), .ZN(G1353gat));
  NAND3_X1  g802(.A1(new_n993), .A2(new_n215), .A3(new_n685), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n685), .B(new_n991), .C1(new_n953), .C2(new_n954), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1005), .B2(G211gat), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(G1354gat));
  OAI21_X1  g807(.A(G218gat), .B1(new_n996), .B2(new_n718), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n993), .A2(new_n216), .A3(new_n584), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(G1355gat));
endmodule


