

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(n752), .A2(n751), .ZN(n753) );
  INV_X1 U554 ( .A(n734), .ZN(n718) );
  NOR2_X2 U555 ( .A1(n700), .A2(n966), .ZN(n706) );
  XOR2_X1 U556 ( .A(KEYINPUT32), .B(n741), .Z(n517) );
  NOR2_X1 U557 ( .A1(n517), .A2(n747), .ZN(n768) );
  INV_X1 U558 ( .A(KEYINPUT88), .ZN(n674) );
  XNOR2_X1 U559 ( .A(n675), .B(n674), .ZN(n688) );
  NOR2_X2 U560 ( .A1(G2104), .A2(n519), .ZN(n870) );
  AND2_X1 U561 ( .A1(n519), .A2(G2104), .ZN(n873) );
  NOR2_X1 U562 ( .A1(G651), .A2(n613), .ZN(n636) );
  XNOR2_X1 U563 ( .A(n521), .B(n520), .ZN(n522) );
  INV_X1 U564 ( .A(G2105), .ZN(n519) );
  NAND2_X1 U565 ( .A1(G125), .A2(n870), .ZN(n518) );
  XOR2_X1 U566 ( .A(KEYINPUT65), .B(n518), .Z(n523) );
  NAND2_X1 U567 ( .A1(G101), .A2(n873), .ZN(n521) );
  XOR2_X1 U568 ( .A(KEYINPUT23), .B(KEYINPUT66), .Z(n520) );
  NAND2_X1 U569 ( .A1(n523), .A2(n522), .ZN(n529) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n871) );
  NAND2_X1 U571 ( .A1(n871), .A2(G113), .ZN(n527) );
  XNOR2_X1 U572 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n525) );
  NOR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XNOR2_X1 U574 ( .A(n525), .B(n524), .ZN(n874) );
  NAND2_X1 U575 ( .A1(n874), .A2(G137), .ZN(n526) );
  NAND2_X1 U576 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U577 ( .A1(n529), .A2(n528), .ZN(G160) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n632) );
  NAND2_X1 U579 ( .A1(G89), .A2(n632), .ZN(n530) );
  XNOR2_X1 U580 ( .A(n530), .B(KEYINPUT4), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n531), .B(KEYINPUT76), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n613) );
  INV_X1 U583 ( .A(G651), .ZN(n535) );
  NOR2_X1 U584 ( .A1(n613), .A2(n535), .ZN(n633) );
  NAND2_X1 U585 ( .A1(G76), .A2(n633), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U587 ( .A(n534), .B(KEYINPUT5), .ZN(n541) );
  NOR2_X1 U588 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n536), .Z(n631) );
  NAND2_X1 U590 ( .A1(G63), .A2(n631), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G51), .A2(n636), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT6), .B(n539), .Z(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U595 ( .A(n542), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U596 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U597 ( .A1(G85), .A2(n632), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G72), .A2(n633), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G60), .A2(n631), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G47), .A2(n636), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U603 ( .A1(n548), .A2(n547), .ZN(G290) );
  AND2_X1 U604 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U605 ( .A(G108), .ZN(G238) );
  INV_X1 U606 ( .A(G82), .ZN(G220) );
  NAND2_X1 U607 ( .A1(n632), .A2(G90), .ZN(n549) );
  XOR2_X1 U608 ( .A(KEYINPUT69), .B(n549), .Z(n551) );
  NAND2_X1 U609 ( .A1(n633), .A2(G77), .ZN(n550) );
  NAND2_X1 U610 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n552), .B(KEYINPUT9), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G64), .A2(n631), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n636), .A2(G52), .ZN(n555) );
  XOR2_X1 U615 ( .A(KEYINPUT68), .B(n555), .Z(n556) );
  NOR2_X1 U616 ( .A1(n557), .A2(n556), .ZN(G171) );
  INV_X1 U617 ( .A(G171), .ZN(G301) );
  NAND2_X1 U618 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U619 ( .A(n558), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U620 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n560) );
  INV_X1 U621 ( .A(G223), .ZN(n817) );
  NAND2_X1 U622 ( .A1(G567), .A2(n817), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n560), .B(n559), .ZN(G234) );
  NAND2_X1 U624 ( .A1(G56), .A2(n631), .ZN(n561) );
  XOR2_X1 U625 ( .A(KEYINPUT14), .B(n561), .Z(n567) );
  NAND2_X1 U626 ( .A1(n632), .A2(G81), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G68), .A2(n633), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT13), .B(n565), .Z(n566) );
  NOR2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n636), .A2(G43), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n966) );
  INV_X1 U634 ( .A(G860), .ZN(n591) );
  OR2_X1 U635 ( .A1(n966), .A2(n591), .ZN(G153) );
  NAND2_X1 U636 ( .A1(G868), .A2(G301), .ZN(n581) );
  NAND2_X1 U637 ( .A1(G92), .A2(n632), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n570), .B(KEYINPUT74), .ZN(n577) );
  NAND2_X1 U639 ( .A1(G79), .A2(n633), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G54), .A2(n636), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G66), .A2(n631), .ZN(n573) );
  XNOR2_X1 U643 ( .A(KEYINPUT73), .B(n573), .ZN(n574) );
  NOR2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT75), .B(KEYINPUT15), .Z(n578) );
  XNOR2_X1 U647 ( .A(n579), .B(n578), .ZN(n707) );
  INV_X1 U648 ( .A(n707), .ZN(n974) );
  INV_X1 U649 ( .A(G868), .ZN(n651) );
  NAND2_X1 U650 ( .A1(n974), .A2(n651), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U652 ( .A1(G91), .A2(n632), .ZN(n583) );
  NAND2_X1 U653 ( .A1(G78), .A2(n633), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n631), .A2(G65), .ZN(n584) );
  XOR2_X1 U656 ( .A(KEYINPUT70), .B(n584), .Z(n585) );
  NOR2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n636), .A2(G53), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(G299) );
  NOR2_X1 U660 ( .A1(G286), .A2(n651), .ZN(n590) );
  NOR2_X1 U661 ( .A1(G868), .A2(G299), .ZN(n589) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(G297) );
  NAND2_X1 U663 ( .A1(n591), .A2(G559), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n592), .A2(n707), .ZN(n593) );
  XNOR2_X1 U665 ( .A(n593), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U666 ( .A1(G868), .A2(n966), .ZN(n596) );
  NAND2_X1 U667 ( .A1(G868), .A2(n707), .ZN(n594) );
  NOR2_X1 U668 ( .A1(G559), .A2(n594), .ZN(n595) );
  NOR2_X1 U669 ( .A1(n596), .A2(n595), .ZN(G282) );
  NAND2_X1 U670 ( .A1(G135), .A2(n874), .ZN(n605) );
  NAND2_X1 U671 ( .A1(G123), .A2(n870), .ZN(n597) );
  XNOR2_X1 U672 ( .A(n597), .B(KEYINPUT18), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G99), .A2(n873), .ZN(n598) );
  XNOR2_X1 U674 ( .A(n598), .B(KEYINPUT78), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G111), .A2(n871), .ZN(n601) );
  XNOR2_X1 U677 ( .A(KEYINPUT77), .B(n601), .ZN(n602) );
  NOR2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n606), .B(KEYINPUT79), .ZN(n922) );
  XNOR2_X1 U681 ( .A(n922), .B(G2096), .ZN(n608) );
  INV_X1 U682 ( .A(G2100), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(G156) );
  NAND2_X1 U684 ( .A1(G49), .A2(n636), .ZN(n610) );
  NAND2_X1 U685 ( .A1(G74), .A2(G651), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U687 ( .A1(n631), .A2(n611), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n612), .B(KEYINPUT82), .ZN(n615) );
  NAND2_X1 U689 ( .A1(G87), .A2(n613), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(G288) );
  NAND2_X1 U691 ( .A1(G62), .A2(n631), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G50), .A2(n636), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U694 ( .A(KEYINPUT83), .B(n618), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G88), .A2(n632), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G75), .A2(n633), .ZN(n619) );
  AND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(G303) );
  INV_X1 U699 ( .A(G303), .ZN(G166) );
  NAND2_X1 U700 ( .A1(G61), .A2(n631), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G86), .A2(n632), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n633), .A2(G73), .ZN(n625) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(n625), .Z(n626) );
  NOR2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n636), .A2(G48), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(G305) );
  NAND2_X1 U708 ( .A1(G559), .A2(n707), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n630), .B(n966), .ZN(n825) );
  NAND2_X1 U710 ( .A1(n631), .A2(G67), .ZN(n641) );
  NAND2_X1 U711 ( .A1(G93), .A2(n632), .ZN(n635) );
  NAND2_X1 U712 ( .A1(G80), .A2(n633), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n636), .A2(G55), .ZN(n637) );
  XOR2_X1 U715 ( .A(KEYINPUT80), .B(n637), .Z(n638) );
  NOR2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U718 ( .A(KEYINPUT81), .B(n642), .Z(n826) );
  XNOR2_X1 U719 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n644) );
  XNOR2_X1 U720 ( .A(G288), .B(KEYINPUT85), .ZN(n643) );
  XNOR2_X1 U721 ( .A(n644), .B(n643), .ZN(n645) );
  XOR2_X1 U722 ( .A(n826), .B(n645), .Z(n647) );
  XNOR2_X1 U723 ( .A(G290), .B(G166), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U725 ( .A(n648), .B(G299), .ZN(n649) );
  XNOR2_X1 U726 ( .A(n649), .B(G305), .ZN(n891) );
  XNOR2_X1 U727 ( .A(n825), .B(n891), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n650), .A2(G868), .ZN(n653) );
  NAND2_X1 U729 ( .A1(n651), .A2(n826), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(G295) );
  NAND2_X1 U731 ( .A1(G2078), .A2(G2084), .ZN(n654) );
  XOR2_X1 U732 ( .A(KEYINPUT20), .B(n654), .Z(n655) );
  NAND2_X1 U733 ( .A1(G2090), .A2(n655), .ZN(n656) );
  XNOR2_X1 U734 ( .A(KEYINPUT21), .B(n656), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n657), .A2(G2072), .ZN(n658) );
  XNOR2_X1 U736 ( .A(KEYINPUT86), .B(n658), .ZN(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U738 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NOR2_X1 U739 ( .A1(G220), .A2(G219), .ZN(n659) );
  XOR2_X1 U740 ( .A(KEYINPUT22), .B(n659), .Z(n660) );
  NOR2_X1 U741 ( .A1(G218), .A2(n660), .ZN(n661) );
  NAND2_X1 U742 ( .A1(G96), .A2(n661), .ZN(n823) );
  NAND2_X1 U743 ( .A1(n823), .A2(G2106), .ZN(n665) );
  NAND2_X1 U744 ( .A1(G120), .A2(G69), .ZN(n662) );
  NOR2_X1 U745 ( .A1(G238), .A2(n662), .ZN(n663) );
  NAND2_X1 U746 ( .A1(G57), .A2(n663), .ZN(n824) );
  NAND2_X1 U747 ( .A1(n824), .A2(G567), .ZN(n664) );
  NAND2_X1 U748 ( .A1(n665), .A2(n664), .ZN(n828) );
  NAND2_X1 U749 ( .A1(G483), .A2(G661), .ZN(n666) );
  NOR2_X1 U750 ( .A1(n828), .A2(n666), .ZN(n822) );
  NAND2_X1 U751 ( .A1(n822), .A2(G36), .ZN(G176) );
  NAND2_X1 U752 ( .A1(G102), .A2(n873), .ZN(n668) );
  NAND2_X1 U753 ( .A1(G138), .A2(n874), .ZN(n667) );
  NAND2_X1 U754 ( .A1(n668), .A2(n667), .ZN(n673) );
  NAND2_X1 U755 ( .A1(G126), .A2(n870), .ZN(n670) );
  NAND2_X1 U756 ( .A1(G114), .A2(n871), .ZN(n669) );
  NAND2_X1 U757 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U758 ( .A(KEYINPUT87), .B(n671), .Z(n672) );
  NOR2_X1 U759 ( .A1(n673), .A2(n672), .ZN(G164) );
  XNOR2_X1 U760 ( .A(G1986), .B(G290), .ZN(n971) );
  NAND2_X1 U761 ( .A1(G160), .A2(G40), .ZN(n675) );
  INV_X1 U762 ( .A(n688), .ZN(n676) );
  NOR2_X1 U763 ( .A1(G164), .A2(G1384), .ZN(n689) );
  NOR2_X1 U764 ( .A1(n676), .A2(n689), .ZN(n812) );
  NAND2_X1 U765 ( .A1(n971), .A2(n812), .ZN(n800) );
  NAND2_X1 U766 ( .A1(G104), .A2(n873), .ZN(n678) );
  NAND2_X1 U767 ( .A1(G140), .A2(n874), .ZN(n677) );
  NAND2_X1 U768 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U769 ( .A(KEYINPUT34), .B(n679), .ZN(n685) );
  NAND2_X1 U770 ( .A1(G128), .A2(n870), .ZN(n681) );
  NAND2_X1 U771 ( .A1(G116), .A2(n871), .ZN(n680) );
  NAND2_X1 U772 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U773 ( .A(KEYINPUT89), .B(n682), .ZN(n683) );
  XNOR2_X1 U774 ( .A(KEYINPUT35), .B(n683), .ZN(n684) );
  NOR2_X1 U775 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U776 ( .A(KEYINPUT36), .B(n686), .ZN(n888) );
  XNOR2_X1 U777 ( .A(KEYINPUT37), .B(G2067), .ZN(n810) );
  NOR2_X1 U778 ( .A1(n888), .A2(n810), .ZN(n913) );
  NAND2_X1 U779 ( .A1(n812), .A2(n913), .ZN(n687) );
  XNOR2_X1 U780 ( .A(KEYINPUT90), .B(n687), .ZN(n808) );
  INV_X1 U781 ( .A(n808), .ZN(n798) );
  INV_X1 U782 ( .A(G299), .ZN(n711) );
  NAND2_X2 U783 ( .A1(n689), .A2(n688), .ZN(n734) );
  XNOR2_X1 U784 ( .A(G1956), .B(KEYINPUT98), .ZN(n998) );
  NAND2_X1 U785 ( .A1(n734), .A2(n998), .ZN(n690) );
  XNOR2_X1 U786 ( .A(KEYINPUT99), .B(n690), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n718), .A2(G2072), .ZN(n691) );
  XNOR2_X1 U788 ( .A(KEYINPUT27), .B(n691), .ZN(n692) );
  NOR2_X1 U789 ( .A1(n693), .A2(n692), .ZN(n710) );
  NOR2_X1 U790 ( .A1(n711), .A2(n710), .ZN(n694) );
  XOR2_X1 U791 ( .A(n694), .B(KEYINPUT28), .Z(n715) );
  AND2_X1 U792 ( .A1(n718), .A2(G1996), .ZN(n697) );
  XOR2_X1 U793 ( .A(KEYINPUT26), .B(KEYINPUT100), .Z(n695) );
  XNOR2_X1 U794 ( .A(KEYINPUT64), .B(n695), .ZN(n696) );
  XNOR2_X1 U795 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U796 ( .A1(n734), .A2(G1341), .ZN(n698) );
  NAND2_X1 U797 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U798 ( .A1(n706), .A2(n707), .ZN(n705) );
  AND2_X1 U799 ( .A1(n718), .A2(G2067), .ZN(n701) );
  XNOR2_X1 U800 ( .A(n701), .B(KEYINPUT101), .ZN(n703) );
  NAND2_X1 U801 ( .A1(n734), .A2(G1348), .ZN(n702) );
  NAND2_X1 U802 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U803 ( .A1(n705), .A2(n704), .ZN(n709) );
  OR2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n717) );
  XOR2_X1 U809 ( .A(KEYINPUT102), .B(KEYINPUT29), .Z(n716) );
  XNOR2_X1 U810 ( .A(n717), .B(n716), .ZN(n723) );
  NAND2_X1 U811 ( .A1(G1961), .A2(n734), .ZN(n720) );
  XOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .Z(n944) );
  NAND2_X1 U813 ( .A1(n718), .A2(n944), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n724) );
  NOR2_X1 U815 ( .A1(G301), .A2(n724), .ZN(n721) );
  XNOR2_X1 U816 ( .A(KEYINPUT97), .B(n721), .ZN(n722) );
  NAND2_X1 U817 ( .A1(n723), .A2(n722), .ZN(n733) );
  NAND2_X1 U818 ( .A1(G301), .A2(n724), .ZN(n725) );
  XNOR2_X1 U819 ( .A(n725), .B(KEYINPUT103), .ZN(n730) );
  NAND2_X1 U820 ( .A1(G8), .A2(n734), .ZN(n765) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n765), .ZN(n746) );
  NOR2_X1 U822 ( .A1(G2084), .A2(n734), .ZN(n742) );
  NOR2_X1 U823 ( .A1(n746), .A2(n742), .ZN(n726) );
  NAND2_X1 U824 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U825 ( .A(KEYINPUT30), .B(n727), .ZN(n728) );
  NOR2_X1 U826 ( .A1(n728), .A2(G168), .ZN(n729) );
  NOR2_X1 U827 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U828 ( .A(KEYINPUT31), .B(n731), .Z(n732) );
  NAND2_X1 U829 ( .A1(n733), .A2(n732), .ZN(n744) );
  NAND2_X1 U830 ( .A1(n744), .A2(G286), .ZN(n739) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n765), .ZN(n736) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n734), .ZN(n735) );
  NOR2_X1 U833 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U834 ( .A1(n737), .A2(G303), .ZN(n738) );
  NAND2_X1 U835 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U836 ( .A1(G8), .A2(n740), .ZN(n741) );
  NAND2_X1 U837 ( .A1(G8), .A2(n742), .ZN(n743) );
  NAND2_X1 U838 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U842 ( .A1(n756), .A2(n748), .ZN(n973) );
  XOR2_X1 U843 ( .A(n973), .B(KEYINPUT104), .Z(n749) );
  NOR2_X1 U844 ( .A1(n768), .A2(n749), .ZN(n752) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n965) );
  NOR2_X1 U846 ( .A1(KEYINPUT105), .A2(n765), .ZN(n750) );
  NAND2_X1 U847 ( .A1(n965), .A2(n750), .ZN(n751) );
  NOR2_X1 U848 ( .A1(KEYINPUT33), .A2(n753), .ZN(n761) );
  INV_X1 U849 ( .A(KEYINPUT105), .ZN(n755) );
  NAND2_X1 U850 ( .A1(n756), .A2(KEYINPUT33), .ZN(n754) );
  NAND2_X1 U851 ( .A1(n755), .A2(n754), .ZN(n758) );
  NAND2_X1 U852 ( .A1(n756), .A2(KEYINPUT105), .ZN(n757) );
  NAND2_X1 U853 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U854 ( .A1(n765), .A2(n759), .ZN(n760) );
  NOR2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U856 ( .A(G1981), .B(G305), .Z(n961) );
  NAND2_X1 U857 ( .A1(n762), .A2(n961), .ZN(n774) );
  NOR2_X1 U858 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XOR2_X1 U859 ( .A(n763), .B(KEYINPUT24), .Z(n764) );
  NOR2_X1 U860 ( .A1(n765), .A2(n764), .ZN(n772) );
  INV_X1 U861 ( .A(n765), .ZN(n770) );
  NAND2_X1 U862 ( .A1(G166), .A2(G8), .ZN(n766) );
  NOR2_X1 U863 ( .A1(G2090), .A2(n766), .ZN(n767) );
  NOR2_X1 U864 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U865 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U866 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n796) );
  NAND2_X1 U868 ( .A1(G95), .A2(n873), .ZN(n776) );
  NAND2_X1 U869 ( .A1(G131), .A2(n874), .ZN(n775) );
  NAND2_X1 U870 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U871 ( .A1(G119), .A2(n870), .ZN(n777) );
  XNOR2_X1 U872 ( .A(KEYINPUT91), .B(n777), .ZN(n778) );
  NOR2_X1 U873 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n871), .A2(G107), .ZN(n780) );
  NAND2_X1 U875 ( .A1(n781), .A2(n780), .ZN(n858) );
  NAND2_X1 U876 ( .A1(G1991), .A2(n858), .ZN(n782) );
  XNOR2_X1 U877 ( .A(KEYINPUT92), .B(n782), .ZN(n794) );
  NAND2_X1 U878 ( .A1(n871), .A2(G117), .ZN(n783) );
  XOR2_X1 U879 ( .A(KEYINPUT93), .B(n783), .Z(n785) );
  NAND2_X1 U880 ( .A1(n870), .A2(G129), .ZN(n784) );
  NAND2_X1 U881 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U882 ( .A(KEYINPUT94), .B(n786), .ZN(n789) );
  NAND2_X1 U883 ( .A1(n873), .A2(G105), .ZN(n787) );
  XOR2_X1 U884 ( .A(KEYINPUT38), .B(n787), .Z(n788) );
  NOR2_X1 U885 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n874), .A2(G141), .ZN(n790) );
  NAND2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n885) );
  NAND2_X1 U888 ( .A1(G1996), .A2(n885), .ZN(n792) );
  XOR2_X1 U889 ( .A(KEYINPUT95), .B(n792), .Z(n793) );
  NAND2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U891 ( .A(KEYINPUT96), .B(n795), .ZN(n935) );
  NAND2_X1 U892 ( .A1(n812), .A2(n935), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n796), .A2(n803), .ZN(n797) );
  NOR2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U895 ( .A1(n800), .A2(n799), .ZN(n815) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n885), .ZN(n927) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n801) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n858), .ZN(n923) );
  NOR2_X1 U899 ( .A1(n801), .A2(n923), .ZN(n802) );
  XOR2_X1 U900 ( .A(KEYINPUT106), .B(n802), .Z(n804) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U902 ( .A(KEYINPUT107), .B(n805), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n927), .A2(n806), .ZN(n807) );
  XNOR2_X1 U904 ( .A(n807), .B(KEYINPUT39), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n888), .A2(n810), .ZN(n912) );
  NAND2_X1 U907 ( .A1(n811), .A2(n912), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n816), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n817), .ZN(G217) );
  NAND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n818) );
  XNOR2_X1 U913 ( .A(KEYINPUT109), .B(n818), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n819), .A2(G661), .ZN(n820) );
  XNOR2_X1 U915 ( .A(KEYINPUT110), .B(n820), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(G188) );
  XNOR2_X1 U918 ( .A(G120), .B(KEYINPUT111), .ZN(G236) );
  XOR2_X1 U919 ( .A(G69), .B(KEYINPUT112), .Z(G235) );
  INV_X1 U921 ( .A(G96), .ZN(G221) );
  NOR2_X1 U922 ( .A1(n824), .A2(n823), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  NOR2_X1 U924 ( .A1(n825), .A2(G860), .ZN(n827) );
  XOR2_X1 U925 ( .A(n827), .B(n826), .Z(G145) );
  INV_X1 U926 ( .A(n828), .ZN(G319) );
  XOR2_X1 U927 ( .A(KEYINPUT114), .B(KEYINPUT43), .Z(n830) );
  XNOR2_X1 U928 ( .A(KEYINPUT113), .B(G2678), .ZN(n829) );
  XNOR2_X1 U929 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U930 ( .A(KEYINPUT42), .B(G2090), .Z(n832) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2072), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U933 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U934 ( .A(G2096), .B(G2100), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n838) );
  XOR2_X1 U936 ( .A(G2078), .B(G2084), .Z(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U938 ( .A(G1961), .B(G1956), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1966), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U941 ( .A(n841), .B(G2474), .Z(n843) );
  XNOR2_X1 U942 ( .A(G1971), .B(G1976), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U944 ( .A(KEYINPUT41), .B(G1981), .Z(n845) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U948 ( .A1(G100), .A2(n873), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n848), .B(KEYINPUT116), .ZN(n852) );
  XOR2_X1 U950 ( .A(KEYINPUT115), .B(KEYINPUT44), .Z(n850) );
  NAND2_X1 U951 ( .A1(G124), .A2(n870), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n851) );
  NAND2_X1 U953 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U954 ( .A1(G136), .A2(n874), .ZN(n854) );
  NAND2_X1 U955 ( .A1(G112), .A2(n871), .ZN(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U957 ( .A1(n856), .A2(n855), .ZN(G162) );
  XOR2_X1 U958 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n869) );
  NAND2_X1 U960 ( .A1(G103), .A2(n873), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G139), .A2(n874), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G127), .A2(n870), .ZN(n862) );
  NAND2_X1 U964 ( .A1(G115), .A2(n871), .ZN(n861) );
  NAND2_X1 U965 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U966 ( .A(KEYINPUT47), .B(n863), .Z(n864) );
  NOR2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n915) );
  XOR2_X1 U968 ( .A(n915), .B(G162), .Z(n867) );
  XNOR2_X1 U969 ( .A(G160), .B(G164), .ZN(n866) );
  XNOR2_X1 U970 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n887) );
  NAND2_X1 U972 ( .A1(G130), .A2(n870), .ZN(n882) );
  NAND2_X1 U973 ( .A1(n871), .A2(G118), .ZN(n872) );
  XNOR2_X1 U974 ( .A(KEYINPUT117), .B(n872), .ZN(n880) );
  NAND2_X1 U975 ( .A1(G106), .A2(n873), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G142), .A2(n874), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(KEYINPUT118), .B(n877), .Z(n878) );
  XNOR2_X1 U979 ( .A(KEYINPUT45), .B(n878), .ZN(n879) );
  NOR2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n883), .B(n922), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n889) );
  XOR2_X1 U985 ( .A(n889), .B(n888), .Z(n890) );
  NOR2_X1 U986 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U987 ( .A(G286), .B(n891), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n966), .B(G171), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n894), .B(n974), .ZN(n895) );
  NOR2_X1 U991 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U992 ( .A(G2438), .B(G2435), .Z(n897) );
  XNOR2_X1 U993 ( .A(G2443), .B(G2430), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(n898), .B(G2454), .Z(n900) );
  XNOR2_X1 U996 ( .A(G1341), .B(G1348), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U998 ( .A(G2451), .B(G2427), .Z(n902) );
  XNOR2_X1 U999 ( .A(KEYINPUT108), .B(G2446), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(n904), .B(n903), .Z(n905) );
  NAND2_X1 U1002 ( .A1(G14), .A2(n905), .ZN(n911) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G57), .ZN(G237) );
  INV_X1 U1011 ( .A(n911), .ZN(G401) );
  INV_X1 U1012 ( .A(KEYINPUT55), .ZN(n957) );
  INV_X1 U1013 ( .A(n912), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n933) );
  XNOR2_X1 U1015 ( .A(G164), .B(G2078), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(G2072), .B(n915), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(KEYINPUT120), .ZN(n917) );
  NAND2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n919), .B(KEYINPUT50), .ZN(n921) );
  XOR2_X1 U1020 ( .A(G2084), .B(G160), .Z(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n925) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n931) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n928), .Z(n929) );
  XNOR2_X1 U1027 ( .A(n929), .B(KEYINPUT119), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n936), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n957), .A2(n937), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n938), .A2(G29), .ZN(n990) );
  XNOR2_X1 U1034 ( .A(KEYINPUT121), .B(G2090), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(n939), .B(G35), .ZN(n955) );
  XNOR2_X1 U1036 ( .A(G2084), .B(G34), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(n940), .B(KEYINPUT54), .ZN(n953) );
  XOR2_X1 U1038 ( .A(G1991), .B(G25), .Z(n941) );
  NAND2_X1 U1039 ( .A1(n941), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(G1996), .B(G32), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(G27), .B(n944), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(n951), .B(KEYINPUT53), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n957), .B(n956), .ZN(n959) );
  INV_X1 U1052 ( .A(G29), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(G11), .A2(n960), .ZN(n988) );
  XNOR2_X1 U1055 ( .A(G1966), .B(G168), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1057 ( .A(KEYINPUT57), .B(n963), .Z(n983) );
  NAND2_X1 U1058 ( .A1(G1971), .A2(G303), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n980) );
  XNOR2_X1 U1060 ( .A(n966), .B(G1341), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(G301), .B(G1961), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n978) );
  XNOR2_X1 U1063 ( .A(G1956), .B(KEYINPUT122), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n969), .B(G299), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(G1348), .B(n974), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(n981), .B(KEYINPUT123), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n985) );
  XOR2_X1 U1073 ( .A(G16), .B(KEYINPUT56), .Z(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(n986), .B(KEYINPUT124), .ZN(n987) );
  NOR2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n1017) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G22), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(G23), .B(G1976), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1081 ( .A(KEYINPUT126), .B(n993), .Z(n995) );
  XNOR2_X1 U1082 ( .A(G1986), .B(G24), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1084 ( .A(KEYINPUT58), .B(n996), .Z(n1012) );
  XOR2_X1 U1085 ( .A(G1961), .B(G5), .Z(n1007) );
  XNOR2_X1 U1086 ( .A(G1348), .B(KEYINPUT59), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(G4), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(n998), .B(G20), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(G19), .B(G1341), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G6), .B(G1981), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G21), .B(G1966), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT125), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(n1013), .B(KEYINPUT127), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(G16), .A2(n1015), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(n1018), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

