

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U556 ( .A(KEYINPUT99), .B(n750), .Z(n522) );
  OR2_X1 U557 ( .A1(n966), .A2(n705), .ZN(n717) );
  NOR2_X1 U558 ( .A1(G1384), .A2(G164), .ZN(n681) );
  XNOR2_X1 U559 ( .A(n744), .B(KEYINPUT32), .ZN(n745) );
  XNOR2_X1 U560 ( .A(n746), .B(n745), .ZN(n747) );
  XOR2_X1 U561 ( .A(KEYINPUT17), .B(n523), .Z(n887) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  NAND2_X1 U563 ( .A1(n887), .A2(G138), .ZN(n526) );
  INV_X1 U564 ( .A(G2105), .ZN(n527) );
  AND2_X1 U565 ( .A1(n527), .A2(G2104), .ZN(n888) );
  NAND2_X1 U566 ( .A1(G102), .A2(n888), .ZN(n524) );
  XOR2_X1 U567 ( .A(KEYINPUT83), .B(n524), .Z(n525) );
  NAND2_X1 U568 ( .A1(n526), .A2(n525), .ZN(n531) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n891) );
  NAND2_X1 U570 ( .A1(G114), .A2(n891), .ZN(n529) );
  NOR2_X1 U571 ( .A1(G2104), .A2(n527), .ZN(n892) );
  NAND2_X1 U572 ( .A1(G126), .A2(n892), .ZN(n528) );
  NAND2_X1 U573 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U574 ( .A1(n531), .A2(n530), .ZN(G164) );
  NOR2_X1 U575 ( .A1(G651), .A2(G543), .ZN(n532) );
  XOR2_X1 U576 ( .A(KEYINPUT65), .B(n532), .Z(n638) );
  NAND2_X1 U577 ( .A1(G85), .A2(n638), .ZN(n535) );
  INV_X1 U578 ( .A(G651), .ZN(n536) );
  NOR2_X1 U579 ( .A1(G543), .A2(n536), .ZN(n533) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n533), .Z(n634) );
  NAND2_X1 U581 ( .A1(G60), .A2(n634), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n535), .A2(n534), .ZN(n541) );
  XOR2_X1 U583 ( .A(KEYINPUT0), .B(G543), .Z(n618) );
  NOR2_X1 U584 ( .A1(n618), .A2(n536), .ZN(n631) );
  NAND2_X1 U585 ( .A1(G72), .A2(n631), .ZN(n539) );
  NOR2_X1 U586 ( .A1(G651), .A2(n618), .ZN(n537) );
  XNOR2_X1 U587 ( .A(KEYINPUT66), .B(n537), .ZN(n635) );
  NAND2_X1 U588 ( .A1(G47), .A2(n635), .ZN(n538) );
  NAND2_X1 U589 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U590 ( .A1(n541), .A2(n540), .ZN(G290) );
  AND2_X1 U591 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U592 ( .A(G57), .ZN(G237) );
  INV_X1 U593 ( .A(G132), .ZN(G219) );
  INV_X1 U594 ( .A(G82), .ZN(G220) );
  NAND2_X1 U595 ( .A1(G7), .A2(G661), .ZN(n542) );
  XNOR2_X1 U596 ( .A(n542), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U597 ( .A(G223), .ZN(n834) );
  NAND2_X1 U598 ( .A1(n834), .A2(G567), .ZN(n543) );
  XOR2_X1 U599 ( .A(KEYINPUT11), .B(n543), .Z(G234) );
  XOR2_X1 U600 ( .A(KEYINPUT14), .B(KEYINPUT68), .Z(n545) );
  NAND2_X1 U601 ( .A1(G56), .A2(n634), .ZN(n544) );
  XNOR2_X1 U602 ( .A(n545), .B(n544), .ZN(n554) );
  NAND2_X1 U603 ( .A1(n638), .A2(G81), .ZN(n546) );
  XNOR2_X1 U604 ( .A(KEYINPUT12), .B(n546), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n631), .A2(G68), .ZN(n547) );
  XOR2_X1 U606 ( .A(KEYINPUT69), .B(n547), .Z(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U608 ( .A(n550), .B(KEYINPUT13), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G43), .A2(n635), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n982) );
  NAND2_X1 U612 ( .A1(n982), .A2(G860), .ZN(G153) );
  NAND2_X1 U613 ( .A1(G64), .A2(n634), .ZN(n555) );
  XNOR2_X1 U614 ( .A(n555), .B(KEYINPUT67), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G90), .A2(n638), .ZN(n557) );
  NAND2_X1 U616 ( .A1(G77), .A2(n631), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U620 ( .A1(G52), .A2(n635), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(G301) );
  NAND2_X1 U622 ( .A1(G868), .A2(G301), .ZN(n571) );
  NAND2_X1 U623 ( .A1(G92), .A2(n638), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G66), .A2(n634), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G79), .A2(n631), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G54), .A2(n635), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT15), .B(n569), .Z(n966) );
  INV_X1 U631 ( .A(n966), .ZN(n845) );
  INV_X1 U632 ( .A(G868), .ZN(n595) );
  NAND2_X1 U633 ( .A1(n845), .A2(n595), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(G284) );
  NAND2_X1 U635 ( .A1(n638), .A2(G89), .ZN(n572) );
  XNOR2_X1 U636 ( .A(n572), .B(KEYINPUT4), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G76), .A2(n631), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(n575), .B(KEYINPUT5), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G51), .A2(n635), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT70), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G63), .A2(n634), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT6), .B(n579), .Z(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U648 ( .A1(G65), .A2(n634), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G53), .A2(n635), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G91), .A2(n638), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G78), .A2(n631), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n972) );
  INV_X1 U655 ( .A(n972), .ZN(G299) );
  NOR2_X1 U656 ( .A1(G286), .A2(n595), .ZN(n590) );
  NOR2_X1 U657 ( .A1(G868), .A2(G299), .ZN(n589) );
  NOR2_X1 U658 ( .A1(n590), .A2(n589), .ZN(G297) );
  INV_X1 U659 ( .A(G860), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n591), .A2(G559), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n592), .A2(n966), .ZN(n593) );
  XNOR2_X1 U662 ( .A(n593), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U663 ( .A1(n966), .A2(G868), .ZN(n594) );
  NOR2_X1 U664 ( .A1(G559), .A2(n594), .ZN(n597) );
  AND2_X1 U665 ( .A1(n595), .A2(n982), .ZN(n596) );
  NOR2_X1 U666 ( .A1(n597), .A2(n596), .ZN(G282) );
  NAND2_X1 U667 ( .A1(G123), .A2(n892), .ZN(n598) );
  XOR2_X1 U668 ( .A(KEYINPUT18), .B(n598), .Z(n599) );
  XNOR2_X1 U669 ( .A(n599), .B(KEYINPUT71), .ZN(n601) );
  NAND2_X1 U670 ( .A1(G111), .A2(n891), .ZN(n600) );
  NAND2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G135), .A2(n887), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G99), .A2(n888), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n922) );
  XNOR2_X1 U676 ( .A(n922), .B(G2096), .ZN(n607) );
  INV_X1 U677 ( .A(G2100), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(G156) );
  NAND2_X1 U679 ( .A1(G93), .A2(n638), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G80), .A2(n631), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n614) );
  NAND2_X1 U682 ( .A1(G67), .A2(n634), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G55), .A2(n635), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U685 ( .A(KEYINPUT73), .B(n612), .Z(n613) );
  NOR2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n649) );
  NAND2_X1 U687 ( .A1(n966), .A2(G559), .ZN(n652) );
  XOR2_X1 U688 ( .A(n982), .B(KEYINPUT72), .Z(n615) );
  XNOR2_X1 U689 ( .A(n652), .B(n615), .ZN(n616) );
  NOR2_X1 U690 ( .A1(G860), .A2(n616), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n649), .B(n617), .ZN(G145) );
  NAND2_X1 U692 ( .A1(G74), .A2(G651), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n618), .A2(G87), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G49), .A2(n635), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U696 ( .A1(n634), .A2(n621), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U698 ( .A(n624), .B(KEYINPUT74), .ZN(G288) );
  NAND2_X1 U699 ( .A1(G88), .A2(n638), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G75), .A2(n631), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U702 ( .A1(G50), .A2(n635), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n634), .A2(G62), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U705 ( .A1(n630), .A2(n629), .ZN(G166) );
  NAND2_X1 U706 ( .A1(n631), .A2(G73), .ZN(n633) );
  XNOR2_X1 U707 ( .A(KEYINPUT76), .B(KEYINPUT2), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n633), .B(n632), .ZN(n643) );
  NAND2_X1 U709 ( .A1(G61), .A2(n634), .ZN(n637) );
  NAND2_X1 U710 ( .A1(G48), .A2(n635), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U712 ( .A1(G86), .A2(n638), .ZN(n639) );
  XNOR2_X1 U713 ( .A(KEYINPUT75), .B(n639), .ZN(n640) );
  NOR2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U715 ( .A1(n643), .A2(n642), .ZN(G305) );
  NOR2_X1 U716 ( .A1(G868), .A2(n649), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n644), .B(KEYINPUT77), .ZN(n655) );
  XNOR2_X1 U718 ( .A(G290), .B(KEYINPUT19), .ZN(n646) );
  XNOR2_X1 U719 ( .A(G166), .B(n972), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U721 ( .A(G288), .B(n647), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n648), .B(G305), .ZN(n651) );
  XOR2_X1 U723 ( .A(n982), .B(n649), .Z(n650) );
  XNOR2_X1 U724 ( .A(n651), .B(n650), .ZN(n841) );
  XNOR2_X1 U725 ( .A(n841), .B(n652), .ZN(n653) );
  NAND2_X1 U726 ( .A1(G868), .A2(n653), .ZN(n654) );
  NAND2_X1 U727 ( .A1(n655), .A2(n654), .ZN(G295) );
  XNOR2_X1 U728 ( .A(KEYINPUT20), .B(KEYINPUT79), .ZN(n658) );
  NAND2_X1 U729 ( .A1(G2084), .A2(G2078), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(KEYINPUT78), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n659), .A2(G2090), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(KEYINPUT21), .ZN(n661) );
  XNOR2_X1 U734 ( .A(KEYINPUT80), .B(n661), .ZN(n662) );
  NAND2_X1 U735 ( .A1(n662), .A2(G2072), .ZN(n663) );
  XOR2_X1 U736 ( .A(KEYINPUT81), .B(n663), .Z(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U738 ( .A1(G220), .A2(G219), .ZN(n664) );
  XOR2_X1 U739 ( .A(KEYINPUT22), .B(n664), .Z(n665) );
  NOR2_X1 U740 ( .A1(G218), .A2(n665), .ZN(n666) );
  NAND2_X1 U741 ( .A1(G96), .A2(n666), .ZN(n839) );
  NAND2_X1 U742 ( .A1(n839), .A2(G2106), .ZN(n670) );
  NAND2_X1 U743 ( .A1(G69), .A2(G120), .ZN(n667) );
  NOR2_X1 U744 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U745 ( .A1(G108), .A2(n668), .ZN(n838) );
  NAND2_X1 U746 ( .A1(n838), .A2(G567), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n670), .A2(n669), .ZN(n848) );
  NAND2_X1 U748 ( .A1(G661), .A2(G483), .ZN(n671) );
  XNOR2_X1 U749 ( .A(KEYINPUT82), .B(n671), .ZN(n672) );
  NOR2_X1 U750 ( .A1(n848), .A2(n672), .ZN(n837) );
  NAND2_X1 U751 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U752 ( .A1(n891), .A2(G113), .ZN(n675) );
  NAND2_X1 U753 ( .A1(G101), .A2(n888), .ZN(n673) );
  XOR2_X1 U754 ( .A(KEYINPUT23), .B(n673), .Z(n674) );
  NAND2_X1 U755 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U756 ( .A1(G125), .A2(n892), .ZN(n677) );
  NAND2_X1 U757 ( .A1(G137), .A2(n887), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U759 ( .A1(n679), .A2(n678), .ZN(G160) );
  XOR2_X1 U760 ( .A(KEYINPUT84), .B(G166), .Z(G303) );
  INV_X1 U761 ( .A(G301), .ZN(G171) );
  NOR2_X1 U762 ( .A1(G1976), .A2(G288), .ZN(n976) );
  NOR2_X1 U763 ( .A1(G303), .A2(G1971), .ZN(n680) );
  NOR2_X1 U764 ( .A1(n976), .A2(n680), .ZN(n749) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n754) );
  INV_X1 U766 ( .A(n754), .ZN(n682) );
  XNOR2_X1 U767 ( .A(n681), .B(KEYINPUT64), .ZN(n753) );
  NAND2_X1 U768 ( .A1(n682), .A2(n753), .ZN(n734) );
  NOR2_X1 U769 ( .A1(G2084), .A2(n734), .ZN(n683) );
  NAND2_X1 U770 ( .A1(n683), .A2(G8), .ZN(n733) );
  NAND2_X1 U771 ( .A1(G8), .A2(n734), .ZN(n796) );
  NOR2_X1 U772 ( .A1(G1966), .A2(n796), .ZN(n731) );
  NOR2_X1 U773 ( .A1(n731), .A2(n683), .ZN(n684) );
  NAND2_X1 U774 ( .A1(G8), .A2(n684), .ZN(n685) );
  XNOR2_X1 U775 ( .A(n685), .B(KEYINPUT30), .ZN(n686) );
  NOR2_X1 U776 ( .A1(G168), .A2(n686), .ZN(n690) );
  XNOR2_X1 U777 ( .A(G1961), .B(KEYINPUT87), .ZN(n1006) );
  NAND2_X1 U778 ( .A1(n734), .A2(n1006), .ZN(n688) );
  INV_X1 U779 ( .A(n734), .ZN(n706) );
  XNOR2_X1 U780 ( .A(G2078), .B(KEYINPUT25), .ZN(n947) );
  NAND2_X1 U781 ( .A1(n706), .A2(n947), .ZN(n687) );
  NAND2_X1 U782 ( .A1(n688), .A2(n687), .ZN(n725) );
  NOR2_X1 U783 ( .A1(G171), .A2(n725), .ZN(n689) );
  NOR2_X1 U784 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U785 ( .A(n691), .B(KEYINPUT31), .ZN(n692) );
  XNOR2_X1 U786 ( .A(n692), .B(KEYINPUT94), .ZN(n729) );
  NAND2_X1 U787 ( .A1(G1956), .A2(n734), .ZN(n693) );
  XOR2_X1 U788 ( .A(KEYINPUT89), .B(n693), .Z(n697) );
  XOR2_X1 U789 ( .A(KEYINPUT88), .B(KEYINPUT27), .Z(n695) );
  NAND2_X1 U790 ( .A1(n706), .A2(G2072), .ZN(n694) );
  XNOR2_X1 U791 ( .A(n695), .B(n694), .ZN(n696) );
  AND2_X1 U792 ( .A1(n697), .A2(n696), .ZN(n718) );
  NOR2_X1 U793 ( .A1(n972), .A2(n718), .ZN(n699) );
  INV_X1 U794 ( .A(KEYINPUT28), .ZN(n698) );
  XNOR2_X1 U795 ( .A(n699), .B(n698), .ZN(n722) );
  NAND2_X1 U796 ( .A1(n734), .A2(G1341), .ZN(n700) );
  XNOR2_X1 U797 ( .A(n700), .B(KEYINPUT90), .ZN(n701) );
  NAND2_X1 U798 ( .A1(n701), .A2(n982), .ZN(n704) );
  AND2_X1 U799 ( .A1(n706), .A2(G1996), .ZN(n702) );
  XNOR2_X1 U800 ( .A(KEYINPUT26), .B(n702), .ZN(n703) );
  NOR2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n705), .A2(n966), .ZN(n715) );
  NAND2_X1 U803 ( .A1(n706), .A2(G2067), .ZN(n707) );
  XNOR2_X1 U804 ( .A(KEYINPUT92), .B(n707), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n734), .A2(G1348), .ZN(n710) );
  NAND2_X1 U806 ( .A1(n708), .A2(n710), .ZN(n709) );
  NOR2_X1 U807 ( .A1(KEYINPUT91), .A2(n709), .ZN(n713) );
  NAND2_X1 U808 ( .A1(KEYINPUT92), .A2(KEYINPUT91), .ZN(n711) );
  NOR2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U810 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U811 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U813 ( .A1(n972), .A2(n718), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n724) );
  XOR2_X1 U816 ( .A(KEYINPUT93), .B(KEYINPUT29), .Z(n723) );
  XNOR2_X1 U817 ( .A(n724), .B(n723), .ZN(n727) );
  AND2_X1 U818 ( .A1(G171), .A2(n725), .ZN(n726) );
  NOR2_X1 U819 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U821 ( .A(KEYINPUT95), .B(n730), .Z(n739) );
  NOR2_X1 U822 ( .A1(n731), .A2(n739), .ZN(n732) );
  NAND2_X1 U823 ( .A1(n733), .A2(n732), .ZN(n748) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n734), .ZN(n735) );
  XNOR2_X1 U825 ( .A(n735), .B(KEYINPUT96), .ZN(n737) );
  NOR2_X1 U826 ( .A1(n796), .A2(G1971), .ZN(n736) );
  NOR2_X1 U827 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U828 ( .A1(G303), .A2(n738), .ZN(n742) );
  INV_X1 U829 ( .A(n739), .ZN(n740) );
  NAND2_X1 U830 ( .A1(n740), .A2(G286), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U832 ( .A1(G8), .A2(n743), .ZN(n746) );
  XOR2_X1 U833 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n744) );
  NAND2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n789) );
  NAND2_X1 U835 ( .A1(n749), .A2(n789), .ZN(n750) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n973) );
  INV_X1 U837 ( .A(n973), .ZN(n751) );
  NOR2_X1 U838 ( .A1(n796), .A2(n751), .ZN(n785) );
  NAND2_X1 U839 ( .A1(n976), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U840 ( .A1(n752), .A2(n796), .ZN(n784) );
  XOR2_X1 U841 ( .A(G1981), .B(G305), .Z(n983) );
  NOR2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n811) );
  INV_X1 U843 ( .A(n811), .ZN(n772) );
  NAND2_X1 U844 ( .A1(G105), .A2(n888), .ZN(n755) );
  XNOR2_X1 U845 ( .A(n755), .B(KEYINPUT38), .ZN(n762) );
  NAND2_X1 U846 ( .A1(G129), .A2(n892), .ZN(n757) );
  NAND2_X1 U847 ( .A1(G141), .A2(n887), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n760) );
  NAND2_X1 U849 ( .A1(G117), .A2(n891), .ZN(n758) );
  XNOR2_X1 U850 ( .A(KEYINPUT85), .B(n758), .ZN(n759) );
  NOR2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n899) );
  NAND2_X1 U853 ( .A1(G1996), .A2(n899), .ZN(n770) );
  NAND2_X1 U854 ( .A1(G107), .A2(n891), .ZN(n764) );
  NAND2_X1 U855 ( .A1(G131), .A2(n887), .ZN(n763) );
  NAND2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n768) );
  NAND2_X1 U857 ( .A1(G119), .A2(n892), .ZN(n766) );
  NAND2_X1 U858 ( .A1(G95), .A2(n888), .ZN(n765) );
  NAND2_X1 U859 ( .A1(n766), .A2(n765), .ZN(n767) );
  OR2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n900) );
  NAND2_X1 U861 ( .A1(G1991), .A2(n900), .ZN(n769) );
  NAND2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n925) );
  XNOR2_X1 U863 ( .A(G1986), .B(G290), .ZN(n968) );
  NOR2_X1 U864 ( .A1(n925), .A2(n968), .ZN(n771) );
  OR2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n798) );
  AND2_X1 U866 ( .A1(n983), .A2(n798), .ZN(n782) );
  XNOR2_X1 U867 ( .A(KEYINPUT37), .B(G2067), .ZN(n809) );
  NAND2_X1 U868 ( .A1(G140), .A2(n887), .ZN(n774) );
  NAND2_X1 U869 ( .A1(G104), .A2(n888), .ZN(n773) );
  NAND2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U871 ( .A(KEYINPUT34), .B(n775), .ZN(n780) );
  NAND2_X1 U872 ( .A1(G116), .A2(n891), .ZN(n777) );
  NAND2_X1 U873 ( .A1(G128), .A2(n892), .ZN(n776) );
  NAND2_X1 U874 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U875 ( .A(KEYINPUT35), .B(n778), .Z(n779) );
  NOR2_X1 U876 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U877 ( .A(KEYINPUT36), .B(n781), .ZN(n909) );
  NOR2_X1 U878 ( .A1(n809), .A2(n909), .ZN(n929) );
  NAND2_X1 U879 ( .A1(n929), .A2(n811), .ZN(n808) );
  NAND2_X1 U880 ( .A1(n782), .A2(n808), .ZN(n783) );
  NOR2_X1 U881 ( .A1(n784), .A2(n783), .ZN(n818) );
  AND2_X1 U882 ( .A1(n785), .A2(n818), .ZN(n786) );
  NAND2_X1 U883 ( .A1(n522), .A2(n786), .ZN(n822) );
  NOR2_X1 U884 ( .A1(G2090), .A2(G303), .ZN(n787) );
  NAND2_X1 U885 ( .A1(G8), .A2(n787), .ZN(n788) );
  NAND2_X1 U886 ( .A1(n789), .A2(n788), .ZN(n792) );
  AND2_X1 U887 ( .A1(n796), .A2(n798), .ZN(n790) );
  AND2_X1 U888 ( .A1(n790), .A2(n808), .ZN(n791) );
  AND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n817) );
  NOR2_X1 U890 ( .A1(G1981), .A2(G305), .ZN(n793) );
  XOR2_X1 U891 ( .A(n793), .B(KEYINPUT86), .Z(n794) );
  XNOR2_X1 U892 ( .A(KEYINPUT24), .B(n794), .ZN(n795) );
  NOR2_X1 U893 ( .A1(n796), .A2(n795), .ZN(n797) );
  AND2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U895 ( .A1(n808), .A2(n799), .ZN(n815) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n899), .ZN(n920) );
  NOR2_X1 U897 ( .A1(G1991), .A2(n900), .ZN(n923) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n800) );
  XNOR2_X1 U899 ( .A(KEYINPUT100), .B(n800), .ZN(n801) );
  NOR2_X1 U900 ( .A1(n923), .A2(n801), .ZN(n802) );
  NOR2_X1 U901 ( .A1(n802), .A2(n925), .ZN(n803) );
  XOR2_X1 U902 ( .A(KEYINPUT101), .B(n803), .Z(n804) );
  NOR2_X1 U903 ( .A1(n920), .A2(n804), .ZN(n805) );
  XOR2_X1 U904 ( .A(KEYINPUT39), .B(n805), .Z(n806) );
  XOR2_X1 U905 ( .A(KEYINPUT102), .B(n806), .Z(n807) );
  NAND2_X1 U906 ( .A1(n808), .A2(n807), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n809), .A2(n909), .ZN(n936) );
  NAND2_X1 U908 ( .A1(n810), .A2(n936), .ZN(n812) );
  NAND2_X1 U909 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U910 ( .A(KEYINPUT103), .B(n813), .Z(n814) );
  NAND2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n818), .A2(KEYINPUT33), .ZN(n819) );
  AND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U916 ( .A(n823), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U917 ( .A(G2430), .B(G2435), .ZN(n832) );
  XNOR2_X1 U918 ( .A(G2454), .B(KEYINPUT104), .ZN(n830) );
  XOR2_X1 U919 ( .A(G2451), .B(G2427), .Z(n825) );
  XNOR2_X1 U920 ( .A(G2438), .B(G2446), .ZN(n824) );
  XNOR2_X1 U921 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U922 ( .A(n826), .B(G2443), .Z(n828) );
  XNOR2_X1 U923 ( .A(G1341), .B(G1348), .ZN(n827) );
  XNOR2_X1 U924 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U925 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n832), .B(n831), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(G14), .ZN(n912) );
  XNOR2_X1 U928 ( .A(KEYINPUT105), .B(n912), .ZN(G401) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U931 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U933 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U935 ( .A(G120), .ZN(G236) );
  INV_X1 U936 ( .A(G96), .ZN(G221) );
  INV_X1 U937 ( .A(G69), .ZN(G235) );
  NOR2_X1 U938 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n840), .B(KEYINPUT106), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  XOR2_X1 U941 ( .A(KEYINPUT114), .B(n841), .Z(n843) );
  XNOR2_X1 U942 ( .A(G286), .B(G171), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U944 ( .A(n845), .B(n844), .Z(n846) );
  NOR2_X1 U945 ( .A1(G37), .A2(n846), .ZN(n847) );
  XOR2_X1 U946 ( .A(KEYINPUT115), .B(n847), .Z(G397) );
  INV_X1 U947 ( .A(n848), .ZN(G319) );
  XOR2_X1 U948 ( .A(G2100), .B(G2096), .Z(n850) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(G2678), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U951 ( .A(KEYINPUT43), .B(G2072), .Z(n852) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U954 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U955 ( .A(G2084), .B(G2078), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(G227) );
  XOR2_X1 U957 ( .A(KEYINPUT108), .B(G1991), .Z(n858) );
  XNOR2_X1 U958 ( .A(G1961), .B(G1996), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U960 ( .A(n859), .B(KEYINPUT41), .Z(n861) );
  XNOR2_X1 U961 ( .A(G1966), .B(G1986), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U963 ( .A(G1976), .B(G1981), .Z(n863) );
  XNOR2_X1 U964 ( .A(G1971), .B(G1956), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U966 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U967 ( .A(KEYINPUT107), .B(G2474), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(G229) );
  NAND2_X1 U969 ( .A1(G124), .A2(n892), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n868), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G112), .A2(n891), .ZN(n869) );
  XOR2_X1 U972 ( .A(KEYINPUT109), .B(n869), .Z(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G136), .A2(n887), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G100), .A2(n888), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U977 ( .A1(n875), .A2(n874), .ZN(G162) );
  NAND2_X1 U978 ( .A1(n891), .A2(G118), .ZN(n876) );
  XNOR2_X1 U979 ( .A(KEYINPUT111), .B(n876), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n892), .A2(G130), .ZN(n877) );
  XOR2_X1 U981 ( .A(KEYINPUT110), .B(n877), .Z(n878) );
  NOR2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U983 ( .A(KEYINPUT112), .B(n880), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G142), .A2(n887), .ZN(n882) );
  NAND2_X1 U985 ( .A1(G106), .A2(n888), .ZN(n881) );
  NAND2_X1 U986 ( .A1(n882), .A2(n881), .ZN(n884) );
  XOR2_X1 U987 ( .A(KEYINPUT113), .B(KEYINPUT45), .Z(n883) );
  XNOR2_X1 U988 ( .A(n884), .B(n883), .ZN(n885) );
  NAND2_X1 U989 ( .A1(n886), .A2(n885), .ZN(n908) );
  NAND2_X1 U990 ( .A1(G139), .A2(n887), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G103), .A2(n888), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G115), .A2(n891), .ZN(n894) );
  NAND2_X1 U994 ( .A1(G127), .A2(n892), .ZN(n893) );
  NAND2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n895), .Z(n896) );
  NOR2_X1 U997 ( .A1(n897), .A2(n896), .ZN(n932) );
  XOR2_X1 U998 ( .A(n932), .B(G162), .Z(n898) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n900), .B(n922), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1003 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1004 ( .A(G160), .B(G164), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1007 ( .A(n910), .B(n909), .Z(n911) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n911), .ZN(G395) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n912), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(G397), .A2(n913), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n914) );
  XOR2_X1 U1012 ( .A(KEYINPUT49), .B(n914), .Z(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(n917), .A2(G395), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(n918), .B(KEYINPUT116), .ZN(G308) );
  INV_X1 U1016 ( .A(G308), .ZN(G225) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1020 ( .A(KEYINPUT51), .B(n921), .Z(n931) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n927) );
  XOR2_X1 U1022 ( .A(G160), .B(G2084), .Z(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n939) );
  XOR2_X1 U1027 ( .A(G2072), .B(n932), .Z(n934) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(n935), .B(KEYINPUT50), .ZN(n937) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n940), .ZN(n942) );
  INV_X1 U1034 ( .A(KEYINPUT55), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n943), .A2(G29), .ZN(n1026) );
  XOR2_X1 U1037 ( .A(G1991), .B(G25), .Z(n944) );
  NAND2_X1 U1038 ( .A1(n944), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1039 ( .A(G2067), .B(G26), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G33), .B(G2072), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n951) );
  XOR2_X1 U1042 ( .A(n947), .B(G27), .Z(n949) );
  XNOR2_X1 U1043 ( .A(G1996), .B(G32), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(n954), .B(KEYINPUT53), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(n955), .B(KEYINPUT117), .ZN(n958) );
  XOR2_X1 U1049 ( .A(G2084), .B(G34), .Z(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT54), .B(n956), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(G35), .B(G2090), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(KEYINPUT55), .B(n961), .ZN(n963) );
  INV_X1 U1055 ( .A(G29), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n964), .A2(G11), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(KEYINPUT118), .B(n965), .ZN(n1024) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XNOR2_X1 U1060 ( .A(n966), .B(G1348), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(G1961), .B(G301), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n981) );
  XOR2_X1 U1064 ( .A(G303), .B(G1971), .Z(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT120), .B(n971), .ZN(n978) );
  XNOR2_X1 U1066 ( .A(n972), .B(G1956), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1070 ( .A(KEYINPUT121), .B(n979), .Z(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n990) );
  XOR2_X1 U1072 ( .A(n982), .B(G1341), .Z(n988) );
  XNOR2_X1 U1073 ( .A(G168), .B(G1966), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(n985), .B(KEYINPUT119), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(KEYINPUT57), .B(n986), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n1021) );
  INV_X1 U1080 ( .A(G16), .ZN(n1019) );
  XOR2_X1 U1081 ( .A(G4), .B(KEYINPUT123), .Z(n994) );
  XNOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT59), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(n994), .B(n993), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(G6), .B(G1981), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(KEYINPUT122), .B(G1956), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(G20), .B(n999), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1091 ( .A(KEYINPUT60), .B(n1002), .Z(n1004) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(KEYINPUT124), .B(n1005), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(n1006), .B(G5), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1016) );
  XNOR2_X1 U1097 ( .A(G1971), .B(G22), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G23), .B(G1976), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G1986), .B(KEYINPUT125), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(n1011), .B(G24), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(n1022), .B(KEYINPUT126), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(n1027), .B(KEYINPUT127), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

