//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n587, new_n589, new_n590, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1115, new_n1116;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n454), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  AND2_X1   g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n475), .A2(G137), .B1(G101), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n475), .A2(G136), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n467), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n483), .B(new_n485), .C1(G124), .C2(new_n487), .ZN(G162));
  INV_X1    g063(.A(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n489), .C1(new_n471), .C2(new_n473), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n467), .A2(G138), .A3(new_n489), .A4(new_n491), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n471), .C2(new_n473), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n499), .A3(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n496), .A2(KEYINPUT69), .A3(new_n500), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n495), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(KEYINPUT71), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n517), .A2(G88), .B1(new_n519), .B2(G50), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT72), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n515), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n526), .B(new_n528), .C1(new_n518), .C2(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n530), .B1(G89), .B2(new_n517), .ZN(G168));
  NAND2_X1  g106(.A1(new_n512), .A2(new_n516), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n518), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n535), .A2(KEYINPUT73), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(KEYINPUT73), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n536), .A2(new_n537), .B1(new_n514), .B2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  AOI22_X1  g115(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n514), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n517), .A2(G81), .ZN(new_n543));
  AOI211_X1 g118(.A(new_n542), .B(new_n543), .C1(G43), .C2(new_n519), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(new_n519), .A2(G53), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT9), .ZN(new_n551));
  NAND2_X1  g126(.A1(G78), .A2(G543), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT74), .ZN(new_n553));
  INV_X1    g128(.A(new_n512), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n556), .A2(G651), .B1(new_n517), .B2(G91), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n551), .A2(new_n557), .ZN(G299));
  INV_X1    g133(.A(G168), .ZN(G286));
  INV_X1    g134(.A(G166), .ZN(G303));
  AOI22_X1  g135(.A1(new_n517), .A2(G87), .B1(new_n519), .B2(G49), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(G288));
  AOI22_X1  g138(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n514), .ZN(new_n565));
  INV_X1    g140(.A(G86), .ZN(new_n566));
  INV_X1    g141(.A(G48), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n532), .A2(new_n566), .B1(new_n518), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G305));
  AOI22_X1  g145(.A1(new_n517), .A2(G85), .B1(new_n519), .B2(G47), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n514), .B2(new_n572), .ZN(G290));
  NAND2_X1  g148(.A1(G301), .A2(G868), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n517), .A2(G92), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT10), .Z(new_n576));
  NAND2_X1  g151(.A1(G79), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G66), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n554), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(G54), .B2(new_n519), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n574), .B1(new_n582), .B2(G868), .ZN(G284));
  OAI21_X1  g158(.A(new_n574), .B1(new_n582), .B2(G868), .ZN(G321));
  MUX2_X1   g159(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g160(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g161(.A(G559), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n582), .B1(new_n587), .B2(G860), .ZN(G148));
  NAND2_X1  g163(.A1(new_n582), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G868), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g166(.A(KEYINPUT75), .B(KEYINPUT11), .ZN(new_n592));
  XNOR2_X1  g167(.A(G323), .B(new_n592), .ZN(G282));
  OAI21_X1  g168(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n594));
  INV_X1    g169(.A(G111), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(G2105), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n487), .A2(G123), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT76), .Z(new_n598));
  AOI211_X1 g173(.A(new_n596), .B(new_n598), .C1(G135), .C2(new_n475), .ZN(new_n599));
  INV_X1    g174(.A(G2096), .ZN(new_n600));
  INV_X1    g175(.A(G2100), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n467), .A2(new_n477), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT13), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n599), .A2(new_n600), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n604), .A2(new_n601), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n605), .B(new_n606), .C1(new_n600), .C2(new_n599), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT77), .Z(G156));
  XOR2_X1   g183(.A(KEYINPUT15), .B(G2435), .Z(new_n609));
  XOR2_X1   g184(.A(KEYINPUT79), .B(G2438), .Z(new_n610));
  XOR2_X1   g185(.A(new_n609), .B(new_n610), .Z(new_n611));
  XNOR2_X1  g186(.A(G2427), .B(G2430), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(KEYINPUT14), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT80), .Z(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n612), .B2(new_n611), .ZN(new_n616));
  XOR2_X1   g191(.A(G1341), .B(G1348), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(G2451), .B(G2454), .Z(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n618), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2443), .B(G2446), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n622), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(G14), .A3(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(G401));
  INV_X1    g203(.A(KEYINPUT18), .ZN(new_n629));
  XOR2_X1   g204(.A(G2084), .B(G2090), .Z(new_n630));
  XNOR2_X1  g205(.A(G2067), .B(G2678), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT17), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n630), .A2(new_n631), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n629), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(new_n601), .ZN(new_n636));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n632), .B2(KEYINPUT18), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(new_n600), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(new_n639), .ZN(G227));
  XOR2_X1   g215(.A(G1971), .B(G1976), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT19), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1956), .B(G2474), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1961), .B(G1966), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT20), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n643), .A2(new_n644), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n642), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n642), .B2(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT81), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1981), .B(G1986), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT82), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1991), .B(G1996), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(G229));
  INV_X1    g236(.A(G16), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G22), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(G166), .B2(new_n662), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT85), .B(G1971), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(KEYINPUT86), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(KEYINPUT86), .ZN(new_n669));
  NOR2_X1   g244(.A1(G6), .A2(G16), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n569), .B2(G16), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT32), .ZN(new_n672));
  INV_X1    g247(.A(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n662), .A2(G23), .ZN(new_n675));
  INV_X1    g250(.A(G288), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n675), .B1(new_n676), .B2(new_n662), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT33), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND4_X1  g254(.A1(new_n668), .A2(new_n669), .A3(new_n674), .A4(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n680), .A2(KEYINPUT34), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(KEYINPUT34), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n662), .A2(G24), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT84), .Z(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G290), .B2(G16), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G1986), .Z(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G25), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT83), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n487), .A2(G119), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n475), .A2(G131), .ZN(new_n691));
  OR2_X1    g266(.A1(G95), .A2(G2105), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n692), .B(G2104), .C1(G107), .C2(new_n489), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n689), .B1(new_n695), .B2(new_n687), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT35), .B(G1991), .Z(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  NOR2_X1   g273(.A1(new_n686), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n681), .A2(new_n682), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT36), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n700), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT30), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT93), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n706), .A2(new_n705), .A3(G28), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n705), .B2(G28), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n687), .B1(new_n705), .B2(G28), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT31), .B(G11), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n599), .B2(G29), .ZN(new_n712));
  INV_X1    g287(.A(G2084), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n479), .A2(new_n687), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G34), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n713), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n714), .A2(new_n713), .A3(new_n717), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n712), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n687), .A2(G35), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G162), .B2(new_n687), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT29), .B(G2090), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n687), .A2(G26), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n487), .A2(G128), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n475), .A2(G140), .ZN(new_n728));
  OR2_X1    g303(.A1(G104), .A2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n729), .B(G2104), .C1(G116), .C2(new_n489), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n726), .B1(new_n732), .B2(new_n687), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2067), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n720), .A2(new_n724), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n544), .A2(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G16), .B2(G19), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT88), .B(G1341), .Z(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G168), .A2(new_n662), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n662), .B2(G21), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n739), .B1(G1966), .B2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G1966), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n737), .A2(new_n738), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n735), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n467), .A2(G127), .ZN(new_n747));
  INV_X1    g322(.A(G115), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n476), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n489), .B1(new_n749), .B2(KEYINPUT89), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(KEYINPUT89), .B2(new_n749), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n489), .A2(G103), .A3(G2104), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT25), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G139), .B2(new_n475), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT90), .Z(new_n756));
  MUX2_X1   g331(.A(G33), .B(new_n756), .S(G29), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2072), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n687), .A2(G32), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n487), .A2(G129), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n475), .A2(G141), .B1(G105), .B2(new_n477), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT26), .Z(new_n763));
  NAND3_X1  g338(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT92), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n759), .B1(new_n766), .B2(new_n687), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n687), .A2(G27), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G164), .B2(new_n687), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT96), .B(G2078), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT97), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n771), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n662), .A2(G4), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n582), .B2(new_n662), .ZN(new_n777));
  INV_X1    g352(.A(G1348), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G5), .A2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT94), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G301), .B2(new_n662), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT95), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n662), .A2(G20), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT23), .Z(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G299), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1956), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n779), .A2(new_n785), .A3(new_n786), .A4(new_n790), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n746), .A2(new_n758), .A3(new_n775), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n704), .A2(new_n792), .ZN(G150));
  INV_X1    g368(.A(G150), .ZN(G311));
  AOI22_X1  g369(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(new_n514), .ZN(new_n796));
  INV_X1    g371(.A(G93), .ZN(new_n797));
  INV_X1    g372(.A(G55), .ZN(new_n798));
  OAI22_X1  g373(.A1(new_n532), .A2(new_n797), .B1(new_n518), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G860), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT37), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n581), .A2(new_n587), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT99), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n544), .B(new_n800), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(KEYINPUT39), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT100), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n801), .B1(new_n810), .B2(KEYINPUT39), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n803), .B1(new_n812), .B2(new_n813), .ZN(G145));
  AOI21_X1  g389(.A(new_n501), .B1(new_n495), .B2(KEYINPUT101), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n493), .A2(new_n494), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n756), .B(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n487), .A2(G130), .B1(G142), .B2(new_n475), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n489), .A2(KEYINPUT102), .A3(G118), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT102), .B1(new_n489), .B2(G118), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n820), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT103), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(new_n603), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n819), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n765), .B(new_n732), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n694), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(G162), .B(new_n479), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n599), .B(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(G37), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n832), .B2(new_n830), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g410(.A(G166), .B(G288), .ZN(new_n836));
  XNOR2_X1  g411(.A(G290), .B(new_n569), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(KEYINPUT104), .B2(KEYINPUT42), .ZN(new_n839));
  NAND2_X1  g414(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n581), .B(G299), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT41), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n808), .B(new_n589), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n842), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(new_n845), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n841), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G868), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(G868), .B2(new_n800), .ZN(G295));
  OAI21_X1  g426(.A(new_n850), .B1(G868), .B2(new_n800), .ZN(G331));
  INV_X1    g427(.A(new_n808), .ZN(new_n853));
  AND2_X1   g428(.A1(G301), .A2(KEYINPUT105), .ZN(new_n854));
  OAI21_X1  g429(.A(G168), .B1(G301), .B2(KEYINPUT105), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n808), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n860), .A3(new_n847), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n859), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n864), .A2(KEYINPUT106), .A3(new_n853), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n863), .A2(new_n865), .B1(new_n808), .B2(new_n859), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n838), .B(new_n861), .C1(new_n866), .C2(new_n844), .ZN(new_n867));
  AOI21_X1  g442(.A(G37), .B1(new_n867), .B2(KEYINPUT107), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n858), .A2(new_n862), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT106), .B1(new_n864), .B2(new_n853), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n843), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n861), .ZN(new_n873));
  INV_X1    g448(.A(new_n838), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n872), .A2(new_n876), .A3(new_n838), .A4(new_n861), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n868), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n847), .B(new_n860), .C1(new_n869), .C2(new_n870), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n858), .A2(new_n860), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(KEYINPUT108), .A3(new_n843), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT108), .B1(new_n882), .B2(new_n843), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n874), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AND4_X1   g461(.A1(KEYINPUT43), .A2(new_n868), .A3(new_n877), .A4(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT44), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n878), .A2(KEYINPUT43), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n868), .A2(new_n879), .A3(new_n886), .A4(new_n877), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(new_n893), .ZN(G397));
  AOI21_X1  g469(.A(G1384), .B1(new_n815), .B2(new_n817), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n895), .A2(KEYINPUT45), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n470), .A2(G40), .A3(new_n478), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT109), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n731), .B(G2067), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT110), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n766), .A2(G1996), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(new_n765), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n899), .A2(G1996), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n697), .A3(new_n695), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n731), .A2(G2067), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n902), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT127), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n908), .A2(new_n914), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n916), .A2(new_n907), .A3(new_n904), .A4(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n918), .B(KEYINPUT47), .Z(new_n919));
  XNOR2_X1  g494(.A(new_n694), .B(new_n697), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT111), .ZN(new_n921));
  AOI211_X1 g496(.A(new_n909), .B(new_n905), .C1(new_n901), .C2(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n899), .A2(G1986), .A3(G290), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n923), .B(KEYINPUT48), .Z(new_n924));
  AOI211_X1 g499(.A(new_n913), .B(new_n919), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT125), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT117), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT114), .B(G8), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(G1384), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n897), .B1(new_n818), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT112), .ZN(new_n932));
  INV_X1    g507(.A(G1384), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n505), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n934), .B2(new_n929), .ZN(new_n935));
  AOI211_X1 g510(.A(KEYINPUT112), .B(KEYINPUT45), .C1(new_n505), .C2(new_n933), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G1971), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n818), .B2(new_n933), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n505), .A2(new_n940), .A3(new_n933), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n898), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G2090), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n928), .B1(new_n939), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n522), .A2(G8), .A3(new_n524), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n948), .B(KEYINPUT55), .Z(new_n949));
  OAI21_X1  g524(.A(new_n927), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n948), .B(KEYINPUT55), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n937), .A2(new_n938), .B1(new_n944), .B2(new_n945), .ZN(new_n952));
  OAI211_X1 g527(.A(KEYINPUT117), .B(new_n951), .C1(new_n952), .C2(new_n928), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n895), .A2(new_n940), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n897), .B1(new_n934), .B2(KEYINPUT50), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n939), .B(new_n955), .C1(G2090), .C2(new_n958), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n493), .A2(new_n494), .B1(new_n501), .B2(new_n502), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n960), .B2(new_n504), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT112), .B1(new_n961), .B2(KEYINPUT45), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n934), .A2(new_n932), .A3(new_n929), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G1971), .B1(new_n964), .B2(new_n931), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n958), .A2(G2090), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT113), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n959), .A2(new_n967), .A3(G8), .A4(new_n949), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n895), .A2(new_n898), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n676), .A2(G1976), .ZN(new_n970));
  INV_X1    g545(.A(new_n928), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT52), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n676), .B2(G1976), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n973), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n569), .A2(new_n673), .ZN(new_n977));
  OAI21_X1  g552(.A(G1981), .B1(new_n565), .B2(new_n568), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(KEYINPUT49), .A3(new_n978), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n969), .A3(new_n971), .A4(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n983), .A2(new_n984), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n976), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n954), .A2(new_n968), .A3(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT124), .B(KEYINPUT51), .Z(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n505), .A2(new_n930), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n898), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n744), .B1(new_n896), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n956), .A2(new_n957), .A3(new_n713), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n991), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(G168), .A2(new_n928), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n995), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n971), .ZN(new_n999));
  OAI221_X1 g574(.A(new_n990), .B1(new_n996), .B2(new_n997), .C1(new_n999), .C2(G168), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n997), .A2(KEYINPUT51), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(G301), .B(KEYINPUT54), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n896), .A2(new_n1004), .A3(G2078), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1003), .B1(new_n931), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1004), .B1(new_n937), .B2(G2078), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n958), .A2(new_n783), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n896), .A2(new_n993), .ZN(new_n1010));
  INV_X1    g585(.A(G2078), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(KEYINPUT53), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1007), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n1003), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1000), .A2(new_n1002), .A3(new_n1009), .A4(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n926), .B1(new_n989), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n999), .A2(G168), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n990), .B1(new_n996), .B2(new_n997), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1002), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1014), .A2(new_n1009), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n988), .A2(new_n968), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(KEYINPUT125), .A4(new_n954), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT123), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1348), .B1(new_n956), .B2(new_n957), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n969), .A2(G2067), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(KEYINPUT60), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT60), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1026), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n582), .B1(new_n1032), .B2(KEYINPUT122), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n958), .A2(new_n778), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1027), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n1035), .A3(KEYINPUT60), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT122), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n581), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1025), .B(new_n1030), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1033), .A2(new_n1038), .B1(KEYINPUT122), .B2(new_n1032), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT123), .B1(new_n1042), .B2(new_n1029), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT61), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT56), .B(G2072), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n931), .B(new_n1046), .C1(new_n935), .C2(new_n936), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n964), .A2(KEYINPUT120), .A3(new_n931), .A4(new_n1046), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g626(.A(G299), .B(KEYINPUT57), .Z(new_n1052));
  INV_X1    g627(.A(G1956), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n941), .B2(new_n943), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(KEYINPUT119), .B(new_n1053), .C1(new_n941), .C2(new_n943), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1051), .A2(new_n1052), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1052), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1045), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1051), .A2(new_n1058), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1052), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1051), .A2(new_n1052), .A3(new_n1058), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(KEYINPUT61), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n969), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT58), .B(G1341), .ZN(new_n1068));
  OAI22_X1  g643(.A1(new_n937), .A2(G1996), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n544), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT59), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1061), .A2(new_n1066), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT121), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1061), .A2(new_n1066), .A3(new_n1074), .A4(new_n1071), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1044), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1028), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n582), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1059), .B1(new_n1064), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1024), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1067), .A2(new_n928), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G288), .A2(G1976), .ZN(new_n1082));
  XOR2_X1   g657(.A(new_n1082), .B(KEYINPUT116), .Z(new_n1083));
  INV_X1    g658(.A(new_n987), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n1084), .B2(new_n985), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n977), .ZN(new_n1086));
  INV_X1    g661(.A(new_n968), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1081), .A2(new_n1086), .B1(new_n1087), .B2(new_n988), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1019), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1002), .B(KEYINPUT62), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1090), .A2(G171), .A3(new_n1013), .A4(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1088), .B1(new_n1092), .B2(new_n989), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n999), .A2(G286), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n954), .A2(new_n968), .A3(new_n988), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT63), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(KEYINPUT63), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n959), .A2(new_n967), .A3(G8), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n951), .B2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1097), .A2(KEYINPUT118), .B1(new_n1022), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1095), .A2(new_n1102), .A3(new_n1096), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1093), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1080), .A2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(G290), .B(G1986), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n898), .A3(new_n896), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n922), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT126), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT126), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1111), .B(new_n1108), .C1(new_n1080), .C2(new_n1104), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n925), .B1(new_n1110), .B2(new_n1112), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g688(.A1(G227), .A2(new_n465), .ZN(new_n1115));
  NOR3_X1   g689(.A1(G401), .A2(G229), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n1116), .A3(new_n834), .ZN(G225));
  INV_X1    g691(.A(G225), .ZN(G308));
endmodule


