//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n210), .A2(G20), .A3(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n208), .B(new_n213), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G250), .B(G257), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT64), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n229), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G150), .ZN(new_n244));
  NOR3_X1   g0044(.A1(new_n244), .A2(G20), .A3(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G20), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G50), .A2(G58), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n246), .B1(new_n247), .B2(new_n215), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G58), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT8), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT8), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G58), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI211_X1 g0055(.A(new_n245), .B(new_n248), .C1(new_n250), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n211), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n258), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(G20), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G50), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G50), .B2(new_n262), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G222), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  OAI221_X1 g0075(.A(new_n272), .B1(new_n273), .B2(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n278), .A2(G274), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n283), .A2(G226), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G190), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(G200), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n269), .A2(new_n291), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n290), .A2(G169), .B1(new_n260), .B2(new_n267), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n289), .A2(G179), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n263), .A2(new_n215), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT12), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G20), .A2(G33), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n303), .A2(G50), .B1(G20), .B2(new_n215), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n273), .B2(new_n249), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n264), .A2(G68), .A3(new_n265), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n302), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT11), .B1(new_n305), .B2(new_n258), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT71), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n287), .A2(new_n278), .A3(G274), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n216), .B2(new_n282), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n270), .A2(G232), .A3(G1698), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n270), .A2(G226), .A3(new_n271), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n314), .B1(new_n318), .B2(new_n279), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT14), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(new_n322), .A3(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n320), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n324), .B(G179), .C1(new_n325), .C2(new_n319), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n322), .B1(new_n321), .B2(G169), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n312), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n324), .B(G190), .C1(new_n325), .C2(new_n319), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n310), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT70), .B1(new_n321), .B2(G200), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n321), .A2(KEYINPUT70), .A3(G200), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT17), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT7), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n270), .A2(new_n340), .A3(G20), .ZN(new_n341));
  INV_X1    g0141(.A(G33), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT3), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT3), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G33), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT7), .B1(new_n346), .B2(new_n246), .ZN(new_n347));
  OAI21_X1  g0147(.A(G68), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g0148(.A(G58), .B(G68), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G20), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT72), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n303), .A2(new_n351), .A3(G159), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(new_n303), .B2(G159), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n339), .B1(new_n348), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n340), .B1(new_n270), .B2(G20), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n346), .A2(KEYINPUT7), .A3(new_n246), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n215), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n360), .A2(KEYINPUT16), .A3(new_n355), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n258), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n264), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n255), .A2(new_n265), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n363), .A2(new_n364), .B1(new_n262), .B2(new_n255), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n343), .A2(new_n345), .A3(G223), .A4(new_n271), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n343), .A2(new_n345), .A3(G226), .A4(G1698), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G87), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n279), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n278), .A2(G232), .A3(new_n281), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n313), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  AND4_X1   g0176(.A1(KEYINPUT73), .A2(new_n372), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n374), .B1(new_n279), .B2(new_n371), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n376), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT73), .B1(new_n378), .B2(G200), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n338), .B1(new_n367), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT18), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n372), .A2(new_n375), .ZN(new_n384));
  INV_X1    g0184(.A(G169), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G179), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n378), .A2(new_n387), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n367), .A2(new_n383), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n348), .A2(new_n356), .A3(new_n339), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT16), .B1(new_n360), .B2(new_n355), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n365), .B1(new_n393), .B2(new_n258), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n386), .A2(new_n388), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT18), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n378), .A2(KEYINPUT73), .A3(new_n376), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT73), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n384), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n384), .A2(G190), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n394), .A2(new_n402), .A3(KEYINPUT17), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n382), .A2(new_n390), .A3(new_n396), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n255), .A2(new_n303), .B1(G20), .B2(G77), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT15), .B(G87), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT67), .B1(new_n407), .B2(new_n249), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n407), .A2(KEYINPUT67), .A3(new_n249), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n258), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT68), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n411), .B(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n273), .B1(new_n261), .B2(G20), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n264), .A2(new_n414), .B1(new_n273), .B2(new_n263), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n283), .A2(G244), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n313), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT66), .ZN(new_n419));
  INV_X1    g0219(.A(G107), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n274), .A2(new_n216), .B1(new_n420), .B2(new_n270), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n346), .A2(new_n231), .A3(G1698), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n279), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT66), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n417), .A2(new_n424), .A3(new_n313), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n419), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n385), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n426), .A2(G179), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n416), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(G200), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n376), .B2(new_n426), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n416), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n300), .A2(new_n337), .A3(new_n405), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT78), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT5), .B(G41), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n286), .A2(G1), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n437), .A2(new_n438), .B1(new_n212), .B2(new_n277), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G257), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n261), .A2(G45), .ZN(new_n441));
  NOR2_X1   g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n284), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT77), .ZN(new_n448));
  INV_X1    g0248(.A(G244), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(G1698), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n343), .A3(new_n345), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT76), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n450), .A2(new_n343), .A3(new_n345), .A4(KEYINPUT4), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n343), .A2(new_n345), .A3(G250), .A4(G1698), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G283), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n452), .B1(new_n451), .B2(new_n453), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n454), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n448), .B1(new_n460), .B2(new_n278), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n451), .A2(new_n453), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT76), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(KEYINPUT77), .A3(new_n279), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n447), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n436), .B1(new_n468), .B2(new_n399), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n440), .A2(new_n446), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n466), .A2(KEYINPUT77), .A3(new_n279), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT77), .B1(new_n466), .B2(new_n279), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(KEYINPUT78), .A3(G200), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n420), .A2(KEYINPUT6), .A3(G97), .ZN(new_n475));
  AND2_X1   g0275(.A1(G97), .A2(G107), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n202), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n477), .B2(KEYINPUT6), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G20), .B1(G77), .B2(new_n303), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n420), .B1(new_n358), .B2(new_n359), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT74), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI211_X1 g0282(.A(KEYINPUT74), .B(new_n420), .C1(new_n358), .C2(new_n359), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n258), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n262), .A2(G97), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n261), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n262), .A2(new_n486), .A3(new_n211), .A4(new_n257), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n485), .B1(new_n488), .B2(G97), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n470), .B1(new_n460), .B2(new_n278), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n376), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n469), .A2(new_n474), .A3(new_n493), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n484), .A2(new_n489), .B1(new_n491), .B2(new_n385), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n387), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n439), .A2(G270), .B1(new_n284), .B2(new_n445), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n344), .A2(G33), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n342), .A2(KEYINPUT3), .ZN(new_n501));
  OAI21_X1  g0301(.A(G303), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n343), .A2(new_n345), .A3(G264), .A4(G1698), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n343), .A2(new_n345), .A3(G257), .A4(new_n271), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n279), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G116), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n263), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n259), .A2(G116), .A3(new_n262), .A4(new_n486), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n257), .A2(new_n211), .B1(G20), .B2(new_n508), .ZN(new_n511));
  INV_X1    g0311(.A(G97), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n457), .B(new_n246), .C1(G33), .C2(new_n512), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n511), .A2(KEYINPUT20), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT20), .B1(new_n511), .B2(new_n513), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n509), .B(new_n510), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n507), .A2(KEYINPUT21), .A3(G169), .A4(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n385), .B1(new_n499), .B2(new_n506), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n520), .A2(KEYINPUT81), .A3(KEYINPUT21), .A4(new_n516), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n516), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT21), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n499), .A2(new_n506), .A3(G179), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n516), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n516), .B1(new_n507), .B2(G200), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n376), .B2(new_n507), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n522), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n343), .A2(new_n345), .A3(new_n246), .A4(G87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT22), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT22), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n270), .A2(new_n533), .A3(new_n246), .A4(G87), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT23), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n536), .A2(new_n246), .A3(G107), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT23), .B1(new_n420), .B2(G20), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G116), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n537), .A2(new_n538), .B1(G20), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(KEYINPUT82), .B(new_n530), .C1(new_n535), .C2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n532), .B2(new_n534), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT82), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT24), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI211_X1 g0344(.A(KEYINPUT82), .B(new_n540), .C1(new_n532), .C2(new_n534), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n541), .B(new_n258), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n420), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT25), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n262), .B2(G107), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n488), .A2(G107), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n343), .A2(new_n345), .A3(G257), .A4(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n343), .A2(new_n345), .A3(G250), .A4(new_n271), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G294), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n279), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT84), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n439), .A2(new_n557), .A3(G264), .ZN(new_n558));
  INV_X1    g0358(.A(new_n444), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n438), .B1(new_n559), .B2(new_n442), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(G264), .A3(new_n278), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT84), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n556), .A2(new_n558), .A3(new_n562), .A4(new_n446), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n563), .A2(new_n387), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n556), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n555), .A2(KEYINPUT83), .A3(new_n279), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n446), .A2(new_n561), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G169), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n551), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n343), .A2(new_n345), .A3(G244), .A4(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n343), .A2(new_n345), .A3(G238), .A4(new_n271), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n574), .A3(new_n539), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n279), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n438), .A2(new_n218), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n284), .A2(new_n438), .B1(new_n577), .B2(new_n278), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n387), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(new_n578), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n385), .ZN(new_n583));
  INV_X1    g0383(.A(new_n407), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(new_n262), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n246), .B1(new_n317), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G87), .B2(new_n203), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n343), .A2(new_n345), .A3(new_n246), .A4(G68), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n586), .B1(new_n249), .B2(new_n512), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n585), .B1(new_n591), .B2(new_n258), .ZN(new_n592));
  OR3_X1    g0392(.A1(new_n487), .A2(KEYINPUT80), .A3(new_n407), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT80), .B1(new_n487), .B2(new_n407), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n576), .A2(new_n578), .A3(KEYINPUT79), .A4(new_n387), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n581), .A2(new_n583), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n582), .A2(G200), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n487), .A2(new_n217), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n600), .B(new_n585), .C1(new_n591), .C2(new_n258), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n576), .A2(G190), .A3(new_n578), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n563), .A2(new_n399), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n569), .B2(G190), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n546), .A3(new_n550), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n572), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  NOR4_X1   g0408(.A1(new_n435), .A2(new_n498), .A3(new_n529), .A4(new_n608), .ZN(G372));
  INV_X1    g0409(.A(new_n435), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT86), .ZN(new_n611));
  INV_X1    g0411(.A(new_n578), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT85), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n576), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n575), .A2(KEYINPUT85), .A3(new_n279), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n611), .B1(new_n616), .B2(G169), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n575), .A2(KEYINPUT85), .A3(new_n279), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT85), .B1(new_n575), .B2(new_n279), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n578), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(KEYINPUT86), .A3(new_n385), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n596), .A2(new_n579), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n602), .B(new_n601), .C1(new_n616), .C2(new_n399), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n623), .A2(new_n607), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n572), .A2(new_n522), .A3(new_n526), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(new_n494), .A4(new_n497), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n495), .A2(new_n496), .A3(new_n603), .A4(new_n598), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n621), .A2(new_n622), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n628), .A2(KEYINPUT26), .B1(new_n617), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n601), .A2(new_n602), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(G200), .B2(new_n620), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n629), .B2(new_n617), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n495), .A2(new_n496), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n627), .B(new_n630), .C1(KEYINPUT26), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n610), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n298), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n390), .A2(new_n396), .ZN(new_n639));
  INV_X1    g0439(.A(new_n335), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n310), .B(new_n331), .C1(new_n640), .C2(new_n333), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n330), .B1(new_n641), .B2(new_n430), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n382), .A2(new_n403), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n639), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n638), .B1(new_n645), .B2(new_n295), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n637), .A2(new_n646), .ZN(G369));
  NAND2_X1  g0447(.A1(new_n522), .A2(new_n526), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n261), .A2(new_n246), .A3(G13), .ZN(new_n649));
  OAI21_X1  g0449(.A(G213), .B1(new_n649), .B2(KEYINPUT27), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT87), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n649), .B2(KEYINPUT27), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n649), .A2(new_n651), .A3(KEYINPUT27), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G343), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n657), .A2(new_n516), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n529), .B2(new_n658), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n660), .A2(G330), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n572), .A2(new_n607), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n656), .B1(new_n546), .B2(new_n550), .ZN(new_n663));
  OAI22_X1  g0463(.A1(new_n662), .A2(new_n663), .B1(new_n572), .B2(new_n656), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n657), .B1(new_n522), .B2(new_n526), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT88), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n664), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n546), .A2(new_n550), .B1(new_n564), .B2(new_n570), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n656), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n665), .A2(new_n668), .A3(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n206), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G1), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n209), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n627), .A2(KEYINPUT90), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n648), .A2(new_n669), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n623), .A2(new_n607), .A3(new_n624), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n484), .B(new_n489), .C1(new_n376), .C2(new_n491), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n461), .A2(new_n467), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n399), .B1(new_n685), .B2(new_n470), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n684), .B1(new_n686), .B2(KEYINPUT78), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n634), .B1(new_n687), .B2(new_n469), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT90), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n683), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n623), .B1(new_n628), .B2(KEYINPUT26), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(KEYINPUT26), .B2(new_n635), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n680), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n679), .B1(new_n693), .B2(new_n656), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n636), .A2(new_n679), .A3(new_n656), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n556), .A2(new_n558), .A3(new_n562), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n582), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n447), .B1(new_n466), .B2(new_n279), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(new_n699), .A3(new_n525), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT30), .A4(new_n525), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n620), .A2(new_n387), .A3(new_n507), .A4(new_n563), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n468), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT89), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n563), .A2(new_n387), .A3(new_n507), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n473), .A2(new_n620), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT89), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(new_n702), .A4(new_n703), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n657), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n608), .A2(new_n529), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n688), .A3(new_n656), .ZN(new_n716));
  OAI211_X1 g0516(.A(KEYINPUT31), .B(new_n657), .C1(new_n704), .C2(new_n706), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n696), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n678), .B1(new_n721), .B2(G1), .ZN(G364));
  AND2_X1   g0522(.A1(new_n246), .A2(G13), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n261), .B1(new_n723), .B2(G45), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n673), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n661), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(G330), .B2(new_n660), .ZN(new_n728));
  INV_X1    g0528(.A(G355), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n270), .A2(new_n206), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n729), .A2(new_n730), .B1(G116), .B2(new_n206), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n239), .A2(new_n286), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n672), .A2(new_n270), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n286), .B2(new_n210), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n731), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n211), .B1(G20), .B2(new_n385), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT91), .Z(new_n742));
  OAI21_X1  g0542(.A(new_n726), .B1(new_n736), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n740), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n246), .A2(new_n387), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(G190), .A3(new_n399), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G190), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n747), .A2(G58), .B1(new_n750), .B2(G77), .ZN(new_n751));
  INV_X1    g0551(.A(G50), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n745), .A2(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n376), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n751), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n246), .A2(G179), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n748), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G159), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT32), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(new_n376), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n420), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n756), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n376), .A2(G179), .A3(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n246), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n512), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n753), .A2(G190), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(G68), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT93), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n270), .B1(new_n771), .B2(new_n217), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT92), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n764), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G283), .ZN(new_n775));
  INV_X1    g0575(.A(G329), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n762), .A2(new_n775), .B1(new_n758), .B2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT94), .Z(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n346), .B1(new_n746), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(G311), .B2(new_n750), .ZN(new_n781));
  INV_X1    g0581(.A(new_n766), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G294), .A2(new_n782), .B1(new_n754), .B2(G326), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  INV_X1    g0584(.A(new_n771), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n768), .A2(new_n784), .B1(new_n785), .B2(G303), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n778), .A2(new_n781), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n744), .B1(new_n774), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n743), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n739), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n660), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n728), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  INV_X1    g0593(.A(new_n768), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n794), .A2(KEYINPUT95), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(KEYINPUT95), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n762), .A2(new_n217), .B1(new_n758), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n798), .A2(G283), .B1(KEYINPUT96), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n346), .B1(new_n749), .B2(new_n508), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G294), .B2(new_n747), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n771), .A2(new_n420), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n804), .B(new_n767), .C1(G303), .C2(new_n754), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n800), .A2(KEYINPUT96), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n801), .A2(new_n803), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n270), .B1(new_n758), .B2(new_n808), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n752), .A2(new_n771), .B1(new_n762), .B2(new_n215), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(G58), .C2(new_n782), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT97), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n747), .A2(G143), .B1(new_n750), .B2(G159), .ZN(new_n813));
  INV_X1    g0613(.A(G137), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n794), .B2(new_n244), .C1(new_n814), .C2(new_n755), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT34), .Z(new_n816));
  OAI21_X1  g0616(.A(new_n807), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n744), .B1(new_n817), .B2(KEYINPUT98), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(KEYINPUT98), .B2(new_n817), .ZN(new_n819));
  INV_X1    g0619(.A(new_n726), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n740), .A2(new_n737), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(new_n273), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n430), .A2(new_n656), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n656), .B1(new_n413), .B2(new_n415), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n429), .B1(new_n433), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n819), .B(new_n822), .C1(new_n738), .C2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n636), .B2(new_n656), .ZN(new_n828));
  INV_X1    g0628(.A(new_n627), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n630), .B1(new_n635), .B2(KEYINPUT26), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n656), .B(new_n826), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT99), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n636), .A2(KEYINPUT99), .A3(new_n656), .A4(new_n826), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n828), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n719), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n820), .B1(new_n835), .B2(new_n836), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n827), .B1(new_n838), .B2(new_n839), .ZN(G384));
  NAND4_X1  g0640(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n657), .A4(new_n711), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n714), .A2(new_n716), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n823), .A2(new_n825), .ZN(new_n843));
  INV_X1    g0643(.A(new_n328), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n844), .A2(new_n326), .A3(new_n323), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n312), .B(new_n657), .C1(new_n336), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n312), .A2(new_n657), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n641), .A2(new_n329), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n843), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT40), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n259), .B1(new_n391), .B2(new_n392), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n389), .A2(new_n655), .B1(new_n852), .B2(new_n365), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n394), .A2(new_n402), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n856), .A2(KEYINPUT102), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n655), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n394), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n404), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n857), .B1(new_n853), .B2(new_n854), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT102), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n859), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n856), .A2(new_n858), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n862), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n851), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n850), .A2(new_n871), .A3(KEYINPUT103), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT103), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n404), .A2(new_n861), .B1(new_n864), .B2(new_n863), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n874), .B2(new_n859), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n862), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT40), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n842), .A2(new_n849), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n873), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n862), .B2(new_n869), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n842), .A3(new_n849), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n872), .A2(new_n879), .B1(new_n851), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n610), .A2(new_n842), .ZN(new_n885));
  OAI21_X1  g0685(.A(G330), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n885), .B2(new_n884), .ZN(new_n887));
  INV_X1    g0687(.A(new_n823), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n833), .B2(new_n834), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n876), .A2(new_n880), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n846), .A2(new_n848), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT39), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n875), .B2(new_n876), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n881), .B2(new_n894), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n330), .A2(new_n656), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n896), .A2(new_n897), .B1(new_n639), .B2(new_n655), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n646), .B1(new_n696), .B2(new_n435), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n887), .A2(new_n901), .B1(new_n261), .B2(new_n723), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n901), .B2(new_n887), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n211), .A2(new_n246), .A3(new_n508), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n478), .B(KEYINPUT100), .Z(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT35), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n907), .B2(new_n906), .ZN(new_n909));
  XOR2_X1   g0709(.A(KEYINPUT101), .B(KEYINPUT36), .Z(new_n910));
  XNOR2_X1  g0710(.A(new_n909), .B(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n210), .B(G77), .C1(new_n251), .C2(new_n215), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n752), .A2(G68), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n261), .B(G13), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  OR3_X1    g0714(.A1(new_n903), .A2(new_n911), .A3(new_n914), .ZN(G367));
  NOR2_X1   g0715(.A1(new_n601), .A2(new_n656), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT104), .Z(new_n917));
  NAND2_X1  g0717(.A1(new_n633), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n623), .B2(new_n917), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT105), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n490), .A2(new_n657), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n688), .A2(new_n922), .B1(new_n634), .B2(new_n657), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT42), .B1(new_n668), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n688), .A2(new_n669), .A3(new_n922), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n497), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n656), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n668), .A2(new_n923), .A3(KEYINPUT42), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n921), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n665), .A2(new_n923), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n673), .B(KEYINPUT41), .Z(new_n935));
  NAND2_X1  g0735(.A1(new_n668), .A2(new_n670), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n923), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT107), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT44), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n936), .A2(new_n923), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n661), .A3(new_n664), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n661), .B(new_n664), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(new_n667), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n940), .A2(new_n665), .A3(new_n941), .A4(new_n944), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n946), .A2(new_n721), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n935), .B1(new_n950), .B2(new_n721), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n934), .B1(new_n951), .B2(new_n725), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n229), .A2(new_n734), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n741), .B1(new_n206), .B2(new_n407), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n726), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G50), .A2(new_n750), .B1(new_n759), .B2(G137), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n956), .B(new_n270), .C1(new_n244), .C2(new_n746), .ZN(new_n957));
  INV_X1    g0757(.A(new_n762), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n754), .A2(G143), .B1(new_n958), .B2(G77), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n959), .B1(new_n251), .B2(new_n771), .C1(new_n215), .C2(new_n766), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n957), .B(new_n960), .C1(new_n798), .C2(G159), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G107), .A2(new_n782), .B1(new_n754), .B2(G311), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n270), .B1(new_n759), .B2(G317), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n747), .A2(G303), .B1(new_n750), .B2(G283), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n958), .A2(G97), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT108), .B1(new_n771), .B2(new_n508), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT46), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n966), .B(new_n968), .C1(new_n798), .C2(G294), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n961), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n955), .B1(new_n972), .B2(new_n740), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n790), .B2(new_n919), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n952), .A2(KEYINPUT110), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT110), .B1(new_n952), .B2(new_n974), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(G387));
  AOI22_X1  g0778(.A1(new_n747), .A2(G317), .B1(new_n750), .B2(G303), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n779), .B2(new_n755), .C1(new_n797), .C2(new_n799), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT48), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n782), .A2(G283), .B1(new_n785), .B2(G294), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT49), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n762), .A2(new_n508), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n270), .B(new_n989), .C1(G326), .C2(new_n759), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n746), .A2(new_n752), .B1(new_n749), .B2(new_n215), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n346), .B(new_n992), .C1(G150), .C2(new_n759), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n754), .A2(G159), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n768), .A2(new_n255), .B1(new_n785), .B2(G77), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n782), .A2(new_n584), .B1(new_n958), .B2(G97), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n744), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n664), .A2(new_n790), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n675), .A2(new_n730), .B1(G107), .B2(new_n206), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n234), .A2(new_n286), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT111), .Z(new_n1002));
  INV_X1    g0802(.A(new_n675), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1003), .A2(KEYINPUT112), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(KEYINPUT112), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n286), .B1(new_n215), .B2(new_n273), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n255), .A2(new_n752), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT50), .Z(new_n1009));
  AOI21_X1  g0809(.A(new_n734), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1000), .B1(new_n1002), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n726), .B1(new_n1011), .B2(new_n742), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n998), .A2(new_n999), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n948), .B2(new_n725), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n721), .A2(new_n948), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n673), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n721), .A2(new_n948), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT113), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(G393));
  NAND2_X1  g0822(.A1(new_n946), .A2(new_n949), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n923), .A2(new_n739), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n741), .B1(new_n512), .B2(new_n206), .C1(new_n242), .C2(new_n734), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n726), .ZN(new_n1027));
  INV_X1    g0827(.A(G159), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n755), .A2(new_n244), .B1(new_n1028), .B2(new_n746), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT51), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n782), .A2(G77), .B1(new_n750), .B2(new_n255), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n752), .C2(new_n797), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n346), .B1(new_n759), .B2(G143), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n215), .B2(new_n771), .C1(new_n217), .C2(new_n762), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT114), .Z(new_n1035));
  AOI22_X1  g0835(.A1(G317), .A2(new_n754), .B1(new_n747), .B2(G311), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n346), .B1(new_n758), .B2(new_n779), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G294), .B2(new_n750), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n771), .A2(new_n775), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n763), .B(new_n1040), .C1(G116), .C2(new_n782), .ZN(new_n1041));
  INV_X1    g0841(.A(G303), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1039), .B(new_n1041), .C1(new_n797), .C2(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1032), .A2(new_n1035), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT115), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1027), .B1(new_n1045), .B2(new_n740), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1024), .A2(new_n725), .B1(new_n1025), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1023), .A2(new_n1015), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n673), .A3(new_n950), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(G390));
  NAND3_X1  g0850(.A1(new_n693), .A2(new_n656), .A3(new_n825), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n823), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT116), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1051), .A2(KEYINPUT116), .A3(new_n823), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n891), .A3(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n868), .A2(new_n870), .B1(new_n330), .B2(new_n656), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n897), .B1(new_n889), .B2(new_n892), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1056), .A2(new_n1057), .B1(new_n1058), .B2(new_n896), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n842), .A2(new_n849), .A3(G330), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1058), .A2(new_n896), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n718), .A2(G330), .A3(new_n826), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n891), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1062), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1061), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n610), .A2(G330), .A3(new_n842), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n646), .C1(new_n696), .C2(new_n435), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n842), .A2(G330), .A3(new_n826), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n892), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1055), .ZN(new_n1074));
  AOI21_X1  g0874(.A(KEYINPUT116), .B1(new_n1051), .B2(new_n823), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1066), .B(new_n1073), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n889), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1060), .B1(new_n1065), .B2(new_n891), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1071), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(KEYINPUT117), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n674), .B1(new_n1069), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(KEYINPUT117), .B(new_n1081), .C1(new_n1061), .C2(new_n1068), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1067), .B(new_n725), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n821), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n726), .B1(new_n1087), .B2(new_n255), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n771), .A2(new_n244), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT53), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n797), .B2(new_n814), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G159), .A2(new_n782), .B1(new_n754), .B2(G128), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(KEYINPUT54), .B(G143), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n346), .B1(new_n750), .B2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n747), .A2(G132), .B1(new_n759), .B2(G125), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n958), .A2(G50), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1092), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n797), .A2(new_n420), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G77), .A2(new_n782), .B1(new_n754), .B2(G283), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n270), .B1(new_n747), .B2(G116), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G97), .A2(new_n750), .B1(new_n759), .B2(G294), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n785), .A2(G87), .B1(new_n958), .B2(G68), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1091), .A2(new_n1098), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1088), .B1(new_n1105), .B2(new_n740), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n896), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n738), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1086), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1085), .A2(new_n1110), .ZN(G378));
  OR2_X1    g0911(.A1(new_n893), .A2(new_n898), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n882), .A2(new_n851), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT103), .B1(new_n850), .B2(new_n871), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n877), .A2(new_n878), .A3(new_n873), .ZN(new_n1115));
  OAI211_X1 g0915(.A(G330), .B(new_n1113), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT120), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n299), .B(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n268), .A2(new_n860), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT119), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1119), .B(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1116), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1122), .B1(new_n883), .B2(G330), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1112), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1116), .A2(new_n1123), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n883), .A2(G330), .A3(new_n1122), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n899), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n724), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1123), .A2(new_n737), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n726), .B1(new_n1087), .B2(G50), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n752), .B1(G33), .B2(G41), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n346), .B2(new_n285), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n794), .A2(new_n512), .B1(new_n755), .B2(new_n508), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G58), .B2(new_n958), .ZN(new_n1136));
  AOI211_X1 g0936(.A(G41), .B(new_n270), .C1(new_n750), .C2(new_n584), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n747), .A2(G107), .B1(new_n759), .B2(G283), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n782), .A2(G68), .B1(new_n785), .B2(G77), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT58), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1134), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(G33), .B(G41), .C1(new_n759), .C2(G124), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G128), .A2(new_n747), .B1(new_n785), .B2(new_n1094), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT118), .Z(new_n1145));
  AOI22_X1  g0945(.A1(new_n754), .A2(G125), .B1(new_n750), .B2(G137), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G150), .A2(new_n782), .B1(new_n768), .B2(G132), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT59), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1143), .B1(new_n1028), .B2(new_n762), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1142), .B1(new_n1141), .B2(new_n1140), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1132), .B1(new_n1152), .B2(new_n740), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1131), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1130), .A2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1067), .B(new_n1080), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1071), .B(KEYINPUT121), .Z(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT122), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT122), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1159), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1157), .A2(new_n1158), .B1(new_n1129), .B2(new_n1126), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n673), .B1(new_n1167), .B2(KEYINPUT57), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1156), .B1(new_n1166), .B2(new_n1168), .ZN(G375));
  INV_X1    g0969(.A(new_n935), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1076), .A2(new_n1071), .A3(new_n1079), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1081), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n724), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n891), .A2(new_n738), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT123), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n270), .B1(new_n759), .B2(G303), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n420), .B2(new_n749), .C1(new_n775), .C2(new_n746), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n754), .A2(G294), .B1(new_n785), .B2(G97), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n273), .B2(new_n762), .C1(new_n407), .C2(new_n766), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(new_n798), .C2(G116), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n346), .B1(new_n759), .B2(G128), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n814), .B2(new_n746), .C1(new_n244), .C2(new_n749), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n754), .A2(G132), .B1(new_n958), .B2(G58), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n752), .B2(new_n766), .C1(new_n1028), .C2(new_n771), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(new_n798), .C2(new_n1094), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n740), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n820), .B1(new_n215), .B2(new_n821), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1173), .B1(new_n1175), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1172), .A2(new_n1189), .ZN(G381));
  NAND3_X1  g0990(.A1(new_n1020), .A2(new_n792), .A3(new_n1021), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(G390), .A2(G384), .A3(new_n1191), .A4(G381), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n976), .B2(new_n977), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1193), .A2(G378), .A3(G375), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT124), .ZN(G407));
  INV_X1    g0995(.A(G213), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1156), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1159), .A2(new_n1164), .A3(new_n1161), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1164), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1167), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n674), .B1(new_n1201), .B2(new_n1160), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1197), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(G378), .A2(G343), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1196), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1194), .A2(KEYINPUT124), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1194), .A2(KEYINPUT124), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(G409));
  NAND2_X1  g1008(.A1(new_n952), .A2(new_n974), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT110), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OR2_X1    g1011(.A1(G390), .A2(KEYINPUT126), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(G390), .A2(KEYINPUT126), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1211), .A2(new_n975), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n952), .A2(G390), .A3(new_n974), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G393), .A2(G396), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1191), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(G390), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1209), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1215), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1217), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1214), .A2(new_n1218), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT60), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1171), .B1(new_n1080), .B2(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n1071), .A4(new_n1079), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n673), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1189), .ZN(new_n1228));
  INV_X1    g1028(.A(G384), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(G384), .A3(new_n1189), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1196), .A2(G343), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(G2897), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1232), .B(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT125), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1130), .B2(new_n1155), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1159), .A2(new_n1170), .A3(new_n1238), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1127), .A2(new_n899), .A3(new_n1128), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n899), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n725), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(KEYINPUT125), .A3(new_n1154), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1237), .A2(new_n1239), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1109), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1203), .B2(G378), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1235), .B1(new_n1247), .B2(new_n1233), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT61), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G378), .B(new_n1156), .C1(new_n1166), .C2(new_n1168), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1232), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT62), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1233), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1248), .A2(new_n1249), .A3(new_n1256), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1233), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1259), .B2(new_n1253), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1223), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT63), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n1232), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1214), .A2(new_n1218), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT61), .B1(new_n1263), .B2(new_n1235), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1259), .A2(KEYINPUT63), .A3(new_n1253), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1264), .A2(new_n1267), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1261), .A2(new_n1270), .ZN(G405));
  NAND2_X1  g1071(.A1(G375), .A2(new_n1245), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1250), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1253), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(new_n1232), .A3(new_n1250), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(new_n1223), .ZN(G402));
endmodule


