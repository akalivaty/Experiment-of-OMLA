//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(G125), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT65), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT66), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n460), .A2(new_n461), .B1(G113), .B2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(new_n470), .B2(new_n464), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n469), .A2(G137), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n469), .A2(G2104), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n463), .A2(new_n475), .B1(new_n476), .B2(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n458), .A2(new_n459), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(KEYINPUT67), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n463), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(G2105), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n481), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n469), .B1(new_n483), .B2(new_n485), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n488), .B1(G136), .B2(new_n490), .ZN(G162));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n494), .A3(G2104), .ZN(new_n495));
  AND2_X1   g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n458), .B2(new_n459), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n458), .B2(new_n459), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n500), .B(new_n503), .C1(new_n459), .C2(new_n458), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n498), .B1(new_n502), .B2(new_n504), .ZN(G164));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(G50), .A2(new_n508), .B1(new_n514), .B2(G88), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n515), .B1(KEYINPUT68), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n520), .A2(KEYINPUT68), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n507), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n517), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n506), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n528), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n516), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT69), .B(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n507), .A2(new_n536), .B1(new_n513), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G171));
  AOI22_X1  g114(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n516), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n507), .A2(new_n542), .B1(new_n513), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n517), .A2(G65), .ZN(new_n551));
  INV_X1    g126(.A(G78), .ZN(new_n552));
  INV_X1    g127(.A(G543), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT71), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT71), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n551), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n556), .A2(G651), .B1(new_n514), .B2(G91), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n558), .B(new_n559), .C1(new_n507), .C2(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n560), .B1(KEYINPUT70), .B2(KEYINPUT9), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n508), .B(new_n562), .C1(KEYINPUT70), .C2(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n557), .A2(new_n561), .A3(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  AND2_X1   g141(.A1(new_n514), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n568));
  INV_X1    g143(.A(G49), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n569), .B2(new_n507), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G288));
  OAI21_X1  g147(.A(G61), .B1(new_n510), .B2(new_n509), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(KEYINPUT72), .B1(G73), .B2(G543), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n517), .A2(new_n575), .A3(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n516), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n517), .A2(new_n506), .A3(G86), .ZN(new_n578));
  OAI211_X1 g153(.A(G48), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n516), .ZN(new_n584));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n507), .A2(new_n585), .B1(new_n513), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n514), .A2(G92), .ZN(new_n591));
  XOR2_X1   g166(.A(KEYINPUT73), .B(KEYINPUT10), .Z(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n529), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n508), .B2(G54), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n590), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n590), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G299), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G168), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(new_n602), .B2(G168), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  INV_X1    g182(.A(new_n545), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(new_n602), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n598), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n463), .A2(new_n476), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT12), .Z(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT74), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n615), .A2(new_n616), .B1(new_n617), .B2(G2100), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n616), .B2(new_n615), .ZN(new_n619));
  OR3_X1    g194(.A1(new_n619), .A2(new_n617), .A3(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n490), .A2(G135), .ZN(new_n621));
  INV_X1    g196(.A(new_n486), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G123), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT75), .ZN(new_n625));
  INV_X1    g200(.A(G111), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n624), .A2(new_n625), .B1(new_n626), .B2(G2105), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n625), .B2(new_n624), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n621), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n619), .B1(new_n617), .B2(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(G2096), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n620), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT77), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2430), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT78), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT79), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT80), .Z(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(KEYINPUT17), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n658), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n653), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n655), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n656), .A2(new_n659), .A3(new_n653), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT81), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT20), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n669), .A2(new_n671), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n678), .A2(new_n674), .A3(new_n672), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n676), .B(new_n679), .C1(new_n674), .C2(new_n678), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT82), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1981), .B(G1986), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NOR2_X1   g263(.A1(G171), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G5), .B2(new_n688), .ZN(new_n690));
  INV_X1    g265(.A(G1961), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(KEYINPUT30), .A2(G28), .ZN(new_n693));
  NAND2_X1  g268(.A1(KEYINPUT30), .A2(G28), .ZN(new_n694));
  AOI21_X1  g269(.A(G29), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT31), .B(G11), .Z(new_n696));
  NOR3_X1   g271(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n629), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n688), .A2(G21), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G168), .B2(new_n688), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n698), .A2(G29), .B1(G1966), .B2(new_n700), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n697), .B(new_n701), .C1(G1966), .C2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT96), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G33), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n490), .A2(G139), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT25), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n706), .B(new_n709), .C1(new_n469), .C2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT93), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n705), .B1(new_n713), .B2(new_n704), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2072), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n704), .A2(G32), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n490), .A2(G141), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n622), .A2(G129), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT26), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n721), .A2(new_n722), .B1(G105), .B2(new_n476), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n717), .A2(new_n718), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n716), .B1(new_n725), .B2(new_n704), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT27), .ZN(new_n727));
  INV_X1    g302(.A(G1996), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n545), .A2(G16), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G16), .B2(G19), .ZN(new_n731));
  INV_X1    g306(.A(G1341), .ZN(new_n732));
  NOR2_X1   g307(.A1(G164), .A2(new_n704), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G27), .B2(new_n704), .ZN(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  OAI22_X1  g310(.A1(new_n731), .A2(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(new_n734), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n690), .A2(new_n691), .B1(new_n732), .B2(new_n731), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n688), .A2(G4), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n599), .B2(new_n688), .ZN(new_n741));
  INV_X1    g316(.A(G1348), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G29), .A2(G35), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G162), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n739), .B(new_n743), .C1(G2090), .C2(new_n747), .ZN(new_n748));
  NOR4_X1   g323(.A1(new_n703), .A2(new_n715), .A3(new_n729), .A4(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G34), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(KEYINPUT24), .ZN(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n750), .B2(KEYINPUT24), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(KEYINPUT94), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT94), .B2(new_n752), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n478), .B2(new_n704), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT95), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G2084), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n704), .A2(G26), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT90), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  OR2_X1    g335(.A1(G104), .A2(G2105), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n762));
  INV_X1    g337(.A(G140), .ZN(new_n763));
  INV_X1    g338(.A(G128), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n762), .B1(new_n489), .B2(new_n763), .C1(new_n764), .C2(new_n486), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT89), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n760), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT91), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n688), .A2(G20), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT23), .Z(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G299), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT98), .ZN(new_n775));
  INV_X1    g350(.A(G1956), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n747), .A2(G2090), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT99), .Z(new_n780));
  NAND4_X1  g355(.A1(new_n749), .A2(new_n757), .A3(new_n771), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G22), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G166), .B2(G16), .ZN(new_n783));
  INV_X1    g358(.A(G1971), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n688), .A2(G6), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n581), .B2(new_n688), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT32), .B(G1981), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(KEYINPUT86), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(KEYINPUT86), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n688), .A2(G23), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n571), .B2(new_n688), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT33), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1976), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n785), .A2(new_n790), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT87), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT34), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NOR2_X1   g375(.A1(G16), .A2(G24), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n588), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT85), .ZN(new_n803));
  INV_X1    g378(.A(G1986), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n704), .A2(G25), .ZN(new_n806));
  OR2_X1    g381(.A1(G95), .A2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT83), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n622), .B2(G119), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n490), .A2(G131), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n806), .B1(new_n813), .B2(new_n704), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT35), .B(G1991), .Z(new_n815));
  XOR2_X1   g390(.A(new_n814), .B(new_n815), .Z(new_n816));
  OAI21_X1  g391(.A(new_n805), .B1(new_n816), .B2(KEYINPUT84), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(KEYINPUT84), .B2(new_n816), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n799), .A2(new_n800), .A3(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT88), .B(KEYINPUT36), .Z(new_n820));
  OR2_X1    g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n781), .B1(new_n821), .B2(new_n822), .ZN(G311));
  XOR2_X1   g398(.A(G311), .B(KEYINPUT100), .Z(G150));
  NAND2_X1  g399(.A1(new_n599), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n514), .A2(G93), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n508), .A2(G55), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n827), .B(new_n828), .C1(new_n516), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n608), .B(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n826), .B(new_n831), .Z(new_n832));
  AND2_X1   g407(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n833), .A2(new_n834), .A3(G860), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(G860), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT101), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT37), .Z(new_n838));
  OR2_X1    g413(.A1(new_n835), .A2(new_n838), .ZN(G145));
  OAI21_X1  g414(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n463), .A2(new_n496), .B1(new_n841), .B2(new_n494), .ZN(new_n842));
  INV_X1    g417(.A(new_n504), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n503), .B1(new_n463), .B2(new_n500), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n767), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n724), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n711), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n846), .B(new_n725), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(new_n713), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n812), .B(new_n615), .ZN(new_n852));
  OR2_X1    g427(.A1(G106), .A2(G2105), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n854));
  INV_X1    g429(.A(G142), .ZN(new_n855));
  INV_X1    g430(.A(G130), .ZN(new_n856));
  OAI221_X1 g431(.A(new_n854), .B1(new_n489), .B2(new_n855), .C1(new_n856), .C2(new_n486), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n852), .B(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT102), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n851), .A2(new_n858), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n478), .B(new_n629), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(G162), .Z(new_n864));
  AND2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  INV_X1    g441(.A(new_n864), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n861), .B(new_n867), .C1(new_n868), .C2(new_n859), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT103), .B1(new_n851), .B2(new_n858), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n872), .A2(KEYINPUT40), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n865), .A2(new_n874), .A3(new_n871), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(new_n875), .ZN(G395));
  NOR2_X1   g451(.A1(new_n830), .A2(G868), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n571), .B(new_n588), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n878), .A2(KEYINPUT104), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(G166), .B2(G305), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(G166), .B2(G305), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(KEYINPUT104), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n881), .B(new_n882), .Z(new_n883));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(KEYINPUT105), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n831), .B(new_n610), .Z(new_n888));
  XNOR2_X1  g463(.A(new_n598), .B(G299), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(KEYINPUT41), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(new_n888), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n887), .B1(KEYINPUT106), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(KEYINPUT106), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n893), .B(new_n894), .Z(new_n895));
  AOI21_X1  g470(.A(new_n877), .B1(new_n895), .B2(G868), .ZN(G295));
  AOI21_X1  g471(.A(new_n877), .B1(new_n895), .B2(G868), .ZN(G331));
  INV_X1    g472(.A(new_n889), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n831), .B(G301), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(G168), .ZN(new_n900));
  MUX2_X1   g475(.A(new_n891), .B(new_n898), .S(new_n900), .Z(new_n901));
  AOI21_X1  g476(.A(G37), .B1(new_n901), .B2(new_n883), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n883), .B2(new_n901), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT43), .ZN(new_n904));
  NAND2_X1  g479(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n906), .B(new_n907), .Z(G397));
  XNOR2_X1  g483(.A(new_n767), .B(new_n770), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n725), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n477), .A2(G40), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI211_X1 g487(.A(KEYINPUT66), .B(new_n469), .C1(new_n470), .C2(new_n464), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n472), .B1(new_n466), .B2(G2105), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(G164), .B2(G1384), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT46), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n728), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n910), .A2(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n919), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n922), .B(KEYINPUT122), .Z(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT123), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT123), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n924), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT47), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n724), .B(new_n728), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n909), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n812), .B(new_n815), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n918), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n918), .A2(new_n804), .A3(new_n588), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT48), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n813), .A2(new_n815), .ZN(new_n939));
  OAI22_X1  g514(.A1(new_n932), .A2(new_n939), .B1(G2067), .B2(new_n767), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n936), .A2(new_n938), .B1(new_n918), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n927), .A2(new_n930), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT124), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n942), .B(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n918), .ZN(new_n945));
  INV_X1    g520(.A(new_n935), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n588), .B(G1986), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n911), .B1(new_n468), .B2(new_n473), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  NOR3_X1   g529(.A1(G164), .A2(new_n954), .A3(G1384), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT108), .B1(new_n845), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n952), .B(new_n953), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n954), .B1(G164), .B2(G1384), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n845), .A2(KEYINPUT108), .A3(new_n956), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT114), .B1(new_n963), .B2(new_n915), .ZN(new_n964));
  INV_X1    g539(.A(G2090), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n845), .A2(new_n956), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(KEYINPUT50), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n960), .A2(new_n964), .A3(new_n965), .A4(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n845), .A2(KEYINPUT45), .A3(new_n956), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n917), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n784), .B1(new_n915), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT110), .B(G8), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n951), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n974), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n961), .A2(new_n962), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(new_n915), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1976), .ZN(new_n979));
  NOR2_X1   g554(.A1(G288), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n571), .B2(G1976), .ZN(new_n982));
  OR3_X1    g557(.A1(new_n978), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT52), .B1(new_n978), .B2(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n574), .A2(new_n576), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G651), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  INV_X1    g563(.A(new_n580), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n578), .A2(new_n991), .A3(new_n579), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n578), .B2(new_n579), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n577), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT49), .B(new_n990), .C1(new_n994), .C2(new_n988), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT112), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n580), .A2(KEYINPUT111), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n578), .A2(new_n991), .A3(new_n579), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(G1981), .B1(new_n999), .B2(new_n577), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(KEYINPUT49), .A4(new_n990), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n996), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT49), .B1(new_n1000), .B2(new_n990), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n978), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT113), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1003), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n985), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n951), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n961), .A2(new_n959), .A3(new_n962), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n966), .A2(KEYINPUT50), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n953), .A2(new_n1012), .A3(new_n965), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n972), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT109), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n972), .A3(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1011), .A2(new_n1016), .A3(G8), .A4(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n975), .A2(new_n1010), .A3(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n953), .A2(new_n735), .A3(new_n917), .A4(new_n970), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(KEYINPUT118), .A3(new_n1022), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT45), .B1(new_n961), .B2(new_n962), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n970), .B(new_n912), .C1(new_n913), .C2(new_n914), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1022), .A2(G2078), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n953), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1030), .A2(new_n1031), .B1(new_n1032), .B2(new_n691), .ZN(new_n1033));
  AOI21_X1  g608(.A(G301), .B1(new_n1027), .B2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1020), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT62), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G168), .A2(new_n974), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1966), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(G2084), .B2(new_n1032), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT117), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1040), .B(new_n1043), .C1(G2084), .C2(new_n1032), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(G8), .A3(new_n1044), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(new_n1038), .ZN(new_n1048));
  AOI211_X1 g623(.A(KEYINPUT51), .B(new_n1037), .C1(new_n1041), .C2(new_n976), .ZN(new_n1049));
  OAI221_X1 g624(.A(new_n1036), .B1(new_n1038), .B2(new_n1045), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g625(.A1(new_n1048), .A2(new_n1049), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT62), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1035), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1016), .A2(G8), .A3(new_n1018), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(new_n951), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1010), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n990), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1058));
  NOR2_X1   g633(.A1(G288), .A2(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1056), .B1(new_n1060), .B2(new_n978), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1041), .A2(G168), .A3(new_n976), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n975), .A2(new_n1010), .A3(new_n1019), .A4(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(KEYINPUT63), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1054), .B2(new_n951), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1019), .A3(new_n1010), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1061), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n960), .A2(new_n964), .A3(new_n968), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n776), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT56), .B(G2072), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n953), .A2(new_n917), .A3(new_n970), .A4(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(G299), .B(KEYINPUT57), .Z(new_n1074));
  NAND3_X1  g649(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1074), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1032), .A2(new_n742), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n958), .A2(new_n953), .A3(new_n770), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(new_n599), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1076), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT61), .B1(new_n1079), .B2(new_n1075), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n963), .A2(new_n915), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n967), .B1(new_n1089), .B2(new_n952), .ZN(new_n1090));
  AOI21_X1  g665(.A(G1956), .B1(new_n1090), .B2(new_n964), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1074), .A2(new_n1073), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT61), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1074), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n608), .B1(new_n1095), .B2(KEYINPUT59), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT58), .B(G1341), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n958), .B2(new_n953), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n915), .A2(new_n971), .A3(G1996), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1095), .A2(KEYINPUT59), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1104));
  OAI22_X1  g679(.A1(new_n1093), .A2(new_n1094), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1088), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1085), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT60), .B1(new_n1107), .B2(new_n1083), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT60), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1084), .A2(new_n1109), .A3(new_n1085), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(new_n1110), .A3(new_n599), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT60), .B(new_n598), .C1(new_n1107), .C2(new_n1083), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1087), .B1(new_n1106), .B2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1021), .A2(KEYINPUT118), .A3(new_n1022), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT118), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1033), .A2(G301), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT54), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n467), .A2(new_n912), .A3(new_n1031), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n971), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1032), .B2(new_n691), .ZN(new_n1122));
  AOI21_X1  g697(.A(G301), .B1(new_n1027), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT119), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1122), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G171), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1027), .A2(G301), .A3(new_n1033), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(KEYINPUT54), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1027), .A2(G301), .A3(new_n1122), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1133), .B2(new_n1034), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1130), .A2(new_n1051), .A3(new_n1020), .A4(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1069), .B1(new_n1114), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1053), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1069), .B(KEYINPUT120), .C1(new_n1114), .C2(new_n1135), .ZN(new_n1139));
  AOI211_X1 g714(.A(KEYINPUT121), .B(new_n948), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1053), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n948), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1141), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n944), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n944), .B(KEYINPUT125), .C1(new_n1140), .C2(new_n1146), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g726(.A(G319), .ZN(new_n1153));
  OR2_X1    g727(.A1(G227), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n1155));
  AND2_X1   g729(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1157));
  NOR4_X1   g731(.A1(G229), .A2(G401), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g732(.A(new_n1158), .B(KEYINPUT127), .ZN(new_n1159));
  NAND2_X1  g733(.A1(new_n1159), .A2(new_n904), .ZN(new_n1160));
  NOR2_X1   g734(.A1(new_n1160), .A2(new_n872), .ZN(G308));
  OR2_X1    g735(.A1(new_n1160), .A2(new_n872), .ZN(G225));
endmodule


