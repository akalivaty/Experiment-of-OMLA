//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT67), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(G113), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G137), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G101), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI211_X1 g054(.A(KEYINPUT68), .B(G2105), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(G160));
  XNOR2_X1  g056(.A(KEYINPUT3), .B(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(G124), .A3(G2105), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT69), .Z(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G2104), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n485), .A2(G136), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n484), .A2(new_n490), .ZN(G162));
  AOI21_X1  g066(.A(KEYINPUT4), .B1(new_n485), .B2(G138), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G2105), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT4), .A2(G138), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n497), .B(new_n498), .C1(new_n473), .C2(new_n474), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n473), .B2(new_n474), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(new_n502), .C1(new_n473), .C2(new_n474), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(KEYINPUT71), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n496), .A2(new_n499), .ZN(new_n509));
  OAI211_X1 g084(.A(G138), .B(new_n497), .C1(new_n473), .C2(new_n474), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND4_X1   g087(.A1(KEYINPUT71), .A2(new_n507), .A3(new_n509), .A4(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n508), .A2(new_n513), .ZN(G164));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n516), .B(new_n518), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n520), .A2(new_n521), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n524), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(new_n522), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT73), .B1(new_n531), .B2(G62), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(G75), .B2(G543), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n531), .A2(KEYINPUT73), .A3(G62), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n515), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(KEYINPUT74), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n527), .B(KEYINPUT72), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n533), .A2(new_n534), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n536), .A2(new_n541), .ZN(G166));
  INV_X1    g117(.A(new_n525), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G89), .ZN(new_n544));
  AND3_X1   g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT75), .B(G51), .Z(new_n546));
  OAI221_X1 g121(.A(new_n544), .B1(KEYINPUT7), .B2(new_n545), .C1(new_n520), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n531), .A2(G63), .ZN(new_n548));
  NAND3_X1  g123(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n515), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G168));
  AOI22_X1  g126(.A1(new_n531), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n515), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n520), .A2(new_n554), .B1(new_n525), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(G171));
  AOI22_X1  g132(.A1(new_n531), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n515), .ZN(new_n559));
  INV_X1    g134(.A(G43), .ZN(new_n560));
  XOR2_X1   g135(.A(KEYINPUT76), .B(G81), .Z(new_n561));
  OAI22_X1  g136(.A1(new_n520), .A2(new_n560), .B1(new_n525), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  AND2_X1   g143(.A1(new_n543), .A2(G91), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n519), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(new_n573), .A3(G53), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n520), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(new_n531), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n571), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G299));
  INV_X1    g160(.A(G171), .ZN(G301));
  OR2_X1    g161(.A1(new_n547), .A2(new_n550), .ZN(G286));
  INV_X1    g162(.A(G166), .ZN(G303));
  NAND2_X1  g163(.A1(new_n572), .A2(G49), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n543), .A2(G87), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n531), .B2(G74), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G288));
  NAND4_X1  g168(.A1(new_n516), .A2(new_n518), .A3(G48), .A4(G543), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n525), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT78), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n530), .B2(new_n522), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n597), .A2(new_n602), .ZN(G305));
  NAND2_X1  g178(.A1(G72), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G60), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n579), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n515), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(new_n606), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n572), .A2(G47), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n543), .A2(G85), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n525), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n579), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n619), .A2(G651), .B1(new_n572), .B2(G54), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n613), .B1(new_n622), .B2(G868), .ZN(G284));
  OAI21_X1  g198(.A(new_n613), .B1(new_n622), .B2(G868), .ZN(G321));
  NAND3_X1  g199(.A1(G286), .A2(KEYINPUT80), .A3(G868), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT80), .ZN(new_n626));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(G168), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n628), .C1(G868), .C2(new_n584), .ZN(G297));
  OAI211_X1 g204(.A(new_n625), .B(new_n628), .C1(G868), .C2(new_n584), .ZN(G280));
  XNOR2_X1  g205(.A(KEYINPUT81), .B(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n622), .B1(G860), .B2(new_n631), .ZN(G148));
  NAND2_X1  g207(.A1(new_n622), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n485), .A2(G2104), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT13), .Z(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n485), .A2(G135), .ZN(new_n643));
  NOR2_X1   g218(.A1(G99), .A2(G2105), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(new_n497), .B2(G111), .ZN(new_n645));
  INV_X1    g220(.A(G123), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n482), .A2(G2105), .ZN(new_n647));
  OAI221_X1 g222(.A(new_n643), .B1(new_n644), .B2(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2096), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n641), .A2(new_n642), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2443), .B(G2446), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT83), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(G14), .B1(new_n656), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n656), .ZN(G401));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n668), .B(KEYINPUT85), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT17), .ZN(new_n672));
  INV_X1    g247(.A(new_n666), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n672), .A2(new_n667), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n667), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n673), .B1(new_n667), .B2(new_n668), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT84), .Z(new_n677));
  AOI211_X1 g252(.A(new_n670), .B(new_n674), .C1(new_n675), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2096), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2100), .ZN(G227));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT86), .ZN(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n688), .B(new_n691), .C1(new_n682), .C2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT87), .ZN(new_n697));
  INV_X1    g272(.A(G1981), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n695), .B(new_n699), .ZN(G229));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n701), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(G1971), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(G1971), .ZN(new_n705));
  MUX2_X1   g280(.A(G6), .B(G305), .S(G16), .Z(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G23), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT88), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G288), .B2(new_n701), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n704), .A2(new_n705), .A3(new_n708), .A4(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n716));
  OR2_X1    g291(.A1(G16), .A2(G24), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G290), .B2(new_n701), .ZN(new_n718));
  INV_X1    g293(.A(G1986), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n485), .A2(G131), .ZN(new_n722));
  NOR2_X1   g297(.A1(G95), .A2(G2105), .ZN(new_n723));
  OAI21_X1  g298(.A(G2104), .B1(new_n497), .B2(G107), .ZN(new_n724));
  INV_X1    g299(.A(G119), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n722), .B1(new_n723), .B2(new_n724), .C1(new_n725), .C2(new_n647), .ZN(new_n726));
  MUX2_X1   g301(.A(G25), .B(new_n726), .S(G29), .Z(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n727), .B(new_n729), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n720), .A2(new_n721), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n715), .A2(new_n716), .A3(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT36), .Z(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G27), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G164), .B2(new_n734), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G2078), .ZN(new_n737));
  INV_X1    g312(.A(G28), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT30), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n738), .B2(KEYINPUT30), .ZN(new_n740));
  OR2_X1    g315(.A1(KEYINPUT31), .A2(G11), .ZN(new_n741));
  NAND2_X1  g316(.A1(KEYINPUT31), .A2(G11), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n739), .A2(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AND3_X1   g318(.A1(new_n497), .A2(G103), .A3(G2104), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT25), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n485), .A2(G139), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n497), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(new_n734), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n734), .B2(G33), .ZN(new_n752));
  INV_X1    g327(.A(G2072), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n743), .B1(new_n734), .B2(new_n648), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n701), .A2(G19), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n563), .B2(new_n701), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1341), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT91), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n734), .A2(G26), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n760), .B(new_n761), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n485), .A2(G140), .ZN(new_n763));
  NOR2_X1   g338(.A1(G104), .A2(G2105), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(new_n497), .B2(G116), .ZN(new_n765));
  INV_X1    g340(.A(G128), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n763), .B1(new_n764), .B2(new_n765), .C1(new_n766), .C2(new_n647), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n762), .B1(G29), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2067), .ZN(new_n769));
  NOR2_X1   g344(.A1(G168), .A2(new_n701), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n701), .B2(G21), .ZN(new_n771));
  INV_X1    g346(.A(G1966), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n758), .A2(new_n769), .A3(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G1961), .ZN(new_n775));
  NOR2_X1   g350(.A1(G171), .A2(new_n701), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G5), .B2(new_n701), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n775), .A2(new_n777), .B1(new_n752), .B2(new_n753), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n734), .A2(G32), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT26), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  AND2_X1   g358(.A1(G105), .A2(G2104), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n782), .A2(new_n783), .B1(new_n497), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n485), .A2(G141), .ZN(new_n786));
  INV_X1    g361(.A(G129), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n785), .B(new_n786), .C1(new_n787), .C2(new_n647), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT92), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n779), .B1(new_n789), .B2(G29), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT27), .B(G1996), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT93), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT24), .ZN(new_n795));
  INV_X1    g370(.A(G34), .ZN(new_n796));
  AOI21_X1  g371(.A(G29), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G160), .B2(new_n734), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G2084), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n777), .A2(new_n775), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n778), .A2(new_n794), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n734), .A2(G35), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G162), .B2(new_n734), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT29), .B(G2090), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n772), .B2(new_n771), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n774), .A2(new_n802), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n701), .A2(G20), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT96), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT23), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n584), .B2(new_n701), .ZN(new_n812));
  INV_X1    g387(.A(G1956), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n736), .A2(G2078), .ZN(new_n815));
  AND4_X1   g390(.A1(new_n737), .A2(new_n808), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n701), .A2(G4), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n622), .B2(new_n701), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT89), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G1348), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n799), .A2(G2084), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT95), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n791), .A2(new_n793), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT94), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n816), .A2(new_n820), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n733), .A2(new_n825), .ZN(G311));
  INV_X1    g401(.A(G311), .ZN(G150));
  AOI22_X1  g402(.A1(new_n531), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n515), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n520), .A2(new_n830), .B1(new_n525), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G860), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT98), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT37), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n563), .A2(new_n833), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n563), .A2(new_n833), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n622), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT97), .Z(new_n846));
  OAI21_X1  g421(.A(new_n834), .B1(new_n843), .B2(new_n844), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n837), .B1(new_n846), .B2(new_n847), .ZN(G145));
  NAND2_X1  g423(.A1(new_n501), .A2(new_n507), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n750), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n789), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n767), .ZN(new_n852));
  INV_X1    g427(.A(G130), .ZN(new_n853));
  NOR2_X1   g428(.A1(G106), .A2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(new_n497), .B2(G118), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n647), .A2(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(G142), .B2(new_n485), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(new_n726), .Z(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(new_n639), .Z(new_n859));
  OR2_X1    g434(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n852), .A2(new_n859), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(G160), .B(new_n648), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT99), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G162), .ZN(new_n865));
  AOI21_X1  g440(.A(G37), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n860), .A2(new_n861), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n852), .A2(KEYINPUT100), .A3(new_n859), .ZN(new_n869));
  INV_X1    g444(.A(new_n865), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n868), .A2(KEYINPUT101), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT101), .B1(new_n868), .B2(new_n871), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n866), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n876));
  NAND2_X1  g451(.A1(G166), .A2(new_n592), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n536), .A2(new_n541), .A3(G288), .ZN(new_n878));
  XNOR2_X1  g453(.A(G290), .B(G305), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n877), .B2(new_n878), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT42), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n840), .B(new_n633), .Z(new_n889));
  INV_X1    g464(.A(new_n571), .ZN(new_n890));
  INV_X1    g465(.A(new_n583), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n621), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n622), .B1(new_n583), .B2(new_n571), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n894), .B(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n889), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n887), .B1(new_n888), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n888), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT102), .B1(new_n896), .B2(new_n899), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n884), .B(new_n886), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(G868), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n833), .A2(G868), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n876), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AOI211_X1 g484(.A(KEYINPUT103), .B(new_n907), .C1(new_n905), .C2(G868), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(G295));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n908), .ZN(G331));
  NAND2_X1  g487(.A1(G286), .A2(G171), .ZN(new_n913));
  NAND2_X1  g488(.A1(G168), .A2(G301), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n840), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n913), .A2(new_n838), .A3(new_n839), .A4(new_n914), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n894), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n894), .B(KEYINPUT41), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n920), .A2(KEYINPUT104), .A3(new_n918), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  INV_X1    g497(.A(new_n918), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n922), .B1(new_n898), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n882), .B(new_n919), .C1(new_n921), .C2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  INV_X1    g502(.A(new_n919), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT104), .B1(new_n920), .B2(new_n918), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n898), .A2(new_n923), .A3(new_n922), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n927), .B1(new_n931), .B2(new_n882), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n926), .B1(new_n932), .B2(KEYINPUT105), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n934), .B(new_n927), .C1(new_n931), .C2(new_n882), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT43), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n919), .B1(new_n920), .B2(new_n918), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n883), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n883), .A2(KEYINPUT106), .A3(new_n937), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n940), .A2(new_n927), .A3(new_n925), .A4(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT44), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n943), .B1(new_n933), .B2(new_n935), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n949), .ZN(G397));
  INV_X1    g525(.A(KEYINPUT117), .ZN(new_n951));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n508), .B2(new_n513), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(KEYINPUT107), .A3(KEYINPUT50), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT71), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n512), .A2(new_n499), .A3(new_n496), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n505), .B1(new_n482), .B2(new_n502), .ZN(new_n958));
  INV_X1    g533(.A(new_n506), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT71), .A4(new_n512), .ZN(new_n962));
  AOI21_X1  g537(.A(G1384), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n955), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n954), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  AOI21_X1  g542(.A(G1384), .B1(new_n501), .B2(new_n507), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n964), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n482), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT68), .B1(new_n970), .B2(G2105), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n477), .A2(new_n478), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(new_n972), .A3(G40), .A4(new_n472), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G2090), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n966), .A2(new_n967), .A3(new_n969), .A4(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G40), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n479), .A2(new_n976), .A3(new_n480), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n968), .A2(KEYINPUT45), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n977), .B(new_n978), .C1(new_n963), .C2(KEYINPUT45), .ZN(new_n979));
  INV_X1    g554(.A(G1971), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n954), .A2(new_n965), .B1(new_n964), .B2(new_n968), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n967), .B1(new_n983), .B2(new_n974), .ZN(new_n984));
  OAI21_X1  g559(.A(G8), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n536), .A2(G8), .A3(new_n541), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT55), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n986), .B(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(G8), .B(new_n990), .C1(new_n982), .C2(new_n984), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n589), .A2(new_n590), .A3(G1976), .A4(new_n591), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n952), .B1(new_n957), .B2(new_n960), .ZN(new_n993));
  OAI211_X1 g568(.A(G8), .B(new_n992), .C1(new_n973), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n592), .B2(G1976), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT110), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n994), .B2(new_n996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n1002));
  INV_X1    g577(.A(new_n994), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n995), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n994), .A2(KEYINPUT109), .A3(KEYINPUT52), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G8), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n977), .B2(new_n968), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n519), .A2(new_n531), .A3(G86), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n602), .A2(new_n698), .A3(new_n1010), .A4(new_n594), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT111), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n597), .A2(new_n1013), .A3(new_n698), .A4(new_n602), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1012), .A2(new_n1014), .B1(G1981), .B2(G305), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1009), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G305), .A2(G1981), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1018), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1008), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n1022));
  AND4_X1   g597(.A1(new_n1022), .A2(new_n1018), .A3(KEYINPUT49), .A4(new_n1019), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1015), .B2(KEYINPUT49), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1001), .B(new_n1006), .C1(new_n1021), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1029), .B(G1384), .C1(new_n961), .C2(new_n962), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n993), .A2(new_n1029), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n977), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n772), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT116), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n973), .B1(new_n1029), .B2(new_n993), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n953), .B2(new_n1029), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n772), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G2084), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n966), .A2(new_n1040), .A3(new_n977), .A4(new_n969), .ZN(new_n1041));
  AOI211_X1 g616(.A(new_n1007), .B(G286), .C1(new_n1039), .C2(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n991), .A2(new_n1028), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n981), .ZN(new_n1044));
  NOR2_X1   g619(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n508), .B2(new_n513), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(KEYINPUT114), .B(new_n1045), .C1(new_n508), .C2(new_n513), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n973), .B1(KEYINPUT50), .B2(new_n993), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G2090), .B1(new_n1051), .B2(KEYINPUT115), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1048), .A2(new_n1053), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1044), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n987), .B1(new_n1055), .B2(new_n1007), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1026), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1056), .A2(new_n991), .A3(new_n1042), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n988), .A2(new_n1043), .B1(new_n1058), .B2(new_n1027), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n991), .A2(new_n1026), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1061), .A2(G1976), .A3(G288), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1018), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1008), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n951), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1058), .A2(new_n1027), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n988), .A2(new_n991), .A3(new_n1042), .A4(new_n1028), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1065), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(KEYINPUT117), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n584), .B(KEYINPUT57), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1051), .A2(new_n813), .ZN(new_n1073));
  INV_X1    g648(.A(new_n979), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1072), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1348), .B1(new_n983), .B2(new_n977), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n977), .A2(new_n1079), .A3(new_n968), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT118), .B1(new_n973), .B2(new_n993), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G2067), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT119), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(new_n1086), .A3(new_n1083), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n622), .B1(new_n1078), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1072), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1077), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT58), .B(G1341), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n979), .A2(G1996), .B1(new_n1082), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n563), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(KEYINPUT121), .A3(new_n563), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(KEYINPUT59), .A3(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1104));
  NAND3_X1  g679(.A1(new_n1098), .A2(new_n563), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1073), .A2(new_n1076), .A3(new_n1072), .A4(KEYINPUT61), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1103), .A2(new_n1105), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n966), .A2(new_n977), .A3(new_n969), .ZN(new_n1111));
  INV_X1    g686(.A(G1348), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(new_n621), .B(KEYINPUT123), .Z(new_n1114));
  NAND4_X1  g689(.A1(new_n1110), .A2(new_n1113), .A3(KEYINPUT60), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n1078), .B2(new_n1088), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1078), .A2(new_n1088), .A3(new_n1116), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n621), .A2(KEYINPUT123), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1115), .B(new_n1117), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1109), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1096), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1111), .A2(new_n775), .ZN(new_n1123));
  INV_X1    g698(.A(G2078), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT53), .B1(new_n1074), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(KEYINPUT53), .A3(new_n1124), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1123), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G301), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1125), .B1(new_n775), .B2(new_n1111), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1035), .A2(KEYINPUT53), .A3(new_n1124), .A4(new_n978), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(G171), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1130), .A2(new_n1133), .A3(KEYINPUT54), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT54), .B1(new_n1129), .B2(G171), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1123), .A2(new_n1126), .A3(G301), .A4(new_n1132), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1134), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(G168), .A2(new_n1007), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT124), .ZN(new_n1143));
  NAND2_X1  g718(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(new_n1041), .A3(new_n1039), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1007), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1143), .B1(new_n1147), .B2(new_n1144), .ZN(new_n1148));
  AOI211_X1 g723(.A(KEYINPUT51), .B(new_n1007), .C1(new_n1039), .C2(new_n1041), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1056), .A2(new_n991), .A3(new_n1057), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1122), .A2(new_n1141), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1151), .ZN(new_n1156));
  AOI21_X1  g731(.A(G301), .B1(new_n1131), .B2(new_n1128), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1146), .B(KEYINPUT62), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1066), .A2(new_n1071), .A3(new_n1153), .A4(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1031), .A2(new_n973), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n789), .B(G1996), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n767), .B(new_n1083), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n726), .B(new_n728), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(G290), .B(G1986), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1161), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1160), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1161), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n726), .A2(new_n729), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1165), .A2(new_n1172), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n767), .A2(G2067), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1167), .A2(new_n1161), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1171), .A2(G1986), .A3(G290), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1177), .B(KEYINPUT48), .Z(new_n1178));
  AOI21_X1  g753(.A(new_n1175), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT47), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT46), .ZN(new_n1181));
  OR3_X1    g756(.A1(new_n1171), .A2(new_n1181), .A3(G1996), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1161), .B1(new_n1164), .B2(new_n789), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1181), .B1(new_n1171), .B2(G1996), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT127), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1179), .B1(new_n1180), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1180), .B2(new_n1186), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1170), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g764(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1191));
  OAI211_X1 g765(.A(new_n874), .B(new_n1191), .C1(new_n947), .C2(new_n948), .ZN(G225));
  INV_X1    g766(.A(G225), .ZN(G308));
endmodule


