//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT89), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n204), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n205), .A2(new_n206), .B1(KEYINPUT16), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n203), .B(KEYINPUT89), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(new_n207), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n209), .B(new_n211), .C1(KEYINPUT90), .C2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n208), .B1(new_n207), .B2(new_n210), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT90), .ZN(new_n216));
  OAI21_X1  g015(.A(G8gat), .B1(new_n208), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n202), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n217), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n209), .A2(new_n211), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(KEYINPUT91), .A3(new_n213), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT95), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G57gat), .ZN(new_n228));
  INV_X1    g027(.A(G64gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n225), .A2(new_n226), .ZN(new_n231));
  NAND2_X1  g030(.A1(G57gat), .A2(G64gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n227), .A2(new_n230), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(G71gat), .B(G78gat), .Z(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n225), .B(KEYINPUT95), .ZN(new_n236));
  INV_X1    g035(.A(new_n234), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n229), .B1(new_n228), .B2(KEYINPUT96), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n232), .A2(KEYINPUT96), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT97), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT97), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n235), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT21), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n224), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G183gat), .ZN(new_n248));
  AND2_X1   g047(.A1(G231gat), .A2(G233gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G127gat), .B(G155gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G211gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n250), .B(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n245), .A2(KEYINPUT21), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n250), .A2(new_n252), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n250), .A2(new_n252), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n256), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT85), .ZN(new_n265));
  NOR2_X1   g064(.A1(KEYINPUT82), .A2(KEYINPUT14), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G29gat), .ZN(new_n268));
  INV_X1    g067(.A(G36gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(KEYINPUT82), .A2(KEYINPUT14), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n267), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(KEYINPUT82), .A2(KEYINPUT14), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(new_n268), .A3(new_n269), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(KEYINPUT83), .A2(G36gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(KEYINPUT83), .A2(G36gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(G29gat), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT84), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g079(.A1(KEYINPUT83), .A2(G36gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(KEYINPUT83), .A2(G36gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(KEYINPUT84), .A3(G29gat), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n275), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G43gat), .B(G50gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT15), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n265), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n271), .A2(G29gat), .A3(G36gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n266), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n270), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT84), .B1(new_n283), .B2(G29gat), .ZN(new_n292));
  NOR4_X1   g091(.A1(new_n281), .A2(new_n282), .A3(new_n279), .A4(new_n268), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n287), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT85), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n286), .A2(KEYINPUT15), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n285), .A2(new_n287), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT86), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n284), .ZN(new_n301));
  AOI211_X1 g100(.A(new_n265), .B(new_n287), .C1(new_n301), .C2(new_n291), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT85), .B1(new_n294), .B2(new_n295), .ZN(new_n303));
  OAI211_X1 g102(.A(KEYINPUT86), .B(new_n299), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n264), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT88), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT86), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n304), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT88), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(new_n264), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G99gat), .B(G106gat), .Z(new_n315));
  INV_X1    g114(.A(KEYINPUT99), .ZN(new_n316));
  INV_X1    g115(.A(G85gat), .ZN(new_n317));
  INV_X1    g116(.A(G92gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(KEYINPUT7), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT7), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n316), .B(new_n322), .C1(new_n317), .C2(new_n318), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G99gat), .A2(G106gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT8), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT100), .B(G85gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(G92gat), .ZN(new_n328));
  OAI211_X1 g127(.A(KEYINPUT101), .B(new_n315), .C1(new_n324), .C2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  INV_X1    g129(.A(new_n315), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n330), .A2(new_n331), .A3(new_n323), .A4(new_n321), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n315), .B1(new_n324), .B2(new_n328), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT101), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n297), .A2(KEYINPUT17), .A3(new_n299), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n314), .A2(new_n329), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G134gat), .B(G162gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(new_n329), .ZN(new_n340));
  NAND2_X1  g139(.A1(G232gat), .A2(G233gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n341), .B(KEYINPUT98), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n311), .A2(new_n340), .B1(KEYINPUT41), .B2(new_n343), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n337), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n339), .B1(new_n337), .B2(new_n344), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n343), .A2(KEYINPUT41), .ZN(new_n347));
  XNOR2_X1  g146(.A(G190gat), .B(G218gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT102), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n347), .B(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  OR3_X1    g150(.A1(new_n345), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n345), .B2(new_n346), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n262), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n332), .A2(new_n333), .A3(new_n235), .A4(new_n240), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n356), .B(new_n357), .C1(new_n245), .C2(new_n340), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n245), .A2(new_n340), .A3(KEYINPUT10), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(new_n359), .B1(G230gat), .B2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n357), .B1(new_n245), .B2(new_n340), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(G230gat), .A3(G233gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(G176gat), .B(G204gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(G148gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT103), .ZN(new_n366));
  INV_X1    g165(.A(G120gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n361), .A2(new_n363), .A3(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT104), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n361), .A2(new_n363), .ZN(new_n371));
  INV_X1    g170(.A(new_n368), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n355), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT11), .B(G169gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(G197gat), .ZN(new_n377));
  XOR2_X1   g176(.A(G113gat), .B(G141gat), .Z(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT12), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n224), .B1(new_n310), .B2(new_n304), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n336), .A2(new_n213), .A3(new_n222), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n384), .B1(new_n314), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G229gat), .A2(G233gat), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n312), .B1(new_n311), .B2(new_n264), .ZN(new_n389));
  AOI211_X1 g188(.A(KEYINPUT88), .B(new_n263), .C1(new_n310), .C2(new_n304), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n224), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n311), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n391), .A2(KEYINPUT18), .A3(new_n387), .A4(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n387), .B(KEYINPUT13), .Z(new_n395));
  NOR2_X1   g194(.A1(new_n392), .A2(new_n311), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(new_n384), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n381), .B1(new_n388), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT93), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n391), .A2(new_n387), .A3(new_n393), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n382), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n402), .A2(new_n380), .A3(new_n394), .A4(new_n397), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(KEYINPUT93), .B(new_n381), .C1(new_n388), .C2(new_n398), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n404), .A2(KEYINPUT94), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT94), .B1(new_n404), .B2(new_n405), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(G155gat), .B(G162gat), .Z(new_n409));
  XOR2_X1   g208(.A(KEYINPUT73), .B(KEYINPUT2), .Z(new_n410));
  XNOR2_X1  g209(.A(G141gat), .B(G148gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT74), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  NAND2_X1  g214(.A1(G155gat), .A2(G162gat), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n409), .B1(KEYINPUT2), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G141gat), .ZN(new_n418));
  OR3_X1    g217(.A1(new_n418), .A2(KEYINPUT75), .A3(G148gat), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT75), .B1(new_n418), .B2(G148gat), .ZN(new_n420));
  INV_X1    g219(.A(G148gat), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n419), .B(new_n420), .C1(G141gat), .C2(new_n421), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n414), .A2(new_n415), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT3), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G197gat), .B(G204gat), .ZN(new_n426));
  INV_X1    g225(.A(G211gat), .ZN(new_n427));
  INV_X1    g226(.A(G218gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n426), .B1(KEYINPUT22), .B2(new_n429), .ZN(new_n430));
  XOR2_X1   g229(.A(G211gat), .B(G218gat), .Z(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT71), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n425), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT29), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n423), .B1(new_n424), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(G50gat), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n438), .ZN(new_n440));
  INV_X1    g239(.A(G50gat), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n440), .B(new_n441), .C1(new_n425), .C2(new_n434), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT31), .B(G22gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(G228gat), .A2(G233gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G78gat), .B(G106gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n446), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n439), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n448), .B1(new_n447), .B2(new_n450), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n412), .B(new_n413), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n417), .A2(new_n422), .ZN(new_n456));
  XNOR2_X1  g255(.A(G127gat), .B(G134gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(KEYINPUT68), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT67), .B(G120gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(G113gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n367), .A2(G113gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT1), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT1), .ZN(new_n464));
  INV_X1    g263(.A(G113gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(G120gat), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(G127gat), .A2(G134gat), .ZN(new_n468));
  XOR2_X1   g267(.A(KEYINPUT66), .B(G127gat), .Z(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(G134gat), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n458), .A2(new_n463), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT4), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n456), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n423), .A2(new_n424), .ZN(new_n476));
  INV_X1    g275(.A(new_n471), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G225gat), .A2(G233gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(KEYINPUT5), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n473), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n472), .A2(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT76), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT77), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n472), .B2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n423), .A2(KEYINPUT77), .A3(new_n487), .A4(new_n471), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT76), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n489), .A3(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n484), .A2(new_n486), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(new_n479), .A3(new_n478), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT5), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n477), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n472), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n493), .B1(new_n495), .B2(new_n480), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n482), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  XOR2_X1   g296(.A(G1gat), .B(G29gat), .Z(new_n498));
  XNOR2_X1  g297(.A(G57gat), .B(G85gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  NOR2_X1   g301(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n479), .B1(new_n473), .B2(new_n478), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n495), .A2(new_n480), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT39), .ZN(new_n507));
  INV_X1    g306(.A(new_n502), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT39), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n503), .B1(new_n511), .B2(KEYINPUT40), .ZN(new_n512));
  XNOR2_X1  g311(.A(G8gat), .B(G36gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(new_n229), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(new_n318), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G183gat), .A2(G190gat), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n517), .A2(KEYINPUT24), .ZN(new_n518));
  OR2_X1    g317(.A1(G183gat), .A2(G190gat), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n518), .A2(new_n519), .B1(G169gat), .B2(G176gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(G169gat), .A2(G176gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT23), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n520), .B(new_n523), .C1(KEYINPUT24), .C2(new_n517), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT25), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G183gat), .ZN(new_n527));
  INV_X1    g326(.A(G190gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(KEYINPUT28), .Z(new_n530));
  INV_X1    g329(.A(KEYINPUT64), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT26), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n521), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G169gat), .A2(G176gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n521), .A2(new_n532), .ZN(new_n535));
  OAI211_X1 g334(.A(KEYINPUT64), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n538), .A2(KEYINPUT65), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(KEYINPUT65), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n530), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G226gat), .A2(G233gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n436), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n543), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n526), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n544), .A2(new_n434), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n434), .B1(new_n544), .B2(new_n546), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n516), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT72), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT72), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n552), .B(new_n516), .C1(new_n547), .C2(new_n548), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n434), .ZN(new_n555));
  AOI211_X1 g354(.A(KEYINPUT29), .B(new_n545), .C1(new_n526), .C2(new_n541), .ZN(new_n556));
  INV_X1    g355(.A(new_n546), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n544), .A2(new_n434), .A3(new_n546), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n515), .A3(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n549), .A2(new_n551), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n554), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n512), .B(new_n562), .C1(KEYINPUT40), .C2(new_n511), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT38), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT81), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT37), .B1(new_n547), .B2(new_n548), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT37), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n558), .A2(new_n567), .A3(new_n559), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n565), .B1(new_n569), .B2(new_n515), .ZN(new_n570));
  AOI211_X1 g369(.A(KEYINPUT81), .B(new_n516), .C1(new_n566), .C2(new_n568), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n564), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT80), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n492), .A2(new_n496), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n508), .B1(new_n574), .B2(new_n482), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT6), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n503), .A2(KEYINPUT80), .A3(KEYINPUT6), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n497), .A2(new_n502), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n572), .A2(new_n577), .A3(new_n578), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n569), .A2(new_n515), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT81), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n569), .A2(new_n565), .A3(new_n515), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(KEYINPUT38), .A3(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n550), .A2(new_n553), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n454), .B(new_n563), .C1(new_n581), .C2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT32), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT69), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(new_n542), .B2(new_n477), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n542), .A2(new_n477), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n526), .A2(new_n541), .A3(KEYINPUT69), .A4(new_n471), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G227gat), .A2(G233gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n589), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n591), .A2(new_n592), .A3(new_n595), .A4(new_n593), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(KEYINPUT34), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(KEYINPUT34), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n594), .A2(new_n596), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G71gat), .B(G99gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT70), .ZN(new_n608));
  XNOR2_X1  g407(.A(G15gat), .B(G43gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n602), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n597), .B1(new_n612), .B2(new_n600), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n603), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n611), .B1(new_n613), .B2(new_n603), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT36), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n614), .B2(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT79), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n575), .A2(new_n622), .A3(new_n576), .A4(new_n579), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n577), .A2(new_n578), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n562), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n588), .B(new_n620), .C1(new_n626), .C2(new_n454), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT35), .ZN(new_n628));
  NOR4_X1   g427(.A1(new_n614), .A2(new_n615), .A3(new_n453), .A4(new_n628), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n614), .A2(new_n615), .A3(new_n453), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n631));
  INV_X1    g430(.A(new_n562), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n626), .A2(new_n629), .B1(new_n633), .B2(new_n628), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n408), .B1(new_n627), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n375), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n624), .A2(new_n625), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(new_n207), .ZN(G1324gat));
  NOR2_X1   g438(.A1(new_n636), .A2(new_n632), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT42), .Z(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n212), .B2(new_n640), .ZN(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n636), .A2(new_n645), .A3(new_n620), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n375), .A2(new_n635), .A3(new_n616), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n645), .B2(new_n647), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n636), .A2(new_n454), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT43), .B(G22gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  NAND2_X1  g450(.A1(new_n627), .A2(new_n634), .ZN(new_n652));
  INV_X1    g451(.A(new_n354), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n408), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n262), .A2(new_n374), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n637), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n268), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT45), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n354), .B1(new_n627), .B2(new_n634), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(KEYINPUT44), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664));
  AOI211_X1 g463(.A(new_n664), .B(new_n354), .C1(new_n627), .C2(new_n634), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n404), .A2(new_n405), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n668), .A3(new_n656), .ZN(new_n669));
  OAI21_X1  g468(.A(G29gat), .B1(new_n669), .B2(new_n637), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n661), .A2(new_n670), .ZN(G1328gat));
  NOR3_X1   g470(.A1(new_n657), .A2(new_n283), .A3(new_n632), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT46), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n283), .B1(new_n669), .B2(new_n632), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(G1329gat));
  INV_X1    g474(.A(new_n616), .ZN(new_n676));
  OR3_X1    g475(.A1(new_n657), .A2(G43gat), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT105), .ZN(new_n678));
  OAI21_X1  g477(.A(G43gat), .B1(new_n669), .B2(new_n620), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT47), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n678), .A2(KEYINPUT47), .A3(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(G1330gat));
  OAI21_X1  g483(.A(new_n441), .B1(new_n657), .B2(new_n454), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n669), .A2(new_n441), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n686), .B2(new_n454), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g487(.A1(new_n355), .A2(new_n668), .ZN(new_n689));
  INV_X1    g488(.A(new_n374), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n627), .B2(new_n634), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n637), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n228), .ZN(G1332gat));
  NOR2_X1   g493(.A1(new_n692), .A2(new_n632), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT49), .B(G64gat), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n695), .B2(new_n698), .ZN(G1333gat));
  INV_X1    g498(.A(new_n620), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n689), .A2(new_n691), .A3(G71gat), .A4(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n692), .A2(new_n676), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(G71gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g503(.A1(new_n692), .A2(new_n454), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(G78gat), .Z(G1335gat));
  INV_X1    g505(.A(new_n262), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(KEYINPUT106), .A3(new_n667), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n262), .B2(new_n668), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT51), .B1(new_n711), .B2(new_n662), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n662), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT109), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n714), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n716), .A2(new_n712), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  OR4_X1    g518(.A1(new_n637), .A2(new_n719), .A3(new_n327), .A4(new_n690), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n654), .A2(new_n664), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n662), .A2(KEYINPUT44), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n722), .A2(new_n374), .A3(new_n723), .A4(new_n711), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT107), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n666), .A2(new_n726), .A3(new_n374), .A4(new_n711), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n721), .B1(new_n729), .B2(new_n637), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(KEYINPUT108), .A3(new_n659), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n327), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n720), .A2(new_n732), .ZN(G1336gat));
  NOR3_X1   g532(.A1(new_n663), .A2(new_n665), .A3(new_n690), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n726), .B1(new_n734), .B2(new_n711), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n724), .A2(KEYINPUT107), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n562), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(KEYINPUT110), .A3(G92gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n632), .B1(new_n725), .B2(new_n727), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(new_n318), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n690), .B1(new_n713), .B2(new_n714), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(new_n318), .A3(new_n562), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT52), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746));
  OAI21_X1  g545(.A(G92gat), .B1(new_n724), .B2(new_n632), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n743), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(G1337gat));
  OAI21_X1  g548(.A(G99gat), .B1(new_n729), .B2(new_n620), .ZN(new_n750));
  INV_X1    g549(.A(G99gat), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n374), .C1(new_n715), .C2(new_n718), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n752), .B2(new_n676), .ZN(G1338gat));
  INV_X1    g552(.A(G106gat), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(new_n728), .B2(new_n453), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n374), .B(new_n453), .C1(new_n716), .C2(new_n712), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(G106gat), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT53), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT111), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n760), .B(KEYINPUT53), .C1(new_n755), .C2(new_n757), .ZN(new_n761));
  OR3_X1    g560(.A1(new_n756), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n734), .A2(new_n453), .A3(new_n711), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT53), .B1(new_n763), .B2(G106gat), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT112), .B1(new_n756), .B2(G106gat), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n759), .A2(new_n761), .A3(new_n766), .ZN(G1339gat));
  NAND2_X1  g566(.A1(new_n659), .A2(new_n632), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n358), .A2(new_n359), .ZN(new_n769));
  NAND2_X1  g568(.A1(G230gat), .A2(G233gat), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(KEYINPUT54), .A3(new_n361), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n773), .A3(new_n770), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n774), .A2(KEYINPUT113), .A3(new_n372), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT113), .B1(new_n774), .B2(new_n372), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g578(.A(KEYINPUT55), .B(new_n772), .C1(new_n775), .C2(new_n776), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n370), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT114), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n779), .A2(new_n783), .A3(new_n370), .A4(new_n780), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n404), .A2(new_n782), .A3(new_n405), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n386), .A2(new_n387), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n396), .A2(new_n384), .A3(new_n395), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n379), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(new_n374), .A3(new_n403), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n785), .A2(KEYINPUT116), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT116), .B1(new_n785), .B2(new_n789), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n790), .A2(new_n791), .A3(new_n653), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n403), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT115), .Z(new_n794));
  AND2_X1   g593(.A1(new_n782), .A2(new_n784), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n653), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n707), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n355), .A2(new_n374), .A3(new_n668), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n768), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n630), .ZN(new_n802));
  OAI21_X1  g601(.A(G113gat), .B1(new_n802), .B2(new_n408), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n801), .A2(new_n465), .A3(new_n668), .A4(new_n630), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1340gat));
  NOR2_X1   g604(.A1(new_n802), .A2(new_n690), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n459), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n367), .B2(new_n806), .ZN(G1341gat));
  NOR2_X1   g607(.A1(new_n802), .A2(new_n707), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n469), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n469), .A2(new_n810), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n809), .B2(new_n811), .ZN(G1342gat));
  NOR2_X1   g613(.A1(new_n802), .A2(new_n354), .ZN(new_n815));
  INV_X1    g614(.A(G134gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n817), .A2(KEYINPUT56), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(KEYINPUT56), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n818), .B(new_n819), .C1(new_n816), .C2(new_n815), .ZN(G1343gat));
  AOI21_X1  g619(.A(new_n454), .B1(new_n798), .B2(new_n800), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT118), .B1(new_n821), .B2(KEYINPUT57), .ZN(new_n822));
  INV_X1    g621(.A(new_n781), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n406), .B2(new_n407), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n789), .B(KEYINPUT119), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n653), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT120), .B(new_n707), .C1(new_n827), .C2(new_n797), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n800), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT94), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n667), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n404), .A2(KEYINPUT94), .A3(new_n405), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n781), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n354), .B1(new_n833), .B2(new_n825), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n796), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT120), .B1(new_n835), .B2(new_n707), .ZN(new_n836));
  OAI211_X1 g635(.A(KEYINPUT57), .B(new_n453), .C1(new_n829), .C2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n791), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n785), .A2(KEYINPUT116), .A3(new_n789), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n354), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n262), .B1(new_n840), .B2(new_n796), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n453), .B1(new_n841), .B2(new_n799), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n822), .A2(new_n837), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n408), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n768), .A2(new_n700), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(G141gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n821), .A2(new_n848), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n851), .A2(G141gat), .A3(new_n408), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(KEYINPUT58), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n846), .A2(new_n668), .A3(new_n848), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n852), .B1(new_n856), .B2(G141gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n854), .B1(new_n855), .B2(new_n857), .ZN(G1344gat));
  NAND4_X1  g657(.A1(new_n821), .A2(new_n421), .A3(new_n374), .A4(new_n848), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n846), .A2(new_n374), .A3(new_n848), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n860), .A2(new_n861), .A3(G148gat), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n653), .A2(KEYINPUT121), .A3(new_n823), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n354), .B2(new_n781), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n864), .A2(new_n794), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n863), .B1(new_n827), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n794), .A3(new_n866), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n834), .A2(KEYINPUT122), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(new_n870), .A3(new_n707), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n375), .A2(new_n408), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n844), .A3(new_n453), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n842), .A2(KEYINPUT57), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n874), .A2(new_n374), .A3(new_n848), .A4(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n861), .B1(new_n876), .B2(G148gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n859), .B1(new_n862), .B2(new_n877), .ZN(G1345gat));
  AND2_X1   g677(.A1(new_n846), .A2(new_n848), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(G155gat), .A3(new_n262), .ZN(new_n880));
  INV_X1    g679(.A(G155gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n851), .B2(new_n707), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(G1346gat));
  NAND3_X1  g682(.A1(new_n879), .A2(G162gat), .A3(new_n653), .ZN(new_n884));
  INV_X1    g683(.A(G162gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n885), .B1(new_n851), .B2(new_n354), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n884), .A2(new_n886), .ZN(G1347gat));
  NAND2_X1  g686(.A1(new_n798), .A2(new_n800), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n659), .A2(new_n632), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n630), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G169gat), .B1(new_n890), .B2(new_n408), .ZN(new_n891));
  INV_X1    g690(.A(new_n890), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT123), .ZN(new_n893));
  INV_X1    g692(.A(G169gat), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n893), .A2(new_n894), .A3(new_n668), .A4(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n891), .B1(new_n899), .B2(new_n900), .ZN(G1348gat));
  AND2_X1   g700(.A1(new_n893), .A2(new_n896), .ZN(new_n902));
  AOI21_X1  g701(.A(G176gat), .B1(new_n902), .B2(new_n374), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n890), .A2(new_n690), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(G176gat), .B2(new_n904), .ZN(G1349gat));
  NAND3_X1  g704(.A1(new_n892), .A2(new_n262), .A3(new_n527), .ZN(new_n906));
  OAI21_X1  g705(.A(G183gat), .B1(new_n890), .B2(new_n707), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(KEYINPUT125), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n908), .B(new_n910), .ZN(G1350gat));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n913));
  OAI221_X1 g712(.A(G190gat), .B1(new_n912), .B2(new_n913), .C1(new_n890), .C2(new_n354), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n902), .A2(new_n528), .A3(new_n653), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1351gat));
  NAND2_X1  g717(.A1(new_n889), .A2(new_n620), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n874), .A2(new_n875), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G197gat), .B1(new_n921), .B2(new_n408), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n821), .A2(new_n920), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n667), .A2(G197gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(G1352gat));
  NOR3_X1   g724(.A1(new_n923), .A2(G204gat), .A3(new_n690), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT62), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n874), .A2(new_n374), .A3(new_n875), .ZN(new_n928));
  OAI21_X1  g727(.A(G204gat), .B1(new_n928), .B2(new_n919), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1353gat));
  INV_X1    g729(.A(new_n923), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n427), .A3(new_n262), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n874), .A2(new_n262), .A3(new_n875), .A4(new_n920), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n933), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT63), .B1(new_n933), .B2(G211gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(G1354gat));
  NAND4_X1  g735(.A1(new_n874), .A2(new_n653), .A3(new_n875), .A4(new_n920), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G218gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n931), .A2(new_n428), .A3(new_n653), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n938), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1355gat));
endmodule


