//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT64), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(G143), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT68), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G146), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n187), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n191), .A2(G128), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT69), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n205), .B1(new_n202), .B2(G143), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n193), .A2(new_n195), .A3(G128), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT69), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n204), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT71), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n216), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n217));
  INV_X1    g031(.A(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G134), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n219), .A2(KEYINPUT66), .A3(KEYINPUT11), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT11), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n221), .A2(new_n222), .B1(new_n218), .B2(G134), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n217), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G131), .ZN(new_n225));
  INV_X1    g039(.A(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n216), .A2(G137), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(new_n219), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n208), .A2(new_n209), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n211), .A2(KEYINPUT69), .A3(new_n212), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(new_n204), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n215), .A2(new_n229), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G116), .B(G119), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT2), .B(G113), .Z(new_n239));
  XOR2_X1   g053(.A(new_n238), .B(new_n239), .Z(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT67), .A2(G131), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n224), .B(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n191), .A2(KEYINPUT0), .A3(G128), .A4(new_n206), .ZN(new_n245));
  INV_X1    g059(.A(new_n203), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n235), .A2(new_n241), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT28), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT28), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n235), .A2(new_n253), .A3(new_n241), .A4(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G237), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(G210), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n258), .B(KEYINPUT27), .Z(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n248), .A2(KEYINPUT65), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n245), .B(new_n264), .C1(new_n246), .C2(new_n247), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n244), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n214), .A2(new_n229), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n241), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n255), .A2(new_n262), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT73), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n268), .B1(new_n252), .B2(new_n254), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n274), .A3(new_n262), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n271), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n235), .A2(KEYINPUT30), .A3(new_n250), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n266), .A2(new_n267), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n280), .A3(new_n240), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n251), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n261), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n262), .B1(new_n281), .B2(new_n251), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT74), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT75), .B1(new_n276), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n286), .B(new_n284), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n261), .B(new_n268), .C1(new_n252), .C2(new_n254), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT29), .B1(new_n291), .B2(new_n274), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n290), .A2(new_n292), .A3(new_n293), .A4(new_n271), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n235), .A2(new_n250), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n240), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n255), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n261), .A2(new_n272), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n289), .A2(new_n294), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G472), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n281), .A2(new_n262), .A3(new_n251), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT31), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT31), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n281), .A2(new_n304), .A3(new_n262), .A4(new_n251), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n303), .B(new_n305), .C1(new_n262), .C2(new_n273), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT72), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT32), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n301), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G217), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(G234), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT25), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT82), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G128), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n321));
  OAI211_X1 g135(.A(G119), .B(new_n320), .C1(new_n321), .C2(KEYINPUT23), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n323));
  INV_X1    g137(.A(G119), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(G128), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT77), .B1(new_n324), .B2(G128), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G110), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT78), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT24), .B(G110), .Z(new_n330));
  XNOR2_X1  g144(.A(G119), .B(G128), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n332), .B(KEYINPUT76), .Z(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  OR3_X1    g148(.A1(new_n334), .A2(KEYINPUT16), .A3(G140), .ZN(new_n335));
  XOR2_X1   g149(.A(G125), .B(G140), .Z(new_n336));
  INV_X1    g150(.A(KEYINPUT16), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(G146), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n329), .A2(new_n333), .A3(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(G146), .B(new_n335), .C1(new_n336), .C2(new_n337), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n342), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n345), .A2(KEYINPUT80), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(KEYINPUT80), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n202), .A3(new_n347), .ZN(new_n348));
  OAI22_X1  g162(.A1(new_n327), .A2(G110), .B1(new_n331), .B2(new_n330), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n343), .A2(new_n344), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n350), .A2(new_n351), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n340), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT22), .B(G137), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n355), .B(new_n356), .Z(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n340), .B(new_n357), .C1(new_n352), .C2(new_n353), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n319), .B1(new_n361), .B2(G902), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n359), .A2(new_n360), .A3(new_n314), .A4(new_n318), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n316), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n315), .A2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n312), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n256), .A2(new_n257), .A3(G214), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT91), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(G143), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n372), .B1(KEYINPUT90), .B2(G143), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n375), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n226), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT17), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT90), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT91), .B1(new_n382), .B2(new_n199), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(new_n373), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n377), .B1(new_n384), .B2(new_n371), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G131), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n380), .A2(new_n381), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT93), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(new_n386), .B2(new_n381), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n385), .A2(KEYINPUT93), .A3(KEYINPUT17), .A4(G131), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n339), .A4(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n348), .B1(new_n187), .B2(new_n345), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT18), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n379), .B1(new_n393), .B2(new_n226), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n392), .B(new_n394), .C1(new_n393), .C2(new_n386), .ZN(new_n395));
  XNOR2_X1  g209(.A(G113), .B(G122), .ZN(new_n396));
  INV_X1    g210(.A(G104), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n398), .B(KEYINPUT92), .Z(new_n399));
  AND3_X1   g213(.A1(new_n391), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n341), .B(KEYINPUT79), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n380), .A2(new_n386), .ZN(new_n402));
  INV_X1    g216(.A(new_n202), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT19), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n346), .A2(new_n404), .A3(new_n347), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n404), .B2(new_n345), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n401), .B(new_n402), .C1(new_n403), .C2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n398), .B1(new_n407), .B2(new_n395), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(G475), .A2(G902), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT94), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT94), .B1(G475), .B2(G902), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT95), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n410), .B1(new_n400), .B2(new_n408), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT20), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT95), .ZN(new_n419));
  INV_X1    g233(.A(new_n415), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n419), .B(new_n420), .C1(new_n400), .C2(new_n408), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n416), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n398), .B1(new_n391), .B2(new_n395), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n314), .B1(new_n400), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT96), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT96), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n426), .B(new_n314), .C1(new_n400), .C2(new_n423), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(G475), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n199), .A2(G128), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n199), .A2(G128), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT13), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT98), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n432), .B2(new_n430), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n433), .A2(KEYINPUT98), .ZN(new_n436));
  OAI21_X1  g250(.A(G134), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G116), .B(G122), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G107), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT83), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G107), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n441), .A3(new_n443), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT97), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT97), .ZN(new_n450));
  INV_X1    g264(.A(new_n430), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n451), .A2(new_n431), .A3(G134), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT99), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n437), .A2(new_n449), .A3(new_n450), .A4(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G116), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(KEYINPUT14), .A3(G122), .ZN(new_n456));
  OAI211_X1 g270(.A(G107), .B(new_n456), .C1(new_n439), .C2(KEYINPUT14), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n451), .A2(new_n431), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n216), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n457), .B(new_n446), .C1(new_n452), .C2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT9), .B(G234), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n461), .A2(new_n313), .A3(G953), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n454), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n454), .B2(new_n460), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n314), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT100), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n454), .A2(new_n460), .ZN(new_n468));
  INV_X1    g282(.A(new_n462), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n470), .B2(new_n463), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT100), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G478), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT15), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n467), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n471), .B1(KEYINPUT15), .B2(new_n474), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n429), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n257), .A2(G952), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(G234), .B2(G237), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n314), .B(new_n257), .C1(G234), .C2(G237), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT21), .B(G898), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G214), .B1(G237), .B2(G902), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT3), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n440), .B1(new_n486), .B2(G104), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(G104), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n397), .A2(KEYINPUT3), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n441), .A3(new_n443), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G101), .ZN(new_n493));
  INV_X1    g307(.A(G101), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n493), .A2(KEYINPUT84), .A3(KEYINPUT4), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT84), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n494), .B1(new_n489), .B2(new_n491), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n240), .B(new_n496), .C1(new_n497), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n494), .B1(G104), .B2(G107), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n444), .B2(G104), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT85), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n495), .A2(KEYINPUT85), .A3(new_n504), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n239), .A2(new_n236), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n236), .A2(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n324), .A2(G116), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n510), .B(G113), .C1(KEYINPUT5), .C2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n502), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(G110), .B(G122), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n502), .A2(new_n515), .A3(new_n513), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(KEYINPUT6), .A3(new_n518), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n230), .A2(new_n231), .B1(new_n198), .B2(new_n203), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n334), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n248), .A2(G125), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G224), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(G953), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n523), .B(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT6), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n514), .A2(new_n527), .A3(new_n516), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n519), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT7), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n521), .A2(new_n522), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n521), .B2(new_n522), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n515), .B(KEYINPUT8), .Z(new_n534));
  NAND2_X1  g348(.A1(new_n512), .A2(new_n509), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n505), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n513), .B2(new_n536), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(G902), .B1(new_n538), .B2(new_n518), .ZN(new_n539));
  OAI21_X1  g353(.A(G210), .B1(G237), .B2(G902), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n529), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n529), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n485), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(KEYINPUT89), .B(new_n485), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n484), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n495), .A2(KEYINPUT85), .A3(new_n504), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT85), .B1(new_n495), .B2(new_n504), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n215), .A2(KEYINPUT10), .A3(new_n234), .A4(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n244), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n320), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n211), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n232), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n505), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT10), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n249), .B(new_n496), .C1(new_n497), .C2(new_n501), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n551), .A2(new_n552), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  XOR2_X1   g375(.A(G110), .B(G140), .Z(new_n562));
  NAND2_X1  g376(.A1(new_n257), .A2(G227), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT88), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT88), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n551), .A2(new_n559), .A3(new_n560), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n244), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n561), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n505), .B1(new_n232), .B2(new_n554), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n232), .B(new_n204), .C1(new_n548), .C2(new_n549), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(KEYINPUT86), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT86), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n520), .B(new_n579), .C1(new_n549), .C2(new_n548), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n575), .B(new_n552), .C1(new_n578), .C2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT86), .B1(new_n550), .B2(new_n214), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n580), .A3(new_n557), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n244), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n575), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT87), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n581), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(KEYINPUT87), .A3(new_n575), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n574), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(G469), .B(new_n573), .C1(new_n589), .C2(new_n565), .ZN(new_n590));
  INV_X1    g404(.A(G469), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n566), .B1(new_n587), .B2(new_n588), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n565), .B1(new_n572), .B2(new_n561), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n591), .B(new_n314), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n591), .A2(new_n314), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n590), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(G221), .B1(new_n461), .B2(G902), .ZN(new_n598));
  AND4_X1   g412(.A1(new_n479), .A2(new_n547), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n370), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n494), .ZN(G3));
  INV_X1    g415(.A(G472), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n306), .B2(new_n314), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n604), .A2(new_n310), .A3(new_n368), .ZN(new_n605));
  INV_X1    g419(.A(new_n598), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n552), .B1(new_n578), .B2(new_n580), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n586), .B1(new_n607), .B2(KEYINPUT12), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(KEYINPUT12), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n588), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n593), .B1(new_n610), .B2(new_n567), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(G902), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n595), .B1(new_n612), .B2(new_n591), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n606), .B1(new_n613), .B2(new_n590), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n605), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT101), .ZN(new_n616));
  INV_X1    g430(.A(new_n485), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n529), .A2(new_n539), .ZN(new_n618));
  INV_X1    g432(.A(new_n540), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n529), .A2(new_n539), .A3(new_n540), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n467), .A2(new_n473), .A3(new_n474), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n464), .A2(KEYINPUT33), .A3(new_n465), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n470), .B2(new_n463), .ZN(new_n626));
  OAI211_X1 g440(.A(G478), .B(new_n314), .C1(new_n624), .C2(new_n626), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n422), .A2(new_n428), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n484), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n622), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n616), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n428), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n417), .B(KEYINPUT20), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n478), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n622), .A2(new_n629), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n616), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  INV_X1    g458(.A(new_n354), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT36), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n645), .B1(new_n646), .B2(new_n357), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n354), .A2(KEYINPUT36), .A3(new_n358), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n647), .A2(new_n366), .A3(new_n648), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n364), .A2(new_n649), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n604), .A2(new_n310), .A3(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n651), .A2(new_n614), .A3(new_n479), .A4(new_n547), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  NAND2_X1  g468(.A1(new_n650), .A2(new_n622), .ZN(new_n655));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n481), .B1(new_n482), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n636), .A2(new_n478), .A3(new_n637), .A4(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n299), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n292), .A2(new_n285), .A3(new_n287), .A4(new_n271), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(KEYINPUT75), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n602), .B1(new_n663), .B2(new_n294), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT32), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n310), .B(new_n665), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n614), .B(new_n660), .C1(new_n664), .C2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n312), .A2(KEYINPUT103), .A3(new_n614), .A4(new_n660), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XOR2_X1   g486(.A(new_n657), .B(KEYINPUT39), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n614), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT40), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n296), .A2(new_n261), .A3(new_n251), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n314), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n261), .B1(new_n281), .B2(new_n251), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n311), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n620), .A2(new_n621), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT38), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n364), .A2(new_n649), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n422), .A2(new_n428), .ZN(new_n686));
  INV_X1    g500(.A(new_n478), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n684), .A2(new_n485), .A3(new_n685), .A4(new_n688), .ZN(new_n689));
  OR3_X1    g503(.A1(new_n675), .A2(new_n682), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  NAND2_X1  g505(.A1(new_n597), .A2(new_n598), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n301), .B2(new_n311), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n628), .A2(new_n658), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n655), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  OAI21_X1  g511(.A(G469), .B1(new_n611), .B2(G902), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n594), .A2(new_n698), .A3(KEYINPUT105), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n700), .B(G469), .C1(new_n611), .C2(G902), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n606), .B(new_n630), .C1(new_n699), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n370), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND2_X1  g519(.A1(new_n699), .A2(new_n701), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n598), .A3(new_n622), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n311), .B2(new_n301), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n368), .A2(new_n638), .A3(new_n478), .A4(new_n629), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NOR4_X1   g525(.A1(new_n685), .A2(new_n478), .A3(new_n429), .A4(new_n484), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  AOI21_X1  g528(.A(new_n606), .B1(new_n699), .B2(new_n701), .ZN(new_n715));
  INV_X1    g529(.A(new_n305), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n255), .A2(new_n296), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n717), .A2(new_n261), .B1(new_n302), .B2(KEYINPUT31), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n303), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n262), .B1(new_n255), .B2(new_n296), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT106), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n308), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n603), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n640), .A2(new_n686), .A3(new_n687), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n715), .A2(new_n725), .A3(new_n368), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n303), .B1(new_n297), .B2(new_n262), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n305), .B1(new_n730), .B2(KEYINPUT106), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n718), .A2(new_n719), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n309), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n694), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n604), .A3(new_n650), .A4(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n729), .B1(new_n707), .B2(new_n735), .ZN(new_n736));
  AOI211_X1 g550(.A(new_n606), .B(new_n543), .C1(new_n699), .C2(new_n701), .ZN(new_n737));
  NOR4_X1   g551(.A1(new_n724), .A2(new_n603), .A3(new_n694), .A4(new_n685), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(KEYINPUT107), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  NAND3_X1  g555(.A1(new_n620), .A2(new_n485), .A3(new_n621), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT108), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n743), .A2(new_n597), .A3(new_n598), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n312), .A2(new_n744), .A3(new_n368), .A4(new_n734), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n745), .A2(KEYINPUT109), .A3(KEYINPUT42), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT42), .B1(new_n745), .B2(KEYINPUT109), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  INV_X1    g563(.A(new_n659), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n312), .A2(new_n744), .A3(new_n368), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  NAND2_X1  g566(.A1(new_n623), .A2(new_n627), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n686), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n685), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n604), .A2(new_n310), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n754), .B(KEYINPUT43), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT111), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n573), .B1(new_n589), .B2(new_n565), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n591), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n767), .A2(KEYINPUT110), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT110), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n596), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n594), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n598), .B(new_n673), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n743), .B1(new_n762), .B2(new_n763), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT112), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(KEYINPUT112), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n764), .B(new_n776), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n218), .ZN(G39));
  INV_X1    g595(.A(new_n743), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n312), .A2(new_n368), .A3(new_n694), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n598), .B1(new_n774), .B2(new_n775), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g601(.A(KEYINPUT47), .B(new_n598), .C1(new_n774), .C2(new_n775), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g603(.A(KEYINPUT113), .B(G140), .Z(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G42));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n312), .B(new_n368), .C1(new_n599), .C2(new_n702), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n312), .B(new_n737), .C1(new_n709), .C2(new_n712), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n628), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n687), .B2(new_n429), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n605), .A2(new_n614), .A3(new_n547), .A4(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n652), .A2(new_n798), .A3(new_n727), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n685), .A2(new_n478), .A3(new_n657), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n312), .A2(new_n744), .A3(new_n638), .A4(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n751), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n614), .A2(new_n743), .ZN(new_n803));
  OR3_X1    g617(.A1(new_n803), .A2(new_n735), .A3(KEYINPUT115), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT115), .B1(new_n803), .B2(new_n735), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n795), .A2(new_n799), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n747), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n745), .A2(KEYINPUT109), .A3(KEYINPUT42), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n792), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n802), .A2(new_n806), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n799), .A2(new_n793), .A3(new_n794), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n812), .A2(new_n748), .A3(new_n814), .A4(KEYINPUT116), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n736), .A2(new_n739), .B1(new_n693), .B2(new_n695), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n688), .A2(new_n622), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n650), .A3(new_n657), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n680), .A2(new_n614), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n671), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n671), .A2(new_n817), .A3(KEYINPUT52), .A4(new_n820), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT117), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(KEYINPUT117), .A3(new_n824), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n816), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n823), .A2(new_n824), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n816), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n829), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n823), .A2(KEYINPUT117), .A3(new_n824), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n825), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT53), .B1(new_n835), .B2(new_n816), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n807), .A2(new_n810), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n831), .A3(KEYINPUT53), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n836), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n756), .A2(new_n481), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT119), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n368), .A3(new_n725), .ZN(new_n844));
  INV_X1    g658(.A(new_n715), .ZN(new_n845));
  OR3_X1    g659(.A1(new_n845), .A2(new_n485), .A3(new_n684), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT50), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n706), .B(KEYINPUT114), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n606), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n787), .A2(new_n788), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n844), .A2(new_n782), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n845), .A2(new_n782), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n682), .A2(new_n368), .A3(new_n481), .A4(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n855), .A2(new_n429), .A3(new_n753), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n650), .A2(new_n843), .A3(new_n725), .A4(new_n854), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n848), .A2(new_n853), .A3(KEYINPUT51), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n843), .A2(new_n370), .A3(new_n854), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT48), .Z(new_n861));
  NOR2_X1   g675(.A1(new_n855), .A2(new_n796), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n844), .A2(new_n707), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n861), .A2(new_n480), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n787), .A2(new_n788), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT120), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n850), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n866), .A2(KEYINPUT120), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n852), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n848), .A3(new_n858), .ZN(new_n871));
  XNOR2_X1  g685(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n865), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n841), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(G952), .A2(G953), .ZN(new_n875));
  INV_X1    g689(.A(new_n849), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(KEYINPUT49), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n368), .A2(new_n598), .A3(new_n485), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n684), .A2(new_n878), .A3(new_n754), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT49), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n682), .B(new_n879), .C1(new_n880), .C2(new_n849), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n874), .A2(new_n875), .B1(new_n877), .B2(new_n881), .ZN(G75));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n883));
  OAI211_X1 g697(.A(G210), .B(G902), .C1(new_n836), .C2(new_n839), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n519), .A2(new_n528), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(new_n526), .Z(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n884), .A2(new_n885), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n257), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n889), .B1(new_n884), .B2(new_n885), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n883), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n884), .A2(new_n885), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n888), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(KEYINPUT121), .A3(new_n890), .A4(new_n892), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(G51));
  AOI21_X1  g713(.A(new_n839), .B1(new_n828), .B2(new_n830), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n314), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n769), .A2(new_n770), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n595), .B(KEYINPUT57), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n900), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n907), .B1(new_n909), .B2(new_n840), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n592), .B2(new_n593), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n891), .B1(new_n906), .B2(new_n911), .ZN(G54));
  NAND3_X1  g726(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n913), .A2(new_n409), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n409), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n891), .ZN(G60));
  NOR2_X1   g730(.A1(new_n624), .A2(new_n626), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT123), .Z(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT59), .Z(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n909), .B2(new_n840), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(KEYINPUT124), .A3(new_n892), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n924));
  INV_X1    g738(.A(new_n921), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT54), .B1(new_n836), .B2(new_n839), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n828), .A2(new_n830), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n908), .A3(new_n838), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n925), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n924), .B1(new_n929), .B2(new_n891), .ZN(new_n930));
  INV_X1    g744(.A(new_n920), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n833), .B2(new_n840), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n918), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n923), .A2(new_n930), .A3(new_n933), .ZN(G63));
  OAI21_X1  g748(.A(new_n892), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT60), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n900), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n647), .A2(new_n648), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n361), .B1(new_n900), .B2(new_n937), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n940), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(G66));
  OAI21_X1  g759(.A(G953), .B1(new_n483), .B2(new_n524), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n814), .B2(G953), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n886), .B1(G898), .B2(new_n257), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G69));
  NOR2_X1   g763(.A1(new_n780), .A2(new_n789), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n776), .A2(new_n369), .A3(new_n818), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n671), .A2(new_n817), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n748), .A2(new_n952), .A3(new_n751), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n950), .A2(new_n257), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n277), .A2(new_n280), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n406), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n955), .B(new_n957), .C1(new_n656), .C2(new_n257), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n690), .A2(new_n952), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT62), .Z(new_n960));
  INV_X1    g774(.A(new_n674), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n370), .A2(new_n961), .A3(new_n743), .A4(new_n797), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n950), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(new_n257), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n958), .B1(new_n964), .B2(new_n957), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n257), .B1(G227), .B2(G900), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n958), .B2(KEYINPUT126), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n965), .A2(new_n967), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(G72));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n963), .B2(new_n813), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n678), .ZN(new_n974));
  INV_X1    g788(.A(new_n972), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n290), .B2(new_n302), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n829), .A2(new_n832), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n282), .A2(new_n262), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT127), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n950), .A2(new_n814), .A3(new_n954), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n979), .B1(new_n980), .B2(new_n975), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n892), .A2(new_n974), .A3(new_n977), .A4(new_n981), .ZN(G57));
endmodule


