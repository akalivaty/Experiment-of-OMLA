//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT71), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT71), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G211gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT22), .B1(new_n208), .B2(G218gat), .ZN(new_n209));
  XOR2_X1   g008(.A(G197gat), .B(G204gat), .Z(new_n210));
  OAI21_X1  g009(.A(new_n203), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n210), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT71), .B(G211gat), .ZN(new_n213));
  INV_X1    g012(.A(G218gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n202), .B(new_n212), .C1(new_n215), .C2(KEYINPUT22), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT72), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n211), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OAI211_X1 g017(.A(KEYINPUT72), .B(new_n203), .C1(new_n209), .C2(new_n210), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT28), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT27), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G190gat), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n224), .A2(new_n226), .A3(new_n228), .A4(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n232));
  NAND2_X1  g031(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n225), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n221), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT69), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n237), .B(new_n221), .C1(new_n231), .C2(new_n234), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT66), .B(G190gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT27), .B(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT28), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G169gat), .ZN(new_n243));
  INV_X1    g042(.A(G176gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  NOR2_X1   g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(new_n244), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT26), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n248), .A2(new_n250), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n242), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n247), .A2(KEYINPUT23), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(new_n245), .ZN(new_n254));
  OR2_X1    g053(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n255), .A2(KEYINPUT23), .A3(new_n243), .A4(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(KEYINPUT65), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT24), .B1(new_n225), .B2(new_n227), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT24), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(G183gat), .A3(G190gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n225), .A2(new_n227), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT25), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT65), .B1(new_n254), .B2(new_n257), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n239), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n262), .B1(new_n268), .B2(G183gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n247), .A2(KEYINPUT23), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n271), .A2(new_n253), .A3(new_n245), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n265), .A2(new_n267), .B1(KEYINPUT25), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n275));
  INV_X1    g074(.A(G226gat), .ZN(new_n276));
  INV_X1    g075(.A(G233gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n252), .A2(new_n274), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n251), .ZN(new_n281));
  INV_X1    g080(.A(new_n241), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n282), .B1(new_n235), .B2(KEYINPUT69), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n281), .B1(new_n283), .B2(new_n238), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n254), .A2(new_n270), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n239), .A2(new_n225), .B1(new_n259), .B2(new_n261), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT25), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n258), .A2(new_n264), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(new_n266), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n284), .A2(new_n289), .A3(new_n278), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n220), .B1(new_n280), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n252), .A2(new_n274), .A3(new_n279), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n279), .A2(new_n275), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n284), .B2(new_n289), .ZN(new_n295));
  INV_X1    g094(.A(new_n220), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n291), .A2(new_n292), .A3(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(KEYINPUT73), .B(new_n220), .C1(new_n280), .C2(new_n290), .ZN(new_n299));
  XNOR2_X1  g098(.A(G8gat), .B(G36gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(G64gat), .ZN(new_n301));
  INV_X1    g100(.A(G92gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n298), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(new_n298), .B2(new_n299), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n305), .B1(KEYINPUT30), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n297), .A2(new_n292), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n296), .B1(new_n293), .B2(new_n295), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n299), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n303), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT30), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(KEYINPUT74), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(new_n306), .B2(KEYINPUT30), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n307), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT35), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT34), .ZN(new_n319));
  INV_X1    g118(.A(G127gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(G134gat), .ZN(new_n321));
  INV_X1    g120(.A(G134gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(G127gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(G113gat), .B2(G120gat), .ZN(new_n325));
  AND2_X1   g124(.A1(G113gat), .A2(G120gat), .ZN(new_n326));
  OAI22_X1  g125(.A1(new_n321), .A2(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G113gat), .ZN(new_n328));
  INV_X1    g127(.A(G120gat), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT1), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G113gat), .A2(G120gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n322), .A2(G127gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n320), .A2(G134gat), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n327), .A2(new_n334), .A3(KEYINPUT70), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT70), .B1(new_n327), .B2(new_n334), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n252), .A2(new_n274), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n337), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n284), .B2(new_n289), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G227gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(new_n277), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n319), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  AOI211_X1 g144(.A(KEYINPUT34), .B(new_n343), .C1(new_n338), .C2(new_n340), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n338), .A2(new_n340), .A3(new_n343), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT33), .ZN(new_n349));
  XOR2_X1   g148(.A(G15gat), .B(G43gat), .Z(new_n350));
  XNOR2_X1  g149(.A(G71gat), .B(G99gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n348), .B(KEYINPUT32), .C1(new_n349), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n348), .A2(KEYINPUT32), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n348), .A2(new_n349), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n352), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n347), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n220), .B2(KEYINPUT29), .ZN(new_n360));
  NAND3_X1  g159(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT2), .ZN(new_n367));
  INV_X1    g166(.A(G148gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(G141gat), .ZN(new_n369));
  INV_X1    g168(.A(G141gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(G148gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n367), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n368), .B2(G141gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n368), .A2(G141gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n370), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G155gat), .ZN(new_n379));
  INV_X1    g178(.A(G162gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n366), .B1(new_n381), .B2(KEYINPUT2), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n360), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G228gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n365), .A2(new_n372), .B1(new_n378), .B2(new_n382), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n359), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n275), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n220), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n385), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n211), .B2(new_n216), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n384), .B1(new_n394), .B2(KEYINPUT3), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n393), .B1(new_n396), .B2(new_n386), .ZN(new_n397));
  AOI211_X1 g196(.A(KEYINPUT80), .B(new_n387), .C1(new_n391), .C2(new_n395), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n392), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT31), .B(G50gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G22gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(KEYINPUT81), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n404), .B1(new_n406), .B2(new_n402), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n399), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n407), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n392), .B(new_n409), .C1(new_n397), .C2(new_n398), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n345), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n341), .A2(new_n319), .A3(new_n344), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n357), .A2(new_n354), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n358), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT79), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n384), .A2(KEYINPUT3), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n327), .A2(new_n334), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n389), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n420), .B(KEYINPUT77), .Z(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(KEYINPUT5), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(new_n388), .C1(new_n335), .C2(new_n336), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT4), .B1(new_n384), .B2(new_n418), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n424), .A2(KEYINPUT78), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT78), .B1(new_n424), .B2(new_n425), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n419), .B(new_n422), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n388), .A2(new_n327), .A3(new_n334), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n423), .B2(new_n421), .ZN(new_n430));
  OAI211_X1 g229(.A(KEYINPUT4), .B(new_n388), .C1(new_n335), .C2(new_n336), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n419), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n384), .A2(new_n418), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n429), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n421), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(KEYINPUT5), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n428), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT0), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(G57gat), .ZN(new_n440));
  INV_X1    g239(.A(G85gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AND4_X1   g242(.A1(new_n416), .A2(new_n437), .A3(KEYINPUT6), .A4(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n428), .B2(new_n436), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n416), .B1(new_n445), .B2(KEYINPUT6), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT85), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n437), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT79), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n416), .A3(KEYINPUT6), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n445), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n428), .A2(new_n436), .A3(new_n442), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n447), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n317), .A2(new_n318), .A3(new_n415), .A4(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n305), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n306), .A2(KEYINPUT30), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n316), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n456), .A2(new_n451), .A3(new_n449), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n415), .A4(new_n314), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n458), .A2(KEYINPUT87), .B1(KEYINPUT35), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n457), .A2(new_n318), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT87), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n465), .A2(new_n317), .A3(new_n466), .A4(new_n415), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT37), .B1(new_n310), .B2(new_n311), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT37), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n298), .A2(new_n470), .A3(new_n299), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n303), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT38), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n447), .A2(new_n456), .A3(new_n452), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n297), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n297), .A2(new_n476), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(KEYINPUT37), .A3(new_n291), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n471), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n303), .A2(KEYINPUT38), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n306), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n298), .A2(new_n470), .A3(new_n299), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n470), .B1(new_n298), .B2(new_n299), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n304), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(KEYINPUT86), .A3(KEYINPUT38), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n474), .A2(new_n475), .A3(new_n482), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n307), .A2(new_n314), .A3(new_n316), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n419), .B1(new_n426), .B2(new_n427), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT82), .B(KEYINPUT39), .Z(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n421), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n421), .ZN(new_n492));
  INV_X1    g291(.A(new_n427), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT78), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n492), .B1(new_n495), .B2(new_n419), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT39), .B1(new_n434), .B2(new_n421), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n491), .B(new_n442), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n453), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT83), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT83), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n503), .A3(new_n499), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n411), .B1(new_n488), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n307), .A2(new_n462), .A3(new_n314), .A4(new_n316), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n357), .A2(new_n354), .ZN(new_n509));
  INV_X1    g308(.A(new_n347), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n347), .A2(new_n357), .A3(new_n354), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(KEYINPUT36), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n358), .B2(new_n414), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n508), .A2(new_n411), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n464), .A2(new_n467), .B1(new_n507), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G43gat), .B(G50gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n522));
  INV_X1    g321(.A(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(KEYINPUT14), .A3(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n526), .A2(KEYINPUT14), .ZN(new_n528));
  NAND2_X1  g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n521), .B1(new_n530), .B2(KEYINPUT90), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n519), .A2(new_n520), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n530), .B(new_n532), .C1(KEYINPUT90), .C2(new_n521), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT17), .ZN(new_n537));
  INV_X1    g336(.A(G8gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT16), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(G1gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(G1gat), .B2(new_n539), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n543), .B(new_n544), .Z(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n534), .A2(new_n546), .A3(new_n535), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n537), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n536), .A2(new_n545), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  INV_X1    g352(.A(new_n536), .ZN(new_n554));
  INV_X1    g353(.A(new_n545), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(new_n549), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n551), .B(KEYINPUT13), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OAI22_X1  g358(.A1(new_n552), .A2(new_n553), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI221_X1 g361(.A(KEYINPUT92), .B1(new_n557), .B2(new_n559), .C1(new_n552), .C2(new_n553), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n552), .A2(new_n553), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT11), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n243), .ZN(new_n568));
  INV_X1    g367(.A(G197gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT12), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(KEYINPUT88), .Z(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT93), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n564), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n552), .A2(KEYINPUT93), .A3(new_n553), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n571), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n517), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT94), .B(G57gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(G64gat), .ZN(new_n584));
  INV_X1    g383(.A(G64gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(G57gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT9), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n587), .A2(KEYINPUT95), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G57gat), .B(G64gat), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT9), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(new_n588), .A3(new_n590), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT20), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n605), .B(new_n607), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n597), .A2(new_n600), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n555), .B1(new_n609), .B2(KEYINPUT21), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(new_n225), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n608), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G211gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n612), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G134gat), .B(G162gat), .Z(new_n616));
  AND2_X1   g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n616), .B(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(KEYINPUT99), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n619), .A2(KEYINPUT99), .ZN(new_n621));
  NAND2_X1  g420(.A1(G85gat), .A2(G92gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT7), .ZN(new_n623));
  NAND2_X1  g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n624), .B1(new_n441), .B2(new_n302), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G99gat), .B(G106gat), .Z(new_n627));
  OR2_X1    g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n627), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n630), .B(new_n632), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n633), .A2(new_n554), .B1(KEYINPUT41), .B2(new_n617), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n630), .B(new_n631), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n537), .A3(new_n547), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G190gat), .B(G218gat), .Z(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n634), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  AOI211_X1 g440(.A(new_n620), .B(new_n621), .C1(new_n639), .C2(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n639), .A2(new_n620), .A3(new_n641), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G176gat), .ZN(new_n647));
  INV_X1    g446(.A(G204gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(G230gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n277), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n601), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n632), .B1(new_n628), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n626), .A2(new_n654), .A3(new_n627), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n609), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n635), .A2(new_n659), .A3(new_n601), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n652), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n653), .A2(new_n652), .A3(new_n657), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n653), .A2(KEYINPUT101), .A3(new_n657), .A4(new_n652), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n650), .B1(new_n663), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT10), .B1(new_n653), .B2(new_n657), .ZN(new_n670));
  OAI22_X1  g469(.A1(new_n670), .A2(new_n661), .B1(new_n651), .B2(new_n277), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n671), .A2(new_n649), .A3(new_n667), .A4(new_n666), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n615), .A2(new_n645), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n582), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n462), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G1gat), .ZN(G1324gat));
  INV_X1    g478(.A(new_n676), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n317), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  AND2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n683), .A2(KEYINPUT42), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(KEYINPUT42), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n684), .B(new_n685), .C1(new_n538), .C2(new_n681), .ZN(G1325gat));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n515), .A2(new_n687), .A3(new_n513), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n515), .B2(new_n513), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G15gat), .B1(new_n680), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n358), .A2(new_n414), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(G15gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n691), .B1(new_n680), .B2(new_n694), .ZN(G1326gat));
  INV_X1    g494(.A(new_n411), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT103), .B1(new_n680), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n676), .A2(new_n698), .A3(new_n411), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT43), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n697), .A2(new_n702), .A3(new_n699), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n701), .A2(G22gat), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(G22gat), .B1(new_n701), .B2(new_n703), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(G1327gat));
  NOR2_X1   g505(.A1(new_n615), .A2(new_n673), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n644), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n581), .A2(new_n523), .A3(new_n677), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT45), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT44), .B1(new_n517), .B2(new_n645), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n508), .A2(new_n411), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n508), .A2(new_n715), .A3(new_n411), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n507), .A2(new_n690), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n415), .A2(new_n314), .A3(new_n316), .A4(new_n307), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n457), .A2(new_n318), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT87), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n415), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT35), .B1(new_n721), .B2(new_n508), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(new_n467), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n645), .A2(KEYINPUT44), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT105), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n728), .B(new_n725), .C1(new_n717), .C2(new_n723), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n712), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n573), .A2(new_n579), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n707), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n731), .A2(new_n462), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n711), .B1(new_n734), .B2(new_n523), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT106), .Z(G1328gat));
  NAND4_X1  g535(.A1(new_n581), .A2(new_n524), .A3(new_n488), .A4(new_n709), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n731), .A2(new_n317), .A3(new_n733), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(new_n524), .ZN(G1329gat));
  NOR2_X1   g540(.A1(new_n731), .A2(new_n733), .ZN(new_n742));
  INV_X1    g541(.A(new_n690), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G43gat), .ZN(new_n745));
  NOR4_X1   g544(.A1(new_n582), .A2(G43gat), .A3(new_n693), .A4(new_n708), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT108), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1330gat));
  NAND2_X1  g549(.A1(new_n742), .A2(new_n411), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G50gat), .ZN(new_n752));
  OR4_X1    g551(.A1(G50gat), .A2(new_n582), .A3(new_n696), .A4(new_n708), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1331gat));
  INV_X1    g555(.A(new_n615), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n757), .A2(new_n644), .A3(new_n674), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n724), .A2(new_n580), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT109), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n677), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT110), .Z(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n583), .ZN(G1332gat));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n488), .B1(new_n764), .B2(new_n585), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT111), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n585), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1333gat));
  AND2_X1   g568(.A1(new_n760), .A2(new_n692), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n770), .A2(G71gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n760), .A2(G71gat), .A3(new_n743), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n772), .A2(KEYINPUT112), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(KEYINPUT112), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT50), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n771), .B(new_n777), .C1(new_n773), .C2(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1334gat));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n411), .ZN(new_n780));
  XNOR2_X1  g579(.A(KEYINPUT113), .B(G78gat), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1335gat));
  NOR3_X1   g581(.A1(new_n615), .A2(new_n732), .A3(new_n674), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n730), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n441), .B1(new_n784), .B2(new_n677), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n615), .A2(new_n732), .A3(new_n645), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n724), .A2(KEYINPUT51), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT51), .B1(new_n724), .B2(new_n786), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n673), .A2(new_n441), .A3(new_n677), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT114), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n785), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(G1336gat));
  NOR2_X1   g593(.A1(new_n317), .A2(G92gat), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n673), .B(new_n795), .C1(new_n787), .C2(new_n788), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT118), .Z(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n730), .A2(new_n488), .A3(new_n783), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G92gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n796), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n802), .B1(new_n800), .B2(KEYINPUT116), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n799), .A2(new_n804), .A3(G92gat), .ZN(new_n805));
  AOI211_X1 g604(.A(KEYINPUT117), .B(new_n798), .C1(new_n803), .C2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n800), .A2(KEYINPUT116), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n805), .A3(new_n796), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n807), .B1(new_n809), .B2(KEYINPUT52), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n801), .B1(new_n806), .B2(new_n810), .ZN(G1337gat));
  AND2_X1   g610(.A1(new_n789), .A2(new_n673), .ZN(new_n812));
  INV_X1    g611(.A(G99gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n692), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n784), .A2(new_n743), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n813), .ZN(G1338gat));
  INV_X1    g615(.A(G106gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n812), .A2(new_n817), .A3(new_n411), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n784), .A2(new_n411), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n649), .B1(new_n663), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n660), .A2(new_n652), .A3(new_n662), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n671), .A3(KEYINPUT54), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI221_X1 g627(.A(new_n822), .B1(new_n651), .B2(new_n277), .C1(new_n670), .C2(new_n661), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n825), .A2(KEYINPUT55), .A3(new_n650), .A4(new_n829), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n830), .A2(KEYINPUT119), .A3(new_n672), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT119), .B1(new_n830), .B2(new_n672), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n732), .B(new_n828), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n570), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n556), .A2(new_n549), .A3(new_n558), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n551), .B1(new_n548), .B2(new_n550), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT120), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n579), .A2(new_n673), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n644), .B1(new_n833), .B2(new_n839), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n644), .A2(new_n579), .A3(new_n838), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n841), .B(new_n828), .C1(new_n831), .C2(new_n832), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n757), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n675), .A2(new_n732), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n718), .A2(new_n462), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n732), .ZN(new_n851));
  AOI211_X1 g650(.A(new_n462), .B(new_n488), .C1(new_n844), .C2(new_n846), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n852), .A2(new_n415), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n580), .A2(new_n328), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(G1340gat));
  AOI21_X1  g654(.A(G120gat), .B1(new_n850), .B2(new_n673), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n674), .A2(new_n329), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n853), .B2(new_n857), .ZN(G1341gat));
  NOR3_X1   g657(.A1(new_n849), .A2(G127gat), .A3(new_n757), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n853), .A2(new_n615), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(G127gat), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n861), .B(KEYINPUT121), .Z(G1342gat));
  NAND3_X1  g661(.A1(new_n850), .A2(new_n322), .A3(new_n644), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT56), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n322), .B1(new_n853), .B2(new_n644), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n864), .A2(new_n865), .ZN(G1343gat));
  AND3_X1   g665(.A1(new_n852), .A2(new_n411), .A3(new_n690), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n867), .A2(new_n370), .A3(new_n732), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(KEYINPUT58), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n488), .A2(new_n462), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n690), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n696), .B1(new_n844), .B2(new_n846), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n579), .A2(new_n673), .A3(new_n838), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n830), .A2(new_n672), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT55), .B1(new_n823), .B2(new_n825), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n875), .B1(new_n878), .B2(new_n732), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT122), .B1(new_n879), .B2(new_n644), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n828), .A2(new_n672), .A3(new_n830), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n839), .B1(new_n881), .B2(new_n580), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n883), .A3(new_n645), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n884), .A3(new_n842), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n845), .B1(new_n885), .B2(new_n757), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n696), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n874), .A2(new_n887), .A3(new_n732), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n869), .B1(new_n370), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n874), .A2(new_n887), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n874), .B2(new_n887), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n732), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n868), .B1(new_n894), .B2(G141gat), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n889), .B1(new_n895), .B2(new_n896), .ZN(G1344gat));
  NAND2_X1  g696(.A1(new_n368), .A2(KEYINPUT59), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n867), .B2(new_n673), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n891), .A2(new_n892), .A3(new_n674), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n882), .A2(new_n645), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n842), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n845), .B1(new_n902), .B2(new_n757), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(KEYINPUT57), .A3(new_n696), .ZN(new_n904));
  INV_X1    g703(.A(new_n872), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(KEYINPUT57), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n673), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n690), .A2(KEYINPUT59), .A3(new_n870), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n900), .A2(KEYINPUT59), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n899), .B1(new_n909), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g709(.A(new_n379), .B1(new_n893), .B2(new_n615), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n867), .A2(new_n379), .A3(new_n615), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT124), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n891), .A2(new_n892), .A3(new_n757), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n915), .B(new_n912), .C1(new_n916), .C2(new_n379), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(new_n917), .ZN(G1346gat));
  NAND3_X1  g717(.A1(new_n867), .A2(new_n380), .A3(new_n644), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n891), .A2(new_n892), .A3(new_n645), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n380), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n317), .A2(new_n677), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(new_n721), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n847), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(new_n580), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(new_n243), .ZN(G1348gat));
  NOR2_X1   g726(.A1(new_n925), .A2(new_n674), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n255), .A2(new_n256), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(G176gat), .B2(new_n928), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT125), .ZN(G1349gat));
  NAND4_X1  g731(.A1(new_n847), .A2(new_n240), .A3(new_n615), .A4(new_n924), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G183gat), .B1(new_n925), .B2(new_n757), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n934), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g738(.A1(new_n925), .A2(new_n645), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n940), .B2(new_n227), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n942), .B(new_n944), .C1(new_n268), .C2(new_n941), .ZN(G1351gat));
  NOR2_X1   g744(.A1(new_n743), .A2(new_n923), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n872), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n732), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n946), .B(KEYINPUT127), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n949), .A2(new_n569), .A3(new_n580), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n906), .B2(new_n950), .ZN(G1352gat));
  NAND3_X1  g750(.A1(new_n947), .A2(new_n648), .A3(new_n673), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  OAI21_X1  g752(.A(G204gat), .B1(new_n907), .B2(new_n949), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n947), .A2(new_n213), .A3(new_n615), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n906), .A2(new_n615), .A3(new_n946), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1354gat));
  AOI21_X1  g759(.A(G218gat), .B1(new_n947), .B2(new_n644), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n949), .A2(new_n214), .A3(new_n645), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n906), .B2(new_n962), .ZN(G1355gat));
endmodule


