//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT64), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n460), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  AND3_X1   g041(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n460), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(new_n471), .ZN(G160));
  INV_X1    g047(.A(new_n469), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n480));
  OAI221_X1 g055(.A(G2104), .B1(G112), .B2(new_n460), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n474), .A2(new_n477), .A3(new_n481), .ZN(G162));
  INV_X1    g057(.A(G126), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n460), .A2(G114), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n475), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n467), .B2(new_n468), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT68), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(new_n488), .C1(new_n467), .C2(new_n468), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n461), .A2(new_n488), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n486), .B1(new_n493), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT70), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(new_n498), .A3(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(new_n506), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n498), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT7), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n520), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n511), .A2(G51), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n501), .A2(new_n503), .ZN(new_n523));
  INV_X1    g098(.A(new_n499), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n523), .A2(G89), .A3(new_n524), .A4(new_n513), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n523), .A2(G63), .A3(G651), .A4(new_n524), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  INV_X1    g103(.A(G64), .ZN(new_n529));
  AOI211_X1 g104(.A(new_n529), .B(new_n499), .C1(new_n501), .C2(new_n503), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(G651), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n523), .A2(G90), .A3(new_n524), .A4(new_n513), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n511), .A2(G52), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n533), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  AOI211_X1 g114(.A(new_n539), .B(new_n499), .C1(new_n501), .C2(new_n503), .ZN(new_n540));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(G651), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n523), .A2(G81), .A3(new_n524), .A4(new_n513), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n511), .A2(G43), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n523), .A2(G56), .A3(new_n524), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n506), .B1(new_n549), .B2(new_n541), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n544), .A2(new_n545), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT71), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n548), .A2(G860), .A3(new_n552), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(new_n514), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n513), .A2(G53), .A3(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n511), .A2(new_n561), .A3(G53), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n558), .A2(G91), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g138(.A(KEYINPUT72), .B(G65), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n502), .B1(KEYINPUT5), .B2(new_n498), .ZN(new_n565));
  NOR3_X1   g140(.A1(new_n500), .A2(KEYINPUT70), .A3(G543), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n564), .B(new_n524), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(KEYINPUT73), .B1(new_n569), .B2(G651), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n571));
  AOI211_X1 g146(.A(new_n571), .B(new_n506), .C1(new_n567), .C2(new_n568), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n563), .B1(new_n570), .B2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G166), .ZN(G303));
  OAI21_X1  g149(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n511), .A2(G49), .ZN(new_n576));
  INV_X1    g151(.A(G87), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n514), .ZN(G288));
  NAND2_X1  g153(.A1(new_n511), .A2(G48), .ZN(new_n579));
  INV_X1    g154(.A(G86), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  OAI221_X1 g156(.A(new_n579), .B1(new_n514), .B2(new_n580), .C1(new_n581), .C2(new_n506), .ZN(G305));
  AOI22_X1  g157(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n506), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n511), .A2(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n514), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n584), .A2(new_n587), .ZN(G290));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NOR2_X1   g164(.A1(G301), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n511), .A2(G54), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n504), .A2(G66), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n592), .B1(new_n595), .B2(G651), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n504), .A2(G92), .A3(new_n513), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n504), .A2(KEYINPUT10), .A3(G92), .A4(new_n513), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT74), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n590), .B1(new_n604), .B2(new_n589), .ZN(G284));
  AOI21_X1  g180(.A(new_n590), .B1(new_n604), .B2(new_n589), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n548), .A2(new_n552), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n589), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n603), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n589), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g192(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT13), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n473), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n476), .A2(G123), .ZN(new_n623));
  OR2_X1    g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n624), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n621), .A2(new_n627), .ZN(G156));
  XOR2_X1   g203(.A(G1341), .B(G1348), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT75), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n633), .B(new_n639), .Z(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G14), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n640), .B2(new_n641), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  INV_X1    g221(.A(KEYINPUT18), .ZN(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT17), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2096), .B(G2100), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n650), .B2(KEYINPUT18), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT76), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1981), .B(G1986), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n665), .A2(new_n666), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  MUX2_X1   g247(.A(new_n672), .B(new_n671), .S(new_n664), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT77), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n677), .A2(new_n679), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n661), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n677), .A2(new_n679), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n679), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(new_n660), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(G229));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n690), .A2(G35), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G162), .B2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT29), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(G2090), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n696));
  NAND2_X1  g271(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT3), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n701), .A2(G129), .A3(G2105), .ZN(new_n702));
  NAND3_X1  g277(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT26), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g280(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n705), .A2(new_n706), .B1(new_n465), .B2(G105), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n473), .A2(G141), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G32), .B(new_n710), .S(G29), .Z(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT24), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(G34), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(G34), .ZN(new_n717));
  NOR3_X1   g292(.A1(new_n690), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G160), .B2(G29), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G5), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G171), .B2(new_n720), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n714), .B1(G2084), .B2(new_n719), .C1(new_n722), .C2(G1961), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n695), .A2(new_n696), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  MUX2_X1   g302(.A(G19), .B(new_n613), .S(G16), .Z(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(G1341), .Z(new_n729));
  OR2_X1    g304(.A1(new_n711), .A2(new_n713), .ZN(new_n730));
  INV_X1    g305(.A(new_n690), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n626), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT87), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n731), .A2(G27), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n491), .B1(new_n701), .B2(new_n488), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n496), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n486), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n734), .B1(new_n739), .B2(new_n690), .ZN(new_n740));
  INV_X1    g315(.A(G2078), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n719), .A2(G2084), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n730), .A2(new_n733), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G33), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT85), .B(KEYINPUT25), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n749), .A2(new_n750), .B1(new_n473), .B2(G139), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(new_n460), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n746), .B1(new_n754), .B2(G29), .ZN(new_n755));
  INV_X1    g330(.A(G2072), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT86), .Z(new_n758));
  AOI211_X1 g333(.A(new_n744), .B(new_n758), .C1(new_n741), .C2(new_n740), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n727), .A2(new_n729), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT82), .ZN(new_n761));
  OR3_X1    g336(.A1(new_n761), .A2(G4), .A3(G16), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(G4), .B2(G16), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n762), .B(new_n763), .C1(new_n603), .C2(new_n720), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT83), .B(G1348), .Z(new_n765));
  XOR2_X1   g340(.A(new_n764), .B(new_n765), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n720), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G1956), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n731), .A2(G26), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT28), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n473), .A2(G140), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n460), .A2(G116), .ZN(new_n776));
  OAI21_X1  g351(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT84), .ZN(new_n778));
  OR3_X1    g353(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n776), .B2(new_n777), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n476), .A2(G128), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n775), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(G29), .ZN(new_n784));
  INV_X1    g359(.A(G2067), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G1961), .B2(new_n722), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n693), .B2(G2090), .ZN(new_n789));
  NAND2_X1  g364(.A1(G168), .A2(G16), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G16), .B2(G21), .ZN(new_n791));
  INV_X1    g366(.A(G1966), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G28), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT30), .ZN(new_n795));
  AOI21_X1  g370(.A(G29), .B1(new_n794), .B2(KEYINPUT30), .ZN(new_n796));
  OR2_X1    g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  NAND2_X1  g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n795), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  OAI22_X1  g375(.A1(new_n791), .A2(new_n792), .B1(new_n756), .B2(new_n755), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n787), .A2(new_n789), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n693), .A2(G2090), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(KEYINPUT89), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n760), .A2(new_n772), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n760), .A2(KEYINPUT91), .A3(new_n772), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G6), .A2(G16), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G305), .B2(new_n720), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT32), .B(G1981), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n812), .B(new_n814), .C1(G305), .C2(new_n720), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT80), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(KEYINPUT80), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n720), .A2(G22), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G166), .B2(new_n720), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(G1971), .Z(new_n823));
  MUX2_X1   g398(.A(G23), .B(G288), .S(G16), .Z(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT33), .B(G1976), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n819), .A2(new_n820), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n690), .A2(G25), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n473), .A2(G131), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n476), .A2(G119), .ZN(new_n831));
  OR2_X1    g406(.A1(G95), .A2(G2105), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n832), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n829), .B1(new_n835), .B2(new_n690), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT79), .Z(new_n837));
  XOR2_X1   g412(.A(KEYINPUT35), .B(G1991), .Z(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n720), .A2(G24), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n584), .A2(new_n587), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n720), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G1986), .ZN(new_n844));
  NOR4_X1   g419(.A1(new_n828), .A2(new_n839), .A3(new_n840), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(KEYINPUT81), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(KEYINPUT81), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(KEYINPUT36), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n845), .B(new_n851), .C1(new_n847), .C2(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n810), .A2(new_n853), .ZN(G311));
  AND3_X1   g429(.A1(new_n810), .A2(KEYINPUT92), .A3(new_n853), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT92), .B1(new_n810), .B2(new_n853), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(G150));
  NAND3_X1  g432(.A1(new_n523), .A2(G67), .A3(new_n524), .ZN(new_n858));
  NAND2_X1  g433(.A1(G80), .A2(G543), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n506), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n523), .A2(G93), .A3(new_n524), .A4(new_n513), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n511), .A2(G55), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n548), .B2(new_n552), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n543), .A2(new_n546), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n862), .B(new_n861), .C1(new_n867), .C2(new_n506), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n604), .A2(G559), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n874));
  INV_X1    g449(.A(G860), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n864), .A2(new_n875), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(G145));
  OAI211_X1 g455(.A(G130), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n881));
  OR2_X1    g456(.A1(G106), .A2(G2105), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n882), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n883));
  INV_X1    g458(.A(G142), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n881), .B(new_n883), .C1(new_n469), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n619), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n751), .A2(new_n753), .A3(new_n708), .A4(new_n709), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n751), .A2(new_n753), .B1(new_n708), .B2(new_n709), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n754), .A2(new_n710), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n886), .A3(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n783), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(G164), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n739), .A2(new_n783), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n834), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n834), .B1(new_n896), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n894), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n626), .A2(G160), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n626), .A2(G160), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(G162), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n896), .A2(new_n897), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n835), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n907), .A2(new_n898), .A3(new_n893), .A4(new_n891), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT93), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n901), .A2(KEYINPUT93), .A3(new_n908), .A4(new_n905), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n905), .B1(new_n901), .B2(new_n908), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n914), .A2(G37), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT94), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT94), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n913), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(KEYINPUT95), .B(KEYINPUT40), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(G395));
  NAND2_X1  g497(.A1(new_n868), .A2(new_n589), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n615), .A2(new_n865), .A3(new_n869), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n603), .A2(new_n870), .A3(G559), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(G299), .A2(new_n602), .ZN(new_n927));
  INV_X1    g502(.A(new_n568), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n504), .B2(new_n564), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n571), .B1(new_n929), .B2(new_n506), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n569), .A2(KEYINPUT73), .A3(G651), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n932), .A2(new_n563), .B1(new_n596), .B2(new_n601), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n926), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT41), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n927), .B2(new_n933), .ZN(new_n937));
  NAND2_X1  g512(.A1(G299), .A2(new_n602), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n932), .A2(new_n563), .A3(new_n601), .A4(new_n596), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT41), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n937), .B(new_n940), .C1(new_n924), .C2(new_n925), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT96), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n935), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n942), .B2(new_n941), .ZN(new_n944));
  OR2_X1    g519(.A1(G166), .A2(G288), .ZN(new_n945));
  NAND2_X1  g520(.A1(G166), .A2(G288), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n581), .A2(new_n506), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n579), .B1(new_n514), .B2(new_n580), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(G290), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n842), .A2(G305), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n945), .A2(new_n951), .A3(new_n946), .A4(new_n952), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT42), .Z(new_n957));
  XNOR2_X1  g532(.A(new_n944), .B(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n923), .B1(new_n958), .B2(new_n589), .ZN(G295));
  OAI21_X1  g534(.A(new_n923), .B1(new_n958), .B2(new_n589), .ZN(G331));
  AOI21_X1  g535(.A(new_n547), .B1(new_n543), .B2(new_n546), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT71), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n868), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n869), .ZN(new_n964));
  NAND2_X1  g539(.A1(G63), .A2(G651), .ZN(new_n965));
  AOI211_X1 g540(.A(new_n965), .B(new_n499), .C1(new_n501), .C2(new_n503), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n519), .A2(new_n521), .ZN(new_n967));
  AND2_X1   g542(.A1(KEYINPUT6), .A2(G651), .ZN(new_n968));
  NOR2_X1   g543(.A1(KEYINPUT6), .A2(G651), .ZN(new_n969));
  OAI211_X1 g544(.A(G51), .B(G543), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n523), .A2(G64), .A3(new_n524), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n506), .B1(new_n973), .B2(new_n531), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n534), .A2(new_n535), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n972), .B(new_n525), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n533), .A2(new_n536), .A3(G286), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n963), .A2(new_n964), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n977), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n865), .B2(new_n869), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n937), .A2(new_n940), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n978), .B1(new_n963), .B2(new_n964), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n865), .A2(new_n980), .A3(new_n869), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n934), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n985), .A3(new_n956), .ZN(new_n986));
  INV_X1    g561(.A(G37), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n982), .A2(new_n985), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n956), .B1(new_n989), .B2(KEYINPUT98), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT98), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n982), .A2(new_n985), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n988), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT101), .ZN(new_n996));
  INV_X1    g571(.A(new_n988), .ZN(new_n997));
  AOI211_X1 g572(.A(KEYINPUT100), .B(new_n956), .C1(new_n985), .C2(new_n982), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT100), .ZN(new_n999));
  INV_X1    g574(.A(new_n956), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n989), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n997), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n996), .A2(KEYINPUT44), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT99), .B1(new_n993), .B2(new_n994), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT99), .ZN(new_n1006));
  INV_X1    g581(.A(new_n992), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n991), .B1(new_n982), .B2(new_n985), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n956), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1006), .B(KEYINPUT43), .C1(new_n1009), .C2(new_n988), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n997), .B(new_n994), .C1(new_n998), .C2(new_n1001), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1005), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(KEYINPUT97), .B(KEYINPUT44), .Z(new_n1014));
  OAI21_X1  g589(.A(new_n1004), .B1(new_n1013), .B2(new_n1014), .ZN(G397));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1016), .B1(G168), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  AND4_X1   g596(.A1(new_n461), .A2(new_n488), .A3(new_n494), .A4(new_n495), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT4), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n460), .A2(G138), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n699), .B2(new_n700), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n1025), .B2(new_n491), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1022), .B1(new_n1026), .B2(new_n490), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1020), .B(new_n1021), .C1(new_n1027), .C2(new_n486), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n737), .B2(new_n738), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(KEYINPUT107), .A3(new_n1020), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G160), .A2(G40), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n739), .A2(new_n1021), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(KEYINPUT50), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1019), .B1(new_n1037), .B2(G2084), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1031), .A2(KEYINPUT112), .A3(KEYINPUT45), .ZN(new_n1039));
  AND2_X1   g614(.A1(G160), .A2(G40), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(G164), .B2(G1384), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  AOI211_X1 g618(.A(new_n1041), .B(G1384), .C1(new_n737), .C2(new_n738), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(KEYINPUT112), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n792), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G2084), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1033), .A2(KEYINPUT113), .A3(new_n1047), .A4(new_n1036), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1038), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1018), .B1(new_n1049), .B2(G8), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1040), .B1(new_n1031), .B2(new_n1020), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT113), .B1(new_n1054), .B2(new_n1047), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1051), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1038), .A2(KEYINPUT120), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G168), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1050), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G168), .A2(new_n1017), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1056), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1056), .A2(new_n1057), .A3(KEYINPUT121), .A4(new_n1062), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT62), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(G286), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1060), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1049), .A2(G8), .ZN(new_n1071));
  OAI22_X1  g646(.A1(new_n1069), .A2(new_n1070), .B1(new_n1071), .B2(new_n1018), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G303), .A2(G8), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1037), .A2(G2090), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT106), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT45), .B1(new_n739), .B2(new_n1021), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1044), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1034), .B1(new_n1042), .B2(KEYINPUT106), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(G1971), .ZN(new_n1085));
  OAI211_X1 g660(.A(G8), .B(new_n1077), .C1(new_n1079), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1040), .A2(new_n1031), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G8), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1976), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT52), .B1(G288), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1089), .B(new_n1091), .C1(new_n1090), .C2(G288), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G288), .A2(new_n1090), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT52), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(G1981), .B1(new_n948), .B2(KEYINPUT109), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1096), .A2(G305), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(G305), .ZN(new_n1098));
  OR3_X1    g673(.A1(new_n1097), .A2(new_n1098), .A3(KEYINPUT110), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1099), .A2(KEYINPUT49), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1088), .B1(new_n1099), .B2(KEYINPUT49), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1095), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1085), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(new_n1040), .A3(new_n1028), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1105), .A2(G2090), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1017), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1086), .B(new_n1102), .C1(new_n1107), .C2(new_n1077), .ZN(new_n1108));
  INV_X1    g683(.A(G1961), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1037), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1045), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1081), .A2(new_n1034), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n741), .A2(KEYINPUT53), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1111), .A2(new_n1039), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT122), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1110), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1082), .A2(new_n1083), .A3(new_n741), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1116), .A2(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1108), .A2(G301), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1068), .A2(new_n1074), .A3(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(G288), .A2(G1976), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT111), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G305), .A2(G1981), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1089), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1102), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1086), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1071), .A2(G168), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  OAI21_X1  g708(.A(G8), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1077), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1132), .A2(new_n1086), .A3(new_n1102), .A4(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1133), .B1(new_n1108), .B2(new_n1131), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1130), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n613), .B1(new_n1140), .B2(KEYINPUT59), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n1142));
  INV_X1    g717(.A(G1996), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1082), .A2(new_n1083), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT117), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1082), .A2(new_n1083), .A3(KEYINPUT117), .A4(new_n1143), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT58), .B(G1341), .Z(new_n1149));
  AND2_X1   g724(.A1(new_n1087), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1142), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g727(.A(KEYINPUT118), .B(new_n1150), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1141), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI221_X1 g731(.A(new_n1141), .B1(new_n1140), .B2(KEYINPUT59), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1087), .A2(G2067), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(KEYINPUT60), .B(new_n1159), .C1(new_n1054), .C2(G1348), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n603), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1054), .A2(G1348), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1163), .B2(new_n1158), .ZN(new_n1164));
  INV_X1    g739(.A(G1348), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1037), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1166), .A2(KEYINPUT60), .A3(new_n604), .A4(new_n1159), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1161), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT115), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT57), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n608), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1173));
  NOR3_X1   g748(.A1(G299), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1105), .A2(KEYINPUT114), .A3(new_n770), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT114), .B1(new_n1105), .B2(new_n770), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g753(.A(KEYINPUT56), .B(G2072), .Z(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT116), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1082), .A2(new_n1083), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1175), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1105), .A2(new_n770), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT114), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1105), .A2(KEYINPUT114), .A3(new_n770), .ZN(new_n1186));
  AND4_X1   g761(.A1(new_n1175), .A2(new_n1185), .A3(new_n1181), .A4(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT61), .B1(new_n1182), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1185), .A2(new_n1181), .A3(new_n1186), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1189), .B1(new_n1174), .B2(new_n1171), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1178), .A2(new_n1175), .A3(new_n1181), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1168), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1156), .A2(new_n1157), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n603), .B1(new_n1166), .B2(new_n1159), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1192), .B1(new_n1182), .B2(new_n1196), .ZN(new_n1197));
  AND2_X1   g772(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1118), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1117), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1201));
  OAI211_X1 g776(.A(G301), .B(new_n1199), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT54), .ZN(new_n1203));
  OR2_X1    g778(.A1(new_n1081), .A2(new_n1044), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1040), .A2(KEYINPUT124), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1040), .A2(KEYINPUT124), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1205), .A2(new_n1113), .A3(new_n1206), .ZN(new_n1207));
  OAI211_X1 g782(.A(new_n1199), .B(new_n1110), .C1(new_n1204), .C2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1203), .B1(new_n1208), .B2(G171), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1202), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1202), .A2(new_n1209), .A3(KEYINPUT125), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1208), .A2(G171), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1215), .B1(new_n1121), .B2(G301), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1108), .B1(new_n1216), .B2(new_n1203), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1072), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1214), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  OAI211_X1 g794(.A(new_n1123), .B(new_n1139), .C1(new_n1198), .C2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n1042), .A2(new_n1034), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n783), .B(new_n785), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT104), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n710), .A2(G1996), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1221), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1221), .A2(G1996), .A3(new_n710), .ZN(new_n1226));
  OR2_X1    g801(.A1(new_n1226), .A2(KEYINPUT103), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1226), .A2(KEYINPUT103), .ZN(new_n1228));
  AND3_X1   g803(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  XOR2_X1   g804(.A(new_n834), .B(new_n838), .Z(new_n1230));
  XNOR2_X1  g805(.A(new_n1230), .B(KEYINPUT105), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1231), .A2(new_n1221), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g808(.A(G1986), .ZN(new_n1234));
  AOI21_X1  g809(.A(KEYINPUT102), .B1(new_n842), .B2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g810(.A1(new_n842), .A2(new_n1234), .ZN(new_n1236));
  XNOR2_X1  g811(.A(new_n1235), .B(new_n1236), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1233), .B1(new_n1221), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1220), .A2(new_n1238), .ZN(new_n1239));
  OR2_X1    g814(.A1(new_n1223), .A2(new_n710), .ZN(new_n1240));
  INV_X1    g815(.A(new_n1221), .ZN(new_n1241));
  OAI21_X1  g816(.A(KEYINPUT46), .B1(new_n1241), .B2(G1996), .ZN(new_n1242));
  OR3_X1    g817(.A1(new_n1241), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1243));
  AOI22_X1  g818(.A1(new_n1240), .A2(new_n1221), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g819(.A(new_n1244), .B(KEYINPUT47), .ZN(new_n1245));
  NAND3_X1  g820(.A1(new_n1229), .A2(new_n838), .A3(new_n835), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n895), .A2(new_n785), .ZN(new_n1247));
  AOI21_X1  g822(.A(new_n1241), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g823(.A(new_n1233), .ZN(new_n1249));
  NAND3_X1  g824(.A1(new_n1221), .A2(new_n1234), .A3(new_n842), .ZN(new_n1250));
  XNOR2_X1  g825(.A(new_n1250), .B(KEYINPUT48), .ZN(new_n1251));
  AOI211_X1 g826(.A(new_n1245), .B(new_n1248), .C1(new_n1249), .C2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g827(.A1(new_n1239), .A2(new_n1252), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g828(.A1(G227), .A2(new_n458), .ZN(new_n1255));
  NAND4_X1  g829(.A1(new_n682), .A2(new_n685), .A3(new_n645), .A4(new_n1255), .ZN(new_n1256));
  AOI21_X1  g830(.A(new_n1256), .B1(new_n917), .B2(new_n919), .ZN(new_n1257));
  AND3_X1   g831(.A1(new_n1012), .A2(KEYINPUT126), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g832(.A(KEYINPUT126), .B1(new_n1012), .B2(new_n1257), .ZN(new_n1259));
  NOR3_X1   g833(.A1(new_n1258), .A2(new_n1259), .A3(KEYINPUT127), .ZN(new_n1260));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1261));
  NAND2_X1  g835(.A1(new_n989), .A2(KEYINPUT98), .ZN(new_n1262));
  NAND3_X1  g836(.A1(new_n1262), .A2(new_n1000), .A3(new_n992), .ZN(new_n1263));
  AOI21_X1  g837(.A(new_n994), .B1(new_n1263), .B2(new_n997), .ZN(new_n1264));
  OAI21_X1  g838(.A(new_n1011), .B1(new_n1264), .B2(new_n1006), .ZN(new_n1265));
  NOR3_X1   g839(.A1(new_n993), .A2(KEYINPUT99), .A3(new_n994), .ZN(new_n1266));
  OAI21_X1  g840(.A(new_n1257), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g841(.A(KEYINPUT126), .ZN(new_n1268));
  NAND2_X1  g842(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g843(.A1(new_n1012), .A2(KEYINPUT126), .A3(new_n1257), .ZN(new_n1270));
  AOI21_X1  g844(.A(new_n1261), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g845(.A1(new_n1260), .A2(new_n1271), .ZN(G308));
  NAND2_X1  g846(.A1(new_n1269), .A2(new_n1270), .ZN(G225));
endmodule


