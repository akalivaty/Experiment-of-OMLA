

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X2 U322 ( .A(KEYINPUT64), .B(n419), .ZN(n568) );
  NOR2_X1 U323 ( .A1(n561), .A2(n566), .ZN(n563) );
  XOR2_X1 U324 ( .A(n300), .B(n299), .Z(n290) );
  AND2_X1 U325 ( .A1(n523), .A2(n418), .ZN(n419) );
  XNOR2_X1 U326 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U327 ( .A(n385), .B(n384), .ZN(n576) );
  INV_X1 U328 ( .A(G190GAT), .ZN(n457) );
  XNOR2_X1 U329 ( .A(n457), .B(KEYINPUT58), .ZN(n458) );
  XNOR2_X1 U330 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT75), .B(G92GAT), .Z(n292) );
  XNOR2_X1 U332 ( .A(G99GAT), .B(G85GAT), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n378) );
  XOR2_X1 U334 ( .A(G36GAT), .B(G190GAT), .Z(n405) );
  XOR2_X1 U335 ( .A(n405), .B(G218GAT), .Z(n296) );
  XOR2_X1 U336 ( .A(G29GAT), .B(G43GAT), .Z(n294) );
  XNOR2_X1 U337 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n354) );
  XNOR2_X1 U339 ( .A(n354), .B(G134GAT), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U341 ( .A(KEYINPUT9), .B(KEYINPUT79), .Z(n298) );
  NAND2_X1 U342 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U344 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n302) );
  XNOR2_X1 U345 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n303), .B(G106GAT), .ZN(n304) );
  XNOR2_X1 U348 ( .A(n290), .B(n304), .ZN(n305) );
  XNOR2_X1 U349 ( .A(n378), .B(n305), .ZN(n307) );
  XOR2_X1 U350 ( .A(G50GAT), .B(G162GAT), .Z(n306) );
  XNOR2_X1 U351 ( .A(KEYINPUT78), .B(n306), .ZN(n429) );
  XOR2_X1 U352 ( .A(n307), .B(n429), .Z(n552) );
  INV_X1 U353 ( .A(n552), .ZN(n456) );
  XOR2_X1 U354 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n309) );
  XNOR2_X1 U355 ( .A(G148GAT), .B(KEYINPUT93), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U357 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n311) );
  XNOR2_X1 U358 ( .A(G29GAT), .B(G120GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n325) );
  XOR2_X1 U361 ( .A(G155GAT), .B(KEYINPUT5), .Z(n315) );
  XNOR2_X1 U362 ( .A(KEYINPUT91), .B(KEYINPUT4), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U364 ( .A(KEYINPUT97), .B(KEYINPUT95), .Z(n317) );
  XNOR2_X1 U365 ( .A(G127GAT), .B(KEYINPUT96), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n323) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(G57GAT), .ZN(n321) );
  XOR2_X1 U369 ( .A(G113GAT), .B(G134GAT), .Z(n320) );
  XNOR2_X1 U370 ( .A(KEYINPUT0), .B(n320), .ZN(n449) );
  XNOR2_X1 U371 ( .A(n321), .B(n449), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U374 ( .A(G162GAT), .B(n326), .ZN(n332) );
  XOR2_X1 U375 ( .A(KEYINPUT88), .B(KEYINPUT3), .Z(n328) );
  XNOR2_X1 U376 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n421) );
  XOR2_X1 U378 ( .A(n421), .B(G85GAT), .Z(n330) );
  NAND2_X1 U379 ( .A1(G225GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n523) );
  XOR2_X1 U382 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n350) );
  XNOR2_X1 U383 ( .A(KEYINPUT36), .B(KEYINPUT104), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n552), .B(n333), .ZN(n484) );
  XOR2_X1 U385 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n335) );
  NAND2_X1 U386 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U388 ( .A(KEYINPUT14), .B(n336), .ZN(n348) );
  XOR2_X1 U389 ( .A(KEYINPUT82), .B(G78GAT), .Z(n338) );
  XNOR2_X1 U390 ( .A(G183GAT), .B(G71GAT), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U392 ( .A(G57GAT), .B(KEYINPUT13), .Z(n370) );
  XOR2_X1 U393 ( .A(n339), .B(n370), .Z(n343) );
  XOR2_X1 U394 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n341) );
  XNOR2_X1 U395 ( .A(G1GAT), .B(G8GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n353) );
  XOR2_X1 U397 ( .A(G15GAT), .B(G127GAT), .Z(n440) );
  XNOR2_X1 U398 ( .A(n353), .B(n440), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U400 ( .A(G22GAT), .B(G155GAT), .Z(n425) );
  XOR2_X1 U401 ( .A(n344), .B(n425), .Z(n346) );
  XNOR2_X1 U402 ( .A(G211GAT), .B(G64GAT), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n549) );
  NAND2_X1 U405 ( .A1(n484), .A2(n549), .ZN(n349) );
  XOR2_X1 U406 ( .A(n350), .B(n349), .Z(n388) );
  XOR2_X1 U407 ( .A(G22GAT), .B(G15GAT), .Z(n352) );
  XNOR2_X1 U408 ( .A(KEYINPUT69), .B(KEYINPUT72), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n369) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n367) );
  XOR2_X1 U411 ( .A(G141GAT), .B(G113GAT), .Z(n356) );
  XNOR2_X1 U412 ( .A(G50GAT), .B(G36GAT), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U414 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n358) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(G197GAT), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U417 ( .A(n360), .B(n359), .Z(n365) );
  XOR2_X1 U418 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n362) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U421 ( .A(KEYINPUT29), .B(n363), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n571) );
  INV_X1 U425 ( .A(n571), .ZN(n542) );
  XOR2_X1 U426 ( .A(G176GAT), .B(G64GAT), .Z(n402) );
  XOR2_X1 U427 ( .A(n370), .B(n402), .Z(n372) );
  NAND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U430 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n374) );
  XNOR2_X1 U431 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U433 ( .A(n376), .B(n375), .Z(n385) );
  XNOR2_X1 U434 ( .A(G148GAT), .B(G106GAT), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n377), .B(G78GAT), .ZN(n420) );
  XNOR2_X1 U436 ( .A(n378), .B(n420), .ZN(n383) );
  XOR2_X1 U437 ( .A(G120GAT), .B(G71GAT), .Z(n441) );
  XOR2_X1 U438 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n380) );
  XNOR2_X1 U439 ( .A(G204GAT), .B(KEYINPUT32), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n441), .B(n381), .ZN(n382) );
  INV_X1 U442 ( .A(n576), .ZN(n386) );
  NOR2_X1 U443 ( .A1(n542), .A2(n386), .ZN(n387) );
  NAND2_X1 U444 ( .A1(n388), .A2(n387), .ZN(n396) );
  XNOR2_X1 U445 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n390) );
  XNOR2_X1 U446 ( .A(KEYINPUT41), .B(n576), .ZN(n560) );
  NAND2_X1 U447 ( .A1(n542), .A2(n560), .ZN(n389) );
  XOR2_X1 U448 ( .A(n390), .B(n389), .Z(n391) );
  NOR2_X1 U449 ( .A1(n549), .A2(n391), .ZN(n392) );
  NAND2_X1 U450 ( .A1(n456), .A2(n392), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n393), .B(KEYINPUT47), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n394), .B(KEYINPUT113), .ZN(n395) );
  NAND2_X1 U453 ( .A1(n396), .A2(n395), .ZN(n397) );
  XNOR2_X1 U454 ( .A(KEYINPUT48), .B(n397), .ZN(n525) );
  XNOR2_X1 U455 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n398), .B(KEYINPUT85), .ZN(n399) );
  XOR2_X1 U457 ( .A(n399), .B(KEYINPUT19), .Z(n401) );
  XNOR2_X1 U458 ( .A(G169GAT), .B(G183GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n454) );
  XOR2_X1 U460 ( .A(KEYINPUT99), .B(n402), .Z(n404) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n406) );
  XOR2_X1 U463 ( .A(n406), .B(n405), .Z(n414) );
  XOR2_X1 U464 ( .A(G211GAT), .B(G218GAT), .Z(n408) );
  XNOR2_X1 U465 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U467 ( .A(G197GAT), .B(n409), .Z(n436) );
  XOR2_X1 U468 ( .A(KEYINPUT100), .B(KEYINPUT98), .Z(n411) );
  XNOR2_X1 U469 ( .A(G8GAT), .B(G92GAT), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n436), .B(n412), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n454), .B(n415), .ZN(n478) );
  NAND2_X1 U474 ( .A1(n525), .A2(n478), .ZN(n417) );
  XOR2_X1 U475 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n434) );
  XOR2_X1 U478 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n423) );
  XNOR2_X1 U479 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U481 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U484 ( .A(n428), .B(KEYINPUT87), .Z(n432) );
  INV_X1 U485 ( .A(n429), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n430), .B(KEYINPUT23), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n470) );
  NAND2_X1 U490 ( .A1(n568), .A2(n470), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n437), .B(KEYINPUT55), .ZN(n455) );
  XOR2_X1 U492 ( .A(KEYINPUT86), .B(KEYINPUT83), .Z(n439) );
  XNOR2_X1 U493 ( .A(G190GAT), .B(G176GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n445) );
  XOR2_X1 U495 ( .A(G99GAT), .B(n440), .Z(n443) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U498 ( .A(n445), .B(n444), .Z(n447) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U501 ( .A(n448), .B(KEYINPUT20), .Z(n452) );
  INV_X1 U502 ( .A(n449), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n450), .B(KEYINPUT84), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n454), .B(n453), .ZN(n527) );
  NAND2_X1 U506 ( .A1(n455), .A2(n527), .ZN(n566) );
  NOR2_X1 U507 ( .A1(n456), .A2(n566), .ZN(n459) );
  NAND2_X1 U508 ( .A1(n542), .A2(n576), .ZN(n488) );
  INV_X1 U509 ( .A(n549), .ZN(n580) );
  NOR2_X1 U510 ( .A1(n552), .A2(n580), .ZN(n460) );
  XNOR2_X1 U511 ( .A(KEYINPUT16), .B(n460), .ZN(n475) );
  NAND2_X1 U512 ( .A1(n527), .A2(n478), .ZN(n461) );
  NAND2_X1 U513 ( .A1(n470), .A2(n461), .ZN(n462) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(n462), .Z(n463) );
  NAND2_X1 U515 ( .A1(n463), .A2(n523), .ZN(n469) );
  NOR2_X1 U516 ( .A1(n527), .A2(n470), .ZN(n465) );
  XNOR2_X1 U517 ( .A(KEYINPUT103), .B(KEYINPUT26), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U519 ( .A(KEYINPUT102), .B(n466), .ZN(n570) );
  XNOR2_X1 U520 ( .A(KEYINPUT27), .B(KEYINPUT101), .ZN(n467) );
  XNOR2_X1 U521 ( .A(n467), .B(n478), .ZN(n522) );
  NOR2_X1 U522 ( .A1(n570), .A2(n522), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n469), .A2(n468), .ZN(n474) );
  INV_X1 U524 ( .A(n527), .ZN(n516) );
  XNOR2_X1 U525 ( .A(KEYINPUT28), .B(n470), .ZN(n528) );
  NAND2_X1 U526 ( .A1(n516), .A2(n528), .ZN(n471) );
  NOR2_X1 U527 ( .A1(n471), .A2(n522), .ZN(n472) );
  NOR2_X1 U528 ( .A1(n523), .A2(n472), .ZN(n473) );
  NOR2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n485) );
  NAND2_X1 U530 ( .A1(n475), .A2(n485), .ZN(n501) );
  OR2_X1 U531 ( .A1(n488), .A2(n501), .ZN(n482) );
  NOR2_X1 U532 ( .A1(n523), .A2(n482), .ZN(n476) );
  XOR2_X1 U533 ( .A(n476), .B(KEYINPUT34), .Z(n477) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  INV_X1 U535 ( .A(n478), .ZN(n514) );
  NOR2_X1 U536 ( .A1(n514), .A2(n482), .ZN(n479) );
  XOR2_X1 U537 ( .A(G8GAT), .B(n479), .Z(G1325GAT) );
  NOR2_X1 U538 ( .A1(n516), .A2(n482), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NOR2_X1 U541 ( .A1(n528), .A2(n482), .ZN(n483) );
  XOR2_X1 U542 ( .A(G22GAT), .B(n483), .Z(G1327GAT) );
  NAND2_X1 U543 ( .A1(n484), .A2(n485), .ZN(n486) );
  NOR2_X1 U544 ( .A1(n486), .A2(n549), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(KEYINPUT37), .ZN(n511) );
  NOR2_X1 U546 ( .A1(n511), .A2(n488), .ZN(n489) );
  XOR2_X1 U547 ( .A(KEYINPUT38), .B(n489), .Z(n496) );
  NOR2_X1 U548 ( .A1(n496), .A2(n523), .ZN(n491) );
  XNOR2_X1 U549 ( .A(KEYINPUT39), .B(KEYINPUT105), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U551 ( .A(G29GAT), .B(n492), .Z(G1328GAT) );
  NOR2_X1 U552 ( .A1(n514), .A2(n496), .ZN(n493) );
  XOR2_X1 U553 ( .A(G36GAT), .B(n493), .Z(G1329GAT) );
  NOR2_X1 U554 ( .A1(n516), .A2(n496), .ZN(n494) );
  XOR2_X1 U555 ( .A(KEYINPUT40), .B(n494), .Z(n495) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  XNOR2_X1 U557 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n498) );
  NOR2_X1 U558 ( .A1(n528), .A2(n496), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  NAND2_X1 U561 ( .A1(n560), .A2(n571), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT108), .ZN(n512) );
  NOR2_X1 U563 ( .A1(n501), .A2(n512), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(KEYINPUT109), .ZN(n507) );
  NOR2_X1 U565 ( .A1(n523), .A2(n507), .ZN(n503) );
  XOR2_X1 U566 ( .A(KEYINPUT42), .B(n503), .Z(n504) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U568 ( .A1(n514), .A2(n507), .ZN(n505) );
  XOR2_X1 U569 ( .A(G64GAT), .B(n505), .Z(G1333GAT) );
  NOR2_X1 U570 ( .A1(n516), .A2(n507), .ZN(n506) );
  XOR2_X1 U571 ( .A(G71GAT), .B(n506), .Z(G1334GAT) );
  NOR2_X1 U572 ( .A1(n528), .A2(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(n510), .ZN(G1335GAT) );
  OR2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n523), .A2(n518), .ZN(n513) );
  XOR2_X1 U578 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n518), .ZN(n515) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n515), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n516), .A2(n518), .ZN(n517) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n528), .A2(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(KEYINPUT114), .B(n526), .ZN(n541) );
  NAND2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U591 ( .A1(n541), .A2(n529), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n537), .A2(n542), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n530), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U595 ( .A1(n537), .A2(n560), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n536) );
  XOR2_X1 U598 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n534) );
  NAND2_X1 U599 ( .A1(n537), .A2(n549), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U603 ( .A1(n537), .A2(n552), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U605 ( .A(G134GAT), .B(n540), .Z(G1343GAT) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n544) );
  NOR2_X1 U607 ( .A1(n541), .A2(n570), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n542), .A2(n553), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n546) );
  NAND2_X1 U611 ( .A1(n553), .A2(n560), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT119), .Z(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n553), .A2(n549), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(KEYINPUT120), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(n551), .ZN(G1346GAT) );
  XOR2_X1 U618 ( .A(G162GAT), .B(KEYINPUT121), .Z(n555) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1347GAT) );
  NOR2_X1 U621 ( .A1(n566), .A2(n571), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT123), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(n557), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT126), .B(KEYINPUT125), .Z(n559) );
  XNOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n565) );
  INV_X1 U627 ( .A(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n580), .A2(n566), .ZN(n567) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n567), .Z(G1350GAT) );
  INV_X1 U633 ( .A(n568), .ZN(n569) );
  NOR2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n582) );
  INV_X1 U635 ( .A(n582), .ZN(n579) );
  NOR2_X1 U636 ( .A1(n579), .A2(n571), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n579), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n581), .Z(G1354GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n484), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

