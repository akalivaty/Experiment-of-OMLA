//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n210), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n232), .A2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n227), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n239), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n226), .ZN(new_n246));
  XOR2_X1   g0046(.A(KEYINPUT66), .B(G50), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  AOI21_X1  g0054(.A(G1), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n257), .A3(G274), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n259), .B1(G226), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT67), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G222), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n265), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n270), .A2(KEYINPUT67), .A3(G222), .A4(new_n271), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n270), .A2(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G223), .ZN(new_n278));
  INV_X1    g0078(.A(G77), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n277), .A2(new_n278), .B1(new_n279), .B2(new_n270), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n264), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G179), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n280), .B1(new_n274), .B2(new_n275), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n263), .B1(new_n287), .B2(new_n257), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n216), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n208), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(G150), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G50), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n208), .B1(new_n201), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n292), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n292), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n299), .B1(new_n207), .B2(G20), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n304), .A2(new_n305), .B1(new_n299), .B2(new_n303), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n286), .A2(new_n290), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n284), .A2(G190), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT9), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n307), .A2(KEYINPUT71), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT71), .B1(new_n307), .B2(new_n310), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n309), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  INV_X1    g0115(.A(new_n307), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n284), .A2(new_n315), .B1(KEYINPUT9), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT10), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n288), .A2(G200), .B1(new_n310), .B2(new_n307), .ZN(new_n319));
  INV_X1    g0119(.A(new_n311), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n312), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT10), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n319), .A2(new_n321), .A3(new_n322), .A4(new_n309), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n308), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n303), .A2(new_n220), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT12), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n296), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n279), .B2(new_n294), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(KEYINPUT11), .A3(new_n292), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n207), .A2(G20), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n304), .A2(G68), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n326), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT11), .B1(new_n328), .B2(new_n292), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n221), .B1(new_n261), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n257), .A2(KEYINPUT73), .A3(new_n260), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n259), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  AND2_X1   g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  NOR2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  OAI211_X1 g0142(.A(G226), .B(new_n271), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(G232), .B(G1698), .C1(new_n341), .C2(new_n342), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G97), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT72), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(KEYINPUT72), .A2(G33), .A3(G97), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n343), .A2(new_n344), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n283), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n339), .A2(new_n340), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n340), .B1(new_n339), .B2(new_n351), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT14), .B1(new_n354), .B2(new_n289), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(G179), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(G169), .C1(new_n352), .C2(new_n353), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(G200), .B1(new_n352), .B2(new_n353), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n337), .A2(new_n338), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(new_n351), .A3(new_n258), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT13), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n339), .A2(new_n340), .A3(new_n351), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(G190), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n360), .A2(new_n365), .A3(new_n334), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT74), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT74), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n360), .A2(new_n368), .A3(new_n365), .A4(new_n334), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n335), .A2(new_n359), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n270), .A2(G238), .A3(G1698), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n341), .A2(new_n342), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G107), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n371), .B(new_n373), .C1(new_n272), .C2(new_n227), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n283), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n259), .B1(G244), .B2(new_n262), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n375), .A2(KEYINPUT68), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT68), .B1(new_n375), .B2(new_n376), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n285), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT70), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n375), .A2(new_n376), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT68), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n375), .A2(KEYINPUT68), .A3(new_n376), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT70), .A3(new_n285), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n293), .A2(new_n297), .B1(new_n208), .B2(new_n279), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT15), .B(G87), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(new_n294), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n292), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n279), .B1(new_n207), .B2(G20), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n304), .A2(new_n393), .B1(new_n279), .B2(new_n303), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n386), .B2(G169), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n384), .A2(G200), .A3(new_n385), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n395), .B(KEYINPUT69), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n386), .A2(G190), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n388), .A2(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT76), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(KEYINPUT17), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n293), .B1(new_n207), .B2(G20), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(new_n304), .B1(new_n303), .B2(new_n293), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n292), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT7), .B1(new_n372), .B2(new_n208), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  NOR4_X1   g0210(.A1(new_n341), .A2(new_n342), .A3(new_n410), .A4(G20), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n226), .A2(new_n220), .ZN(new_n413));
  OAI21_X1  g0213(.A(G20), .B1(new_n413), .B2(new_n201), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n296), .A2(G159), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n408), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n417), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n407), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n257), .A2(G232), .A3(new_n260), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n258), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT75), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n278), .A2(new_n271), .ZN(new_n427));
  INV_X1    g0227(.A(G226), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G1698), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n427), .B(new_n429), .C1(new_n341), .C2(new_n342), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n257), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G190), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n258), .A2(new_n423), .A3(KEYINPUT75), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n426), .A2(new_n433), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n258), .A2(new_n423), .A3(KEYINPUT75), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT75), .B1(new_n258), .B2(new_n423), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n437), .A2(new_n438), .A3(new_n432), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n436), .B1(new_n439), .B2(G200), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n404), .B1(new_n422), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n410), .B1(new_n270), .B2(G20), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n372), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n220), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n419), .B1(new_n444), .B2(new_n416), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(new_n292), .A3(new_n421), .ZN(new_n446));
  XOR2_X1   g0246(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n447));
  AND4_X1   g0247(.A1(new_n446), .A2(new_n440), .A3(new_n406), .A4(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n441), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n439), .A2(new_n285), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(G169), .B2(new_n439), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT18), .B1(new_n422), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n446), .A2(new_n406), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n438), .A2(new_n432), .ZN(new_n454));
  AOI21_X1  g0254(.A(G169), .B1(new_n454), .B2(new_n435), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n437), .A2(new_n438), .A3(new_n432), .A4(G179), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT18), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n453), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n449), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n324), .A2(new_n370), .A3(new_n402), .A4(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n208), .B(G87), .C1(new_n341), .C2(new_n342), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT22), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT22), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n270), .A2(new_n465), .A3(new_n208), .A4(G87), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT24), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G116), .ZN(new_n469));
  OR3_X1    g0269(.A1(new_n469), .A2(KEYINPUT81), .A3(G20), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT81), .B1(new_n469), .B2(G20), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT23), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n208), .B2(G107), .ZN(new_n473));
  INV_X1    g0273(.A(G107), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(KEYINPUT23), .A3(G20), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n470), .A2(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n467), .A2(new_n468), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n468), .B1(new_n467), .B2(new_n476), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n292), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n207), .A2(G33), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n302), .A2(new_n480), .A3(new_n216), .A4(new_n291), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n303), .A2(KEYINPUT25), .A3(new_n474), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT25), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n302), .B2(G107), .ZN(new_n485));
  AOI22_X1  g0285(.A1(G107), .A2(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n223), .A2(new_n271), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n229), .A2(G1698), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n489), .C1(new_n341), .C2(new_n342), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G294), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n257), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n254), .A2(G1), .ZN(new_n493));
  AND2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  NOR2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(G264), .A3(new_n257), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT82), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT82), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n496), .A2(new_n499), .A3(G264), .A4(new_n257), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n492), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g0301(.A(KEYINPUT5), .B(G41), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(G274), .A3(new_n257), .A4(new_n493), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n490), .A2(new_n491), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n283), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n506), .A2(new_n497), .A3(new_n503), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n504), .A2(new_n315), .B1(new_n434), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT83), .B1(new_n487), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n486), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n467), .A2(new_n476), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT24), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n467), .A2(new_n468), .A3(new_n476), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n510), .B1(new_n514), .B2(new_n292), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT83), .ZN(new_n516));
  INV_X1    g0316(.A(new_n503), .ZN(new_n517));
  AOI211_X1 g0317(.A(new_n492), .B(new_n517), .C1(new_n498), .C2(new_n500), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n506), .A2(new_n497), .A3(new_n503), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n518), .A2(G200), .B1(G190), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n515), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n509), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n498), .A2(new_n500), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n523), .A2(G179), .A3(new_n503), .A4(new_n506), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n519), .A2(G169), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n408), .B1(new_n512), .B2(new_n513), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(new_n510), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n390), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(new_n302), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n481), .A2(new_n222), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n347), .A2(KEYINPUT19), .A3(new_n348), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n208), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT79), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT79), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n533), .A2(new_n536), .A3(new_n208), .ZN(new_n537));
  AND2_X1   g0337(.A1(KEYINPUT77), .A2(G97), .ZN(new_n538));
  NOR2_X1   g0338(.A1(KEYINPUT77), .A2(G97), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n222), .A3(new_n474), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n535), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(G20), .B1(new_n268), .B2(new_n269), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G68), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n540), .A2(new_n294), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(KEYINPUT19), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  AOI211_X1 g0348(.A(new_n531), .B(new_n532), .C1(new_n548), .C2(new_n292), .ZN(new_n549));
  OAI211_X1 g0349(.A(G244), .B(G1698), .C1(new_n341), .C2(new_n342), .ZN(new_n550));
  OAI211_X1 g0350(.A(G238), .B(new_n271), .C1(new_n341), .C2(new_n342), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n551), .A3(new_n469), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n283), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n207), .A2(G45), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n257), .A2(G250), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n257), .A2(G274), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(new_n554), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n553), .A2(new_n558), .A3(new_n434), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(new_n552), .B2(new_n283), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(G200), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n531), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n482), .A2(new_n530), .ZN(new_n563));
  XNOR2_X1  g0363(.A(KEYINPUT77), .B(G97), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n564), .A2(G87), .A3(G107), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n534), .B2(KEYINPUT79), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n546), .B1(new_n566), .B2(new_n537), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n562), .B(new_n563), .C1(new_n567), .C2(new_n408), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n553), .A2(new_n558), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(G179), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n560), .A2(G169), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n549), .A2(new_n561), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT6), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n228), .A2(new_n474), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(new_n204), .ZN(new_n576));
  OAI211_X1 g0376(.A(KEYINPUT6), .B(new_n474), .C1(new_n538), .C2(new_n539), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(G20), .B1(G77), .B2(new_n296), .ZN(new_n579));
  OAI21_X1  g0379(.A(G107), .B1(new_n409), .B2(new_n411), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n292), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n303), .A2(new_n228), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n481), .B2(new_n228), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(G244), .B(new_n271), .C1(new_n341), .C2(new_n342), .ZN(new_n587));
  XNOR2_X1  g0387(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n270), .A2(G250), .A3(G1698), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G283), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n283), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n496), .A2(new_n257), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n503), .B1(new_n595), .B2(new_n229), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n289), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n596), .B1(new_n593), .B2(new_n283), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n285), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n586), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n584), .B1(new_n581), .B2(new_n292), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(G190), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n603), .B(new_n604), .C1(new_n315), .C2(new_n600), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n573), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT21), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n208), .B(new_n592), .C1(new_n540), .C2(G33), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT20), .ZN(new_n609));
  INV_X1    g0409(.A(G116), .ZN(new_n610));
  AOI22_X1  g0410(.A1(KEYINPUT80), .A2(new_n609), .B1(new_n610), .B2(G20), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n292), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n609), .A2(KEYINPUT80), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n608), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n592), .A2(new_n208), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n564), .B2(new_n267), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n614), .B1(new_n618), .B2(new_n612), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n302), .A2(new_n610), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n482), .B2(new_n610), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n616), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n271), .A2(G264), .ZN(new_n623));
  NOR2_X1   g0423(.A1(G257), .A2(G1698), .ZN(new_n624));
  OAI22_X1  g0424(.A1(new_n623), .A2(new_n624), .B1(new_n341), .B2(new_n342), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n625), .B(new_n283), .C1(G303), .C2(new_n270), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n496), .A2(G270), .A3(new_n257), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n503), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G169), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n607), .B1(new_n622), .B2(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(G179), .A2(new_n626), .A3(new_n503), .A4(new_n627), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n616), .A2(new_n619), .A3(new_n621), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(KEYINPUT21), .A3(new_n628), .A4(G169), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n630), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n632), .B1(G200), .B2(new_n628), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n434), .B2(new_n628), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NOR4_X1   g0438(.A1(new_n462), .A2(new_n529), .A3(new_n606), .A4(new_n638), .ZN(G372));
  AND3_X1   g0439(.A1(new_n453), .A2(new_n457), .A3(new_n458), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n458), .B1(new_n453), .B2(new_n457), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n359), .A2(new_n335), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n396), .B1(new_n381), .B2(new_n387), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n366), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n646), .B2(new_n449), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n318), .A2(new_n323), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n308), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n462), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n568), .A2(new_n572), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n531), .B1(new_n548), .B2(new_n292), .ZN(new_n652));
  INV_X1    g0452(.A(new_n532), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(new_n561), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n651), .A2(new_n602), .A3(new_n605), .A4(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n634), .A2(new_n633), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n528), .A2(new_n656), .A3(new_n630), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n522), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n651), .A2(new_n654), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n602), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n408), .B1(new_n579), .B2(new_n580), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n662), .A2(new_n584), .B1(new_n600), .B2(G169), .ZN(new_n663));
  INV_X1    g0463(.A(new_n601), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n573), .A2(KEYINPUT26), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n658), .A2(new_n667), .A3(new_n651), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n650), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n649), .A2(new_n669), .ZN(G369));
  INV_X1    g0470(.A(new_n635), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n529), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n528), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n678), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n622), .A2(new_n678), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n671), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n638), .B2(new_n683), .ZN(new_n685));
  XOR2_X1   g0485(.A(KEYINPUT84), .B(G330), .Z(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n681), .B1(new_n509), .B2(new_n521), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n487), .A2(new_n677), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n688), .A2(new_n689), .B1(new_n681), .B2(new_n677), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n682), .B1(new_n687), .B2(new_n690), .ZN(G399));
  NAND2_X1  g0491(.A1(new_n211), .A2(new_n253), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n207), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n541), .A2(G116), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n694), .A2(new_n695), .B1(new_n215), .B2(new_n693), .ZN(new_n696));
  XOR2_X1   g0496(.A(new_n696), .B(KEYINPUT28), .Z(new_n697));
  NAND4_X1  g0497(.A1(new_n600), .A2(new_n631), .A3(new_n501), .A4(new_n560), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n501), .A2(new_n560), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(KEYINPUT30), .A3(new_n600), .A4(new_n631), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n628), .A2(new_n285), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n504), .A2(new_n703), .A3(new_n598), .A4(new_n569), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n700), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT31), .B1(new_n705), .B2(new_n677), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n638), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n688), .A2(new_n709), .A3(new_n655), .A4(new_n678), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n711), .A2(new_n686), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n668), .A2(new_n678), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n509), .A2(new_n521), .B1(new_n635), .B2(new_n528), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n716), .A2(new_n655), .B1(new_n568), .B2(new_n572), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n661), .A2(new_n666), .A3(KEYINPUT85), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT85), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n573), .A2(new_n719), .A3(KEYINPUT26), .A4(new_n665), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .A3(new_n678), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n712), .B1(new_n715), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n697), .B1(new_n723), .B2(G1), .ZN(G364));
  NAND2_X1  g0524(.A1(new_n208), .A2(G13), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT86), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G45), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n727), .A2(KEYINPUT87), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(KEYINPUT87), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n694), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n685), .B2(new_n686), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n686), .B2(new_n685), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n211), .A2(new_n270), .ZN(new_n736));
  INV_X1    g0536(.A(G355), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n736), .A2(new_n737), .B1(G116), .B2(new_n211), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n211), .A2(new_n372), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n254), .B2(new_n215), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT88), .Z(new_n741));
  NAND2_X1  g0541(.A1(new_n248), .A2(G45), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n738), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n216), .B1(G20), .B2(new_n289), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n733), .B1(new_n743), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n747), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n208), .B1(new_n752), .B2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n228), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n208), .A2(G190), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n752), .ZN(new_n756));
  INV_X1    g0556(.A(G159), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT89), .B(KEYINPUT32), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n208), .A2(new_n285), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n434), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n754), .B(new_n760), .C1(G50), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n208), .A2(new_n434), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n315), .A2(G179), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n270), .B1(new_n767), .B2(new_n222), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT90), .Z(new_n769));
  NAND3_X1  g0569(.A1(new_n761), .A2(new_n434), .A3(G200), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n770), .A2(KEYINPUT91), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(KEYINPUT91), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n769), .B1(new_n774), .B2(G68), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n766), .A2(new_n755), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G107), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n285), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n765), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n755), .A2(new_n779), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G58), .A2(new_n781), .B1(new_n783), .B2(G77), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n764), .A2(new_n775), .A3(new_n778), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n774), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G322), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n780), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G303), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n767), .A2(new_n790), .B1(new_n782), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n756), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n789), .B(new_n792), .C1(G329), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n763), .A2(G326), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n372), .B1(new_n776), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n753), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(G294), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n787), .A2(new_n794), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n751), .B1(new_n785), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n750), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n746), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n685), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n735), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  NAND3_X1  g0606(.A1(new_n388), .A2(new_n397), .A3(new_n678), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n377), .A2(new_n378), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n398), .B(new_n399), .C1(new_n808), .C2(new_n434), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n395), .A2(new_n677), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n807), .B1(new_n811), .B2(new_n645), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n713), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT92), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n677), .B1(new_n717), .B2(new_n667), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT93), .B1(new_n815), .B2(new_n402), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n668), .A2(KEYINPUT93), .A3(new_n402), .A4(new_n678), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n712), .B1(new_n814), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n733), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n814), .A2(new_n820), .A3(new_n712), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n747), .A2(new_n744), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n732), .B1(new_n279), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n767), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n270), .B(new_n754), .C1(G107), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n763), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n790), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n773), .A2(new_n796), .ZN(new_n831));
  INV_X1    g0631(.A(G294), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n780), .A2(new_n832), .B1(new_n776), .B2(new_n222), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n782), .A2(new_n610), .B1(new_n756), .B2(new_n791), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n830), .A2(new_n831), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G143), .A2(new_n781), .B1(new_n783), .B2(G159), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n837), .B2(new_n829), .C1(new_n773), .C2(new_n295), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT34), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n270), .B1(new_n767), .B2(new_n299), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n776), .A2(new_n220), .B1(new_n756), .B2(new_n841), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n840), .B(new_n842), .C1(G58), .C2(new_n798), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n835), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n807), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n388), .A2(new_n397), .B1(new_n809), .B2(new_n810), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n826), .B1(new_n751), .B2(new_n844), .C1(new_n847), .C2(new_n745), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n824), .A2(new_n848), .ZN(G384));
  INV_X1    g0649(.A(KEYINPUT39), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n422), .A2(new_n675), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n449), .B2(new_n460), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT37), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n440), .A2(new_n446), .A3(new_n406), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n422), .B2(new_n451), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n855), .B2(new_n851), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n453), .A2(new_n457), .ZN(new_n857));
  INV_X1    g0657(.A(new_n675), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n453), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n857), .A2(new_n859), .A3(KEYINPUT37), .A4(new_n854), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n852), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT97), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n854), .B1(new_n403), .B2(KEYINPUT17), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n422), .A2(new_n440), .A3(new_n447), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n859), .B1(new_n642), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n856), .A2(new_n860), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT97), .B(new_n862), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n867), .A2(new_n868), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT98), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT38), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n852), .A2(KEYINPUT38), .A3(new_n856), .A4(new_n860), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT98), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n850), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n862), .B1(new_n867), .B2(new_n868), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT96), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(KEYINPUT96), .B(new_n862), .C1(new_n867), .C2(new_n868), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n872), .A2(KEYINPUT95), .A3(KEYINPUT38), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT95), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n875), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n644), .A2(new_n678), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n878), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n807), .B(KEYINPUT94), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n816), .B2(new_n818), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n883), .A2(new_n887), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n334), .A2(new_n678), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n366), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n643), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n359), .B1(new_n367), .B2(new_n369), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n899), .B1(new_n900), .B2(new_n897), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n894), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n642), .A2(new_n858), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n891), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT99), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT99), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n891), .A2(new_n902), .A3(new_n907), .A4(new_n904), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n647), .A2(new_n648), .ZN(new_n910));
  INV_X1    g0710(.A(new_n308), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n722), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n650), .B1(new_n815), .B2(KEYINPUT29), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT100), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n462), .B1(new_n713), .B2(new_n714), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT100), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n917), .A3(new_n722), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n912), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n909), .B(new_n919), .Z(new_n920));
  INV_X1    g0720(.A(KEYINPUT101), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n711), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n367), .A2(new_n369), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n896), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n812), .B1(new_n926), .B2(new_n899), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n708), .A2(new_n710), .A3(KEYINPUT101), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n922), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT102), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT102), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n922), .A2(new_n927), .A3(new_n931), .A4(new_n928), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n895), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT40), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n929), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(KEYINPUT40), .C1(new_n871), .C2(new_n877), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n922), .A2(new_n650), .A3(new_n928), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n686), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n938), .B2(new_n939), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n920), .A2(new_n941), .B1(new_n207), .B2(new_n726), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n920), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n578), .A2(KEYINPUT35), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n578), .A2(KEYINPUT35), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n944), .A2(G116), .A3(new_n217), .A4(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT36), .Z(new_n947));
  OR3_X1    g0747(.A1(new_n214), .A2(new_n279), .A3(new_n413), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n299), .A2(G68), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n207), .B(G13), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  OR3_X1    g0750(.A1(new_n943), .A2(new_n947), .A3(new_n950), .ZN(G367));
  NOR2_X1   g0751(.A1(new_n730), .A2(new_n207), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n602), .B(new_n605), .C1(new_n603), .C2(new_n678), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n602), .B2(new_n678), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n682), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT45), .Z(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT44), .B1(new_n682), .B2(new_n954), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n682), .A2(KEYINPUT44), .A3(new_n954), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n687), .A2(new_n690), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(KEYINPUT109), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n956), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n959), .A2(KEYINPUT109), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT108), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n687), .A2(new_n964), .B1(new_n680), .B2(KEYINPUT107), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT107), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n690), .B2(new_n679), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n965), .B1(new_n680), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n687), .A2(new_n964), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n723), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n963), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n973), .A2(new_n723), .ZN(new_n974));
  XNOR2_X1  g0774(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n692), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n952), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n549), .A2(new_n678), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n651), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n573), .B2(new_n978), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT103), .Z(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT104), .Z(new_n984));
  OR2_X1    g0784(.A1(new_n953), .A2(new_n528), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n677), .B1(new_n985), .B2(new_n602), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n680), .A2(new_n954), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT105), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n986), .B1(new_n988), .B2(KEYINPUT42), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(KEYINPUT42), .B2(new_n988), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n984), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n984), .A2(new_n992), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n959), .A2(new_n954), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n996), .B(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n977), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n981), .A2(new_n746), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n239), .A2(new_n739), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n748), .B1(new_n211), .B2(new_n390), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n733), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n767), .A2(new_n610), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n829), .A2(new_n791), .B1(KEYINPUT46), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(KEYINPUT46), .B2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n774), .A2(G294), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n776), .A2(new_n540), .B1(new_n756), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G303), .B2(new_n781), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n372), .B1(new_n782), .B2(new_n796), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G107), .B2(new_n798), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1007), .A2(new_n1008), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n270), .B1(new_n756), .B2(new_n837), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n777), .A2(G77), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n299), .B2(new_n782), .C1(new_n226), .C2(new_n767), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1015), .B(new_n1017), .C1(G143), .C2(new_n763), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n757), .B2(new_n773), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n753), .A2(new_n220), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G150), .B2(new_n781), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT110), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1014), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT47), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1004), .B1(new_n1024), .B2(new_n747), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1001), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1000), .A2(new_n1026), .ZN(G387));
  INV_X1    g0827(.A(new_n952), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n690), .A2(new_n746), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n695), .A2(new_n736), .B1(G107), .B2(new_n211), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n695), .B(new_n254), .C1(new_n220), .C2(new_n279), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT111), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  OAI21_X1  g0834(.A(KEYINPUT50), .B1(new_n293), .B2(G50), .ZN(new_n1035));
  OR3_X1    g0835(.A1(new_n293), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n739), .B1(new_n243), .B2(G45), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1030), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n733), .B1(new_n1039), .B2(new_n749), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n773), .A2(new_n293), .B1(new_n220), .B2(new_n782), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT113), .Z(new_n1042));
  NAND2_X1  g0842(.A1(new_n777), .A2(G97), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(KEYINPUT112), .B(G150), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n299), .B2(new_n780), .C1(new_n756), .C2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n753), .A2(new_n390), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n270), .B1(new_n279), .B2(new_n767), .C1(new_n829), .C2(new_n757), .ZN(new_n1047));
  OR4_X1    g0847(.A1(new_n1042), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G317), .A2(new_n781), .B1(new_n783), .B2(G303), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n788), .B2(new_n829), .C1(new_n773), .C2(new_n791), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n827), .A2(G294), .B1(new_n798), .B2(G283), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT49), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(KEYINPUT114), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n270), .B1(new_n793), .B2(G326), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n610), .C2(new_n776), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1056), .A2(KEYINPUT114), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1048), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1040), .B1(new_n1061), .B2(new_n747), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n970), .A2(new_n1028), .B1(new_n1029), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n971), .A2(new_n693), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n970), .A2(new_n723), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1066), .A2(KEYINPUT115), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(KEYINPUT115), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(G393));
  NAND2_X1  g0870(.A1(new_n973), .A2(new_n693), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT120), .ZN(new_n1072));
  OR3_X1    g0872(.A1(new_n963), .A2(new_n1072), .A3(new_n972), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1072), .B1(new_n963), .B2(new_n972), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n963), .A2(new_n1028), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n748), .B1(new_n211), .B2(new_n540), .C1(new_n251), .C2(new_n739), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT116), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n733), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n767), .A2(new_n796), .B1(new_n756), .B2(new_n788), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT117), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n372), .B(new_n778), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1083), .B2(new_n1082), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT118), .Z(new_n1086));
  AOI22_X1  g0886(.A1(new_n763), .A2(G317), .B1(new_n781), .B2(G311), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT52), .Z(new_n1088));
  OAI22_X1  g0888(.A1(new_n782), .A2(new_n832), .B1(new_n753), .B2(new_n610), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n774), .B2(G303), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1091), .A2(KEYINPUT119), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n763), .A2(G150), .B1(new_n781), .B2(G159), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT51), .Z(new_n1094));
  NAND2_X1  g0894(.A1(new_n774), .A2(G50), .ZN(new_n1095));
  INV_X1    g0895(.A(G143), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n782), .A2(new_n293), .B1(new_n756), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G68), .B2(new_n827), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n753), .A2(new_n279), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n372), .B(new_n1099), .C1(G87), .C2(new_n777), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1094), .A2(new_n1095), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1091), .A2(KEYINPUT119), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1092), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1081), .B1(new_n1103), .B2(new_n747), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n803), .B2(new_n954), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1076), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1075), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(G390));
  INV_X1    g0908(.A(KEYINPUT121), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n922), .A2(new_n650), .A3(G330), .A4(new_n928), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n916), .A2(new_n917), .A3(new_n722), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n917), .B1(new_n916), .B2(new_n722), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n649), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n922), .A2(new_n927), .A3(G330), .A4(new_n928), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n711), .A2(new_n686), .A3(new_n847), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n901), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n922), .A2(G330), .A3(new_n847), .A4(new_n928), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n1116), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n711), .A2(new_n901), .A3(new_n847), .A4(new_n686), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n846), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n658), .A2(new_n651), .A3(new_n720), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n718), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n678), .B(new_n1122), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1121), .A2(new_n1125), .A3(new_n807), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n894), .A2(new_n1118), .B1(new_n1120), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1109), .B1(new_n1113), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n894), .A2(new_n1118), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1120), .A2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1131), .A2(KEYINPUT121), .A3(new_n919), .A4(new_n1110), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n878), .A2(new_n888), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n487), .A2(new_n508), .A3(KEYINPUT83), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n516), .B1(new_n515), .B2(new_n520), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n657), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n651), .B1(new_n1137), .B2(new_n606), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT26), .B1(new_n573), .B2(new_n665), .ZN(new_n1139));
  AND4_X1   g0939(.A1(KEYINPUT26), .A2(new_n665), .A3(new_n651), .A4(new_n654), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n402), .B(new_n678), .C1(new_n1138), .C2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT93), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n892), .B1(new_n1144), .B2(new_n817), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n889), .B1(new_n1145), .B2(new_n1116), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1134), .A2(new_n1146), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n874), .A2(new_n876), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT97), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n879), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n869), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n890), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1125), .A2(new_n807), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n901), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1147), .A2(new_n1155), .A3(new_n1121), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1134), .A2(new_n1146), .B1(new_n1154), .B2(new_n1152), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n1114), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n692), .B1(new_n1133), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1121), .ZN(new_n1160));
  AOI221_X4 g0960(.A(new_n1160), .B1(new_n1152), .B2(new_n1154), .C1(new_n1134), .C2(new_n1146), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1114), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1159), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1028), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1134), .A2(new_n744), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n732), .B1(new_n293), .B2(new_n825), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT54), .B(G143), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n270), .B1(new_n782), .B2(new_n1170), .C1(new_n829), .C2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G159), .B2(new_n798), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n774), .A2(G137), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n767), .A2(new_n1044), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT53), .ZN(new_n1176));
  INV_X1    g0976(.A(G125), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n780), .A2(new_n841), .B1(new_n756), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G50), .B2(new_n777), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n372), .B1(new_n767), .B2(new_n222), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1099), .B(new_n1181), .C1(G283), .C2(new_n763), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n780), .A2(new_n610), .B1(new_n776), .B2(new_n220), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n782), .A2(new_n540), .B1(new_n756), .B2(new_n832), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1182), .B(new_n1185), .C1(new_n474), .C2(new_n773), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1180), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1168), .B(new_n1169), .C1(new_n751), .C2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1166), .A2(new_n1167), .A3(new_n1188), .ZN(G378));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n316), .A2(new_n675), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n324), .B(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1192), .B(new_n1193), .Z(new_n1194));
  AOI22_X1  g0994(.A1(new_n883), .A2(new_n887), .B1(new_n929), .B2(KEYINPUT102), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT40), .B1(new_n1195), .B2(new_n932), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n937), .A2(G330), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1194), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n935), .A2(G330), .A3(new_n937), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n909), .A2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n906), .A2(new_n1198), .A3(new_n1200), .A4(new_n908), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1113), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1190), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1113), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1133), .B2(new_n1158), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1208), .A2(KEYINPUT57), .A3(new_n1203), .A4(new_n1202), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n693), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1202), .A2(new_n1028), .A3(new_n1203), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n270), .A2(G41), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G50), .B(new_n1212), .C1(new_n267), .C2(new_n253), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n774), .A2(G97), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n780), .A2(new_n474), .B1(new_n782), .B2(new_n390), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n776), .A2(new_n226), .B1(new_n756), .B2(new_n796), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n763), .A2(G116), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1212), .B1(new_n279), .B2(new_n767), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(new_n1020), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1214), .A2(new_n1217), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT58), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1213), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n829), .A2(new_n1177), .B1(new_n837), .B2(new_n782), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G150), .B2(new_n798), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1171), .A2(new_n780), .B1(new_n767), .B2(new_n1170), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT122), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1225), .B(new_n1227), .C1(new_n841), .C2(new_n773), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n267), .B(new_n253), .C1(new_n776), .C2(new_n757), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G124), .B2(new_n793), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1223), .B1(new_n1222), .B2(new_n1221), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n747), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n732), .B1(new_n299), .B2(new_n825), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n1199), .C2(new_n745), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT123), .Z(new_n1238));
  NAND2_X1  g1038(.A1(new_n1211), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1210), .A2(new_n1240), .ZN(G375));
  AOI21_X1  g1041(.A(new_n372), .B1(new_n777), .B2(G58), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n299), .B2(new_n753), .C1(new_n829), .C2(new_n841), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n773), .A2(new_n1170), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n767), .A2(new_n757), .B1(new_n756), .B2(new_n1171), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n780), .A2(new_n837), .B1(new_n782), .B2(new_n295), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n773), .A2(new_n610), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n763), .A2(G294), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1046), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1249), .A2(new_n372), .A3(new_n1016), .A4(new_n1250), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n767), .A2(new_n228), .B1(new_n756), .B2(new_n790), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n780), .A2(new_n796), .B1(new_n782), .B2(new_n474), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(new_n1248), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n747), .B1(new_n1247), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n732), .B1(new_n220), .B2(new_n825), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(new_n901), .C2(new_n745), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1127), .B2(new_n952), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1207), .A2(KEYINPUT124), .A3(new_n1131), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT124), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1113), .B2(new_n1127), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  OR2_X1    g1064(.A1(new_n1164), .A2(new_n976), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1259), .B1(new_n1264), .B2(new_n1265), .ZN(G381));
  NAND3_X1  g1066(.A1(new_n1068), .A2(new_n805), .A3(new_n1069), .ZN(new_n1267));
  NOR4_X1   g1067(.A1(G387), .A2(G390), .A3(G384), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1167), .A2(new_n1188), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1165), .B2(new_n1159), .ZN(new_n1270));
  INV_X1    g1070(.A(G375), .ZN(new_n1271));
  INV_X1    g1071(.A(G381), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1268), .A2(new_n1270), .A3(new_n1271), .A4(new_n1272), .ZN(G407));
  NAND2_X1  g1073(.A1(new_n676), .A2(G213), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1271), .A2(new_n1270), .A3(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(G407), .A2(G213), .A3(new_n1276), .ZN(G409));
  NAND2_X1  g1077(.A1(G387), .A2(new_n1107), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(G390), .A2(new_n1000), .A3(new_n1026), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G393), .A2(G396), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1267), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1280), .B(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1210), .A2(G378), .A3(new_n1240), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1204), .A2(new_n1205), .A3(new_n976), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1270), .B1(new_n1285), .B2(new_n1239), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1275), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n1127), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n693), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1133), .A2(KEYINPUT60), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1290), .B2(new_n1263), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(G384), .A3(new_n1259), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n824), .B(new_n848), .C1(new_n1291), .C2(new_n1258), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1287), .A2(KEYINPUT62), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT62), .B1(new_n1287), .B2(new_n1296), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1287), .A2(new_n1296), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1299), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1274), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1275), .A2(G2897), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1293), .A2(new_n1294), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1306), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT61), .B1(new_n1305), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1303), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1283), .B1(new_n1300), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1282), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1280), .B(new_n1313), .ZN(new_n1314));
  XOR2_X1   g1114(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1315));
  NAND2_X1  g1115(.A1(new_n1301), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1287), .A2(KEYINPUT63), .A3(new_n1296), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1314), .A2(new_n1316), .A3(new_n1317), .A4(new_n1310), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1312), .A2(new_n1318), .ZN(G405));
  OAI21_X1  g1119(.A(new_n1295), .B1(new_n1271), .B2(G378), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1296), .A2(new_n1270), .A3(G375), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT127), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1284), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1320), .A2(new_n1321), .A3(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1323), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1283), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1326), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1314), .A2(new_n1328), .A3(new_n1324), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1327), .A2(new_n1329), .ZN(G402));
endmodule


