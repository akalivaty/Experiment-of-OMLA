//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  XOR2_X1   g030(.A(KEYINPUT66), .B(KEYINPUT67), .Z(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n454), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(G2106), .A2(new_n454), .B1(new_n458), .B2(G567), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n464), .B1(KEYINPUT3), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n463), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n462), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(new_n473), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n471), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  AOI211_X1 g053(.A(KEYINPUT68), .B(new_n478), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  NOR3_X1   g054(.A1(new_n470), .A2(new_n477), .A3(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n462), .A2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n472), .B1(new_n481), .B2(new_n464), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n482), .A2(new_n463), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(new_n478), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(new_n478), .B2(G112), .ZN(new_n487));
  OAI22_X1  g062(.A1(new_n484), .A2(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n483), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n482), .A2(new_n463), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(new_n478), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n488), .B1(G124), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT71), .ZN(G162));
  NAND4_X1  g070(.A1(new_n472), .A2(new_n473), .A3(G138), .A4(new_n478), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n465), .A2(G2105), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n496), .A2(new_n497), .B1(G102), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT4), .A2(G138), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n482), .A2(new_n478), .A3(new_n463), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G126), .B(new_n463), .C1(new_n466), .C2(new_n467), .ZN(new_n503));
  NAND2_X1  g078(.A1(G114), .A2(G2104), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n478), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT73), .A3(G62), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(new_n510), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n512), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT72), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n522), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(KEYINPUT6), .ZN(new_n528));
  NOR3_X1   g103(.A1(new_n527), .A2(new_n515), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G88), .ZN(new_n530));
  INV_X1    g105(.A(G50), .ZN(new_n531));
  INV_X1    g106(.A(new_n528), .ZN(new_n532));
  OAI211_X1 g107(.A(G543), .B(new_n532), .C1(new_n519), .C2(new_n522), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n530), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n521), .A2(new_n534), .ZN(G166));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n529), .A2(G89), .B1(new_n511), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  INV_X1    g114(.A(new_n533), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n537), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT74), .ZN(G168));
  AOI22_X1  g118(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  INV_X1    g119(.A(new_n519), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n529), .A2(G90), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n540), .A2(G52), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(new_n540), .A2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n529), .A2(G81), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n515), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(new_n519), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n551), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  NOR2_X1   g139(.A1(new_n527), .A2(new_n528), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n565), .A2(new_n566), .A3(G53), .A4(G543), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n533), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n529), .A2(G91), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(new_n523), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(G299));
  XOR2_X1   g149(.A(new_n542), .B(KEYINPUT74), .Z(G286));
  OAI211_X1 g150(.A(new_n520), .B(new_n530), .C1(new_n531), .C2(new_n533), .ZN(G303));
  INV_X1    g151(.A(G74), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n523), .B1(new_n515), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n529), .B2(G87), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n540), .A2(G49), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(new_n540), .A2(G48), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n529), .A2(G86), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n508), .A2(new_n510), .A3(G61), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n508), .A2(new_n510), .A3(KEYINPUT75), .A4(G61), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n589), .A2(KEYINPUT76), .A3(new_n519), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT76), .B1(new_n589), .B2(new_n519), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n582), .B(new_n583), .C1(new_n590), .C2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n540), .A2(G47), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n529), .A2(G85), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n593), .B(new_n594), .C1(new_n545), .C2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n529), .A2(G92), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT10), .Z(new_n599));
  AOI22_X1  g174(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G54), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n600), .A2(new_n523), .B1(new_n533), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(new_n605), .B2(G868), .ZN(G284));
  XOR2_X1   g181(.A(G284), .B(KEYINPUT78), .Z(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  XOR2_X1   g183(.A(G299), .B(KEYINPUT79), .Z(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(G868), .B2(new_n609), .ZN(G297));
  OAI21_X1  g185(.A(new_n608), .B1(G868), .B2(new_n609), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT80), .Z(G148));
  NAND2_X1  g189(.A1(new_n605), .A2(new_n612), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  OR3_X1    g192(.A1(new_n616), .A2(KEYINPUT81), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT81), .B1(new_n616), .B2(new_n617), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n618), .B(new_n619), .C1(G868), .C2(new_n558), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g196(.A(KEYINPUT3), .B(G2104), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n498), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2100), .Z(new_n626));
  INV_X1    g201(.A(G135), .ZN(new_n627));
  NOR2_X1   g202(.A1(G99), .A2(G2105), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(new_n478), .B2(G111), .ZN(new_n629));
  OAI22_X1  g204(.A1(new_n484), .A2(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G123), .B2(new_n493), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n626), .A2(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XOR2_X1   g210(.A(G2443), .B(G2446), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT15), .B(G2435), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n639), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G14), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2067), .B(G2678), .Z(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT17), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n656), .B(new_n657), .C1(new_n655), .C2(new_n651), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n657), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2096), .B(G2100), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n663), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  AOI22_X1  g244(.A1(new_n667), .A2(KEYINPUT20), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n671), .A2(new_n663), .A3(new_n666), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n670), .B(new_n672), .C1(KEYINPUT20), .C2(new_n667), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1986), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1991), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G229));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G22), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G166), .B2(new_n680), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT85), .B(G1971), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(G6), .B(G305), .S(G16), .Z(new_n685));
  XOR2_X1   g260(.A(KEYINPUT32), .B(G1981), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G1976), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n680), .A2(G23), .ZN(new_n689));
  INV_X1    g264(.A(G288), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(new_n680), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(KEYINPUT33), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(KEYINPUT33), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n688), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(KEYINPUT33), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(G1976), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n684), .B(new_n687), .C1(new_n694), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT84), .B(KEYINPUT34), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n680), .A2(G24), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G290), .B2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G1986), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G25), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n493), .A2(G119), .ZN(new_n706));
  INV_X1    g281(.A(G131), .ZN(new_n707));
  NOR2_X1   g282(.A1(G95), .A2(G2105), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(new_n478), .B2(G107), .ZN(new_n709));
  OAI22_X1  g284(.A1(new_n484), .A2(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n705), .B1(new_n711), .B2(new_n704), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT35), .B(G1991), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT82), .Z(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT83), .Z(new_n715));
  OR2_X1    g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n712), .A2(new_n715), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n716), .B(new_n717), .C1(new_n702), .C2(new_n701), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n697), .B2(new_n698), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n699), .A2(new_n703), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT86), .B(KEYINPUT36), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n704), .A2(G26), .ZN(new_n724));
  INV_X1    g299(.A(G104), .ZN(new_n725));
  AND3_X1   g300(.A1(new_n725), .A2(new_n478), .A3(KEYINPUT88), .ZN(new_n726));
  AOI21_X1  g301(.A(KEYINPUT88), .B1(new_n725), .B2(new_n478), .ZN(new_n727));
  OAI221_X1 g302(.A(G2104), .B1(G116), .B2(new_n478), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n484), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G140), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n493), .A2(new_n731), .A3(G128), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n493), .B2(G128), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n728), .B(new_n730), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n724), .B1(new_n735), .B2(new_n704), .ZN(new_n736));
  MUX2_X1   g311(.A(new_n724), .B(new_n736), .S(KEYINPUT28), .Z(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(G2067), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n493), .A2(G129), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n498), .A2(G105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT92), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n729), .B2(G141), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n739), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G29), .B2(G32), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n704), .A2(G33), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n498), .A2(G103), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n622), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n757));
  INV_X1    g332(.A(G139), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n756), .B1(new_n478), .B2(new_n757), .C1(new_n484), .C2(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT90), .Z(new_n760));
  AOI21_X1  g335(.A(new_n753), .B1(new_n760), .B2(G29), .ZN(new_n761));
  INV_X1    g336(.A(G2072), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n749), .A2(new_n751), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n752), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n680), .A2(G19), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n558), .B2(new_n680), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(G1341), .ZN(new_n768));
  INV_X1    g343(.A(G34), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(KEYINPUT24), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(KEYINPUT24), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G160), .B2(new_n704), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n768), .B1(G2084), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G5), .A2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G171), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G2078), .ZN(new_n779));
  NOR2_X1   g354(.A1(G27), .A2(G29), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G164), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n776), .B1(G1961), .B2(new_n778), .C1(new_n779), .C2(new_n782), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT31), .B(G11), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n778), .A2(G1961), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n767), .A2(G1341), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n704), .B1(new_n787), .B2(G28), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n787), .B2(G28), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n631), .B2(G29), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n782), .A2(new_n779), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n785), .A2(new_n786), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NOR4_X1   g367(.A1(new_n765), .A2(new_n783), .A3(new_n784), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n680), .A2(G20), .ZN(new_n794));
  INV_X1    g369(.A(G299), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n680), .ZN(new_n796));
  MUX2_X1   g371(.A(new_n794), .B(new_n796), .S(KEYINPUT23), .Z(new_n797));
  XOR2_X1   g372(.A(KEYINPUT98), .B(G1956), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n775), .A2(G2084), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT97), .Z(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n761), .A2(new_n762), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT91), .Z(new_n804));
  NAND3_X1  g379(.A1(new_n793), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n704), .A2(G35), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G162), .B2(new_n704), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT29), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(KEYINPUT29), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G2090), .ZN(new_n811));
  NAND2_X1  g386(.A1(G168), .A2(G16), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(KEYINPUT94), .C1(G16), .C2(G21), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(KEYINPUT94), .B2(new_n812), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT96), .B(G1966), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT95), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(G2090), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n808), .A2(new_n818), .A3(new_n809), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n737), .A2(G2067), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n811), .A2(new_n817), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n680), .A2(G4), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n605), .B2(new_n680), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1348), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n805), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n723), .A2(new_n738), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(G311));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n723), .A2(KEYINPUT99), .A3(new_n825), .A4(new_n738), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(G150));
  NAND2_X1  g406(.A1(new_n599), .A2(new_n604), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(new_n612), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(G80), .A2(G543), .ZN(new_n836));
  INV_X1    g411(.A(G67), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n515), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n519), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT100), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n529), .A2(G93), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n540), .A2(G55), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n557), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n558), .A2(KEYINPUT101), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n843), .A2(new_n845), .A3(new_n557), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n835), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT102), .B(G860), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT103), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n843), .A2(new_n853), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(G162), .B(new_n631), .ZN(new_n859));
  INV_X1    g434(.A(G142), .ZN(new_n860));
  NOR2_X1   g435(.A1(G106), .A2(G2105), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(new_n478), .B2(G118), .ZN(new_n862));
  OAI22_X1  g437(.A1(new_n484), .A2(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(G130), .B2(new_n493), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(G160), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n859), .B(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n734), .A2(G164), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n734), .A2(G164), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n746), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n732), .A2(new_n733), .ZN(new_n870));
  INV_X1    g445(.A(G164), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n728), .A4(new_n730), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n734), .A2(G164), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n747), .A3(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n869), .A2(new_n759), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n760), .B1(new_n869), .B2(new_n874), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n875), .A2(new_n876), .A3(new_n624), .ZN(new_n877));
  INV_X1    g452(.A(new_n624), .ZN(new_n878));
  INV_X1    g453(.A(new_n760), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n867), .A2(new_n868), .A3(new_n746), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n747), .B1(new_n872), .B2(new_n873), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n869), .A2(new_n759), .A3(new_n874), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n711), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n877), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n624), .B1(new_n875), .B2(new_n876), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n878), .A3(new_n883), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n711), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n866), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(KEYINPUT104), .B(G37), .Z(new_n891));
  OAI21_X1  g466(.A(new_n885), .B1(new_n877), .B2(new_n884), .ZN(new_n892));
  INV_X1    g467(.A(new_n866), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n711), .A3(new_n888), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(new_n891), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(G395));
  XNOR2_X1  g473(.A(new_n616), .B(new_n850), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n605), .A2(G299), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n832), .A2(new_n795), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n605), .A2(KEYINPUT106), .A3(G299), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n906), .A3(new_n902), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n899), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n903), .A2(new_n904), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n899), .ZN(new_n913));
  XNOR2_X1  g488(.A(G290), .B(G288), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT108), .ZN(new_n916));
  XNOR2_X1  g491(.A(G305), .B(G166), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n914), .B(KEYINPUT108), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT109), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n922), .B(KEYINPUT42), .Z(new_n923));
  AND2_X1   g498(.A1(new_n913), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n913), .A2(new_n923), .ZN(new_n925));
  OAI21_X1  g500(.A(G868), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n843), .A2(new_n617), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(G295));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n927), .ZN(G331));
  NAND2_X1  g504(.A1(G286), .A2(G171), .ZN(new_n930));
  NAND2_X1  g505(.A1(G168), .A2(G301), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n851), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n850), .A2(new_n930), .A3(new_n931), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n851), .A3(KEYINPUT110), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n936), .A2(new_n905), .A3(new_n907), .A4(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n912), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n933), .A3(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n921), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n920), .A3(new_n940), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n936), .A2(new_n937), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n933), .A2(new_n935), .B1(new_n912), .B2(new_n906), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n900), .A2(new_n902), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT41), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n939), .A2(new_n948), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n891), .B(new_n944), .C1(new_n952), .C2(new_n920), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(new_n946), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT44), .B1(new_n947), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n946), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n942), .A2(KEYINPUT43), .A3(new_n943), .A4(new_n944), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n955), .B1(KEYINPUT44), .B2(new_n958), .ZN(G397));
  XOR2_X1   g534(.A(KEYINPUT111), .B(G1384), .Z(new_n960));
  NAND2_X1  g535(.A1(new_n871), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n468), .A2(new_n469), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n478), .ZN(new_n965));
  INV_X1    g540(.A(new_n475), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n622), .B2(G125), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT68), .B1(new_n967), .B2(new_n478), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n476), .A2(new_n471), .A3(G2105), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n965), .A2(G40), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n963), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT46), .Z(new_n974));
  INV_X1    g549(.A(new_n971), .ZN(new_n975));
  INV_X1    g550(.A(G2067), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n734), .B(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n977), .B2(new_n747), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n979), .B(KEYINPUT47), .Z(new_n980));
  INV_X1    g555(.A(new_n714), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n746), .B(new_n972), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n977), .A2(new_n711), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n735), .A2(new_n976), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n975), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT126), .ZN(new_n986));
  NOR2_X1   g561(.A1(G290), .A2(G1986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n971), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT48), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n977), .B(new_n982), .C1(new_n885), .C2(new_n714), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n885), .B2(new_n714), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n991), .B2(new_n975), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n980), .A2(new_n986), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n502), .B2(new_n505), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n970), .B1(new_n962), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT45), .B(new_n960), .C1(new_n502), .C2(new_n505), .ZN(new_n997));
  AOI21_X1  g572(.A(G1971), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n995), .A2(KEYINPUT50), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n968), .A2(new_n969), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n470), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1003), .B(new_n994), .C1(new_n502), .C2(new_n505), .ZN(new_n1004));
  AND4_X1   g579(.A1(new_n818), .A2(new_n999), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(G8), .B1(new_n998), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(G8), .B1(new_n521), .B2(new_n534), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT113), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n1010));
  NAND4_X1  g585(.A1(G303), .A2(new_n1010), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1006), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G305), .A2(G1981), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n589), .A2(new_n519), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT76), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n589), .A2(KEYINPUT76), .A3(new_n519), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1981), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(new_n582), .A4(new_n583), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT49), .B1(new_n1015), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n499), .A2(new_n501), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n503), .A2(new_n504), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(G2105), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n1002), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1015), .A2(new_n1022), .A3(KEYINPUT49), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1024), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n579), .A2(G1976), .A3(new_n580), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT114), .A4(G1976), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(G288), .B2(new_n688), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1030), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1036), .B(G8), .C1(new_n970), .C2(new_n995), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1035), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT52), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1014), .A2(new_n1032), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1009), .A2(new_n1012), .A3(new_n1011), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n999), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1046));
  OAI22_X1  g621(.A1(new_n998), .A2(KEYINPUT112), .B1(G2090), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n1048), .B(G1971), .C1(new_n996), .C2(new_n997), .ZN(new_n1049));
  OAI211_X1 g624(.A(G8), .B(new_n1045), .C1(new_n1047), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n995), .A2(new_n962), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT45), .B(new_n994), .C1(new_n502), .C2(new_n505), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1002), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n815), .ZN(new_n1055));
  INV_X1    g630(.A(G2084), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n999), .A2(new_n1002), .A3(new_n1056), .A4(new_n1004), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(G168), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1051), .B1(new_n1058), .B2(G8), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(G8), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1046), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1062), .A2(new_n1056), .B1(new_n1054), .B2(new_n815), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT51), .B1(new_n1063), .B2(G168), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1059), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1044), .B(new_n1050), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1052), .A2(new_n1002), .A3(new_n779), .A4(new_n997), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(G2078), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n996), .A2(new_n1053), .A3(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1070), .B(new_n1072), .C1(G1961), .C2(new_n1062), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1060), .A2(KEYINPUT51), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1051), .B1(new_n1077), .B2(G286), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1060), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1075), .B1(new_n1079), .B2(KEYINPUT62), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT124), .B1(new_n1067), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1074), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1015), .A2(new_n1022), .A3(KEYINPUT49), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(new_n1023), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1042), .B1(new_n1085), .B2(new_n1030), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1086), .A2(new_n1050), .A3(new_n1014), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1079), .A2(KEYINPUT62), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1082), .A2(new_n1083), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1081), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1348), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1046), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1029), .A2(KEYINPUT117), .A3(G160), .A4(G40), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n970), .B2(new_n995), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n976), .A3(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1092), .A2(new_n1096), .A3(new_n832), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n832), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT60), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n1100));
  INV_X1    g675(.A(G1956), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1046), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n1103));
  NAND2_X1  g678(.A1(G299), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n570), .A2(KEYINPUT57), .A3(new_n571), .A4(new_n573), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1052), .A2(new_n1002), .A3(new_n997), .A4(new_n1107), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1102), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1106), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1100), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1096), .A2(new_n1092), .A3(new_n605), .A4(new_n1112), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1099), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1110), .B1(new_n1109), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1102), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT120), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1116), .A2(new_n1117), .A3(KEYINPUT61), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1110), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1102), .A2(new_n1115), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1119), .A2(new_n1121), .A3(KEYINPUT61), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT121), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n996), .A2(new_n972), .A3(new_n997), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT58), .B(G1341), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n558), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1129));
  XNOR2_X1  g704(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1114), .A2(new_n1120), .A3(new_n1124), .A4(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1110), .B1(new_n1098), .B2(new_n1118), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(G1961), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1068), .A2(new_n1069), .B1(new_n1046), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(G40), .B1(new_n965), .B2(KEYINPUT122), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(KEYINPUT122), .B2(new_n965), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n997), .A2(new_n1071), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n476), .A2(G2105), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n963), .A2(new_n1137), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1135), .A2(G301), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT123), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1135), .A2(new_n1144), .A3(new_n1140), .A4(G301), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1142), .A2(new_n1143), .A3(new_n1074), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1073), .A2(G301), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1135), .A2(G171), .A3(new_n1140), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(KEYINPUT54), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1150), .A2(new_n1087), .A3(new_n1079), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1133), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1032), .A2(new_n688), .A3(new_n690), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n1022), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1050), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1154), .A2(new_n1030), .B1(new_n1155), .B2(new_n1086), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1063), .A2(new_n1025), .A3(G286), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1086), .A2(new_n1050), .A3(new_n1014), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT115), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT115), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1044), .A2(new_n1160), .A3(new_n1050), .A4(new_n1157), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(G8), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1045), .A2(KEYINPUT116), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1162), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1166), .A2(new_n1167), .A3(new_n1086), .A4(new_n1157), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1090), .A2(new_n1152), .A3(new_n1156), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(G290), .A2(G1986), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n991), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n971), .B1(new_n1172), .B2(new_n987), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1170), .A2(KEYINPUT125), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT125), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n993), .B1(new_n1174), .B2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g751(.A(new_n958), .ZN(new_n1178));
  INV_X1    g752(.A(G229), .ZN(new_n1179));
  INV_X1    g753(.A(G227), .ZN(new_n1180));
  NAND4_X1  g754(.A1(new_n1179), .A2(G319), .A3(new_n646), .A4(new_n1180), .ZN(new_n1181));
  XOR2_X1   g755(.A(new_n1181), .B(KEYINPUT127), .Z(new_n1182));
  AND3_X1   g756(.A1(new_n1178), .A2(new_n896), .A3(new_n1182), .ZN(G308));
  NAND3_X1  g757(.A1(new_n1178), .A2(new_n896), .A3(new_n1182), .ZN(G225));
endmodule


