

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738;

  NOR2_X1 U376 ( .A1(n605), .A2(n604), .ZN(n356) );
  XNOR2_X1 U377 ( .A(n421), .B(n705), .ZN(n430) );
  XNOR2_X1 U378 ( .A(G146), .B(G125), .ZN(n432) );
  XNOR2_X1 U379 ( .A(n379), .B(KEYINPUT18), .ZN(n376) );
  BUF_X1 U380 ( .A(G953), .Z(n355) );
  XNOR2_X1 U381 ( .A(KEYINPUT15), .B(G902), .ZN(n594) );
  NOR2_X2 U382 ( .A1(n618), .A2(n704), .ZN(n620) );
  NOR2_X2 U383 ( .A1(n626), .A2(n704), .ZN(n627) );
  XNOR2_X1 U384 ( .A(n356), .B(KEYINPUT91), .ZN(n520) );
  INV_X1 U385 ( .A(G902), .ZN(n441) );
  AND2_X1 U386 ( .A1(n574), .A2(n573), .ZN(n576) );
  INV_X1 U387 ( .A(n355), .ZN(n724) );
  XNOR2_X1 U388 ( .A(n547), .B(KEYINPUT83), .ZN(n635) );
  NOR2_X2 U389 ( .A1(n601), .A2(n704), .ZN(n603) );
  XNOR2_X2 U390 ( .A(n396), .B(n395), .ZN(n502) );
  OR2_X1 U391 ( .A1(n520), .A2(n522), .ZN(n362) );
  OR2_X1 U392 ( .A1(n568), .A2(n684), .ZN(n569) );
  XNOR2_X1 U393 ( .A(n427), .B(n426), .ZN(n669) );
  XNOR2_X1 U394 ( .A(n722), .B(n383), .ZN(n425) );
  XNOR2_X1 U395 ( .A(n390), .B(n476), .ZN(n722) );
  XNOR2_X1 U396 ( .A(n429), .B(n384), .ZN(n476) );
  INV_X2 U397 ( .A(G128), .ZN(n378) );
  BUF_X1 U398 ( .A(n621), .Z(n696) );
  NOR2_X1 U399 ( .A1(n669), .A2(n500), .ZN(n455) );
  BUF_X1 U400 ( .A(n622), .Z(n357) );
  XNOR2_X2 U401 ( .A(n502), .B(n397), .ZN(n673) );
  XNOR2_X2 U402 ( .A(KEYINPUT70), .B(G101), .ZN(n421) );
  XNOR2_X2 U403 ( .A(G110), .B(G104), .ZN(n705) );
  INV_X1 U404 ( .A(KEYINPUT67), .ZN(n516) );
  NOR2_X1 U405 ( .A1(n735), .A2(KEYINPUT44), .ZN(n521) );
  XNOR2_X1 U406 ( .A(n425), .B(n380), .ZN(n597) );
  XNOR2_X1 U407 ( .A(n382), .B(n381), .ZN(n380) );
  XNOR2_X1 U408 ( .A(n420), .B(n424), .ZN(n381) );
  XNOR2_X1 U409 ( .A(n422), .B(n359), .ZN(n382) );
  INV_X1 U410 ( .A(G134), .ZN(n384) );
  AND2_X1 U411 ( .A1(n564), .A2(n660), .ZN(n565) );
  XNOR2_X1 U412 ( .A(n411), .B(KEYINPUT25), .ZN(n412) );
  XNOR2_X1 U413 ( .A(n490), .B(n366), .ZN(n377) );
  NOR2_X1 U414 ( .A1(G237), .A2(G953), .ZN(n423) );
  INV_X1 U415 ( .A(KEYINPUT90), .ZN(n372) );
  XNOR2_X1 U416 ( .A(G131), .B(G116), .ZN(n418) );
  XOR2_X1 U417 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n419) );
  XNOR2_X1 U418 ( .A(G113), .B(G122), .ZN(n456) );
  XNOR2_X1 U419 ( .A(G113), .B(KEYINPUT3), .ZN(n417) );
  INV_X1 U420 ( .A(KEYINPUT48), .ZN(n575) );
  XNOR2_X1 U421 ( .A(n469), .B(n387), .ZN(n494) );
  XNOR2_X1 U422 ( .A(G116), .B(G122), .ZN(n436) );
  XNOR2_X1 U423 ( .A(n466), .B(n465), .ZN(n615) );
  INV_X1 U424 ( .A(n721), .ZN(n465) );
  XNOR2_X1 U425 ( .A(n462), .B(n461), .ZN(n466) );
  XNOR2_X1 U426 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U427 ( .A(G146), .ZN(n383) );
  INV_X1 U428 ( .A(KEYINPUT66), .ZN(n388) );
  NAND2_X1 U429 ( .A1(n363), .A2(n586), .ZN(n723) );
  AND2_X1 U430 ( .A1(n736), .A2(n585), .ZN(n586) );
  XOR2_X1 U431 ( .A(n576), .B(n575), .Z(n363) );
  INV_X1 U432 ( .A(n649), .ZN(n585) );
  XNOR2_X1 U433 ( .A(n480), .B(n479), .ZN(n497) );
  XNOR2_X1 U434 ( .A(n566), .B(KEYINPUT40), .ZN(n738) );
  XNOR2_X1 U435 ( .A(n483), .B(KEYINPUT87), .ZN(n484) );
  XNOR2_X1 U436 ( .A(n511), .B(KEYINPUT107), .ZN(n604) );
  XOR2_X1 U437 ( .A(n444), .B(n443), .Z(n358) );
  XOR2_X1 U438 ( .A(n419), .B(n418), .Z(n359) );
  XOR2_X1 U439 ( .A(KEYINPUT12), .B(G104), .Z(n360) );
  AND2_X1 U440 ( .A1(n377), .A2(n673), .ZN(n361) );
  AND2_X1 U441 ( .A1(n513), .A2(n551), .ZN(n364) );
  AND2_X1 U442 ( .A1(n673), .A2(n510), .ZN(n365) );
  XOR2_X1 U443 ( .A(KEYINPUT76), .B(KEYINPUT22), .Z(n366) );
  XOR2_X1 U444 ( .A(n523), .B(KEYINPUT65), .Z(n367) );
  XNOR2_X2 U445 ( .A(n368), .B(n358), .ZN(n537) );
  NAND2_X1 U446 ( .A1(n622), .A2(n594), .ZN(n368) );
  XNOR2_X1 U447 ( .A(n369), .B(n707), .ZN(n622) );
  XNOR2_X1 U448 ( .A(n374), .B(n435), .ZN(n369) );
  XNOR2_X1 U449 ( .A(n439), .B(n438), .ZN(n707) );
  XNOR2_X2 U450 ( .A(n370), .B(n367), .ZN(n710) );
  NAND2_X1 U451 ( .A1(n371), .A2(n362), .ZN(n370) );
  XNOR2_X1 U452 ( .A(n373), .B(n372), .ZN(n371) );
  NAND2_X1 U453 ( .A1(n518), .A2(n519), .ZN(n373) );
  XNOR2_X1 U454 ( .A(n375), .B(n430), .ZN(n374) );
  XNOR2_X1 U455 ( .A(n376), .B(n429), .ZN(n375) );
  XNOR2_X2 U456 ( .A(n378), .B(G143), .ZN(n429) );
  NAND2_X1 U457 ( .A1(n377), .A2(n365), .ZN(n511) );
  AND2_X1 U458 ( .A1(n377), .A2(n364), .ZN(n514) );
  NAND2_X1 U459 ( .A1(n428), .A2(G224), .ZN(n379) );
  BUF_X1 U460 ( .A(n488), .Z(n503) );
  XOR2_X1 U461 ( .A(n543), .B(KEYINPUT28), .Z(n385) );
  XOR2_X1 U462 ( .A(KEYINPUT41), .B(KEYINPUT109), .Z(n386) );
  XOR2_X1 U463 ( .A(n468), .B(n467), .Z(n387) );
  INV_X1 U464 ( .A(KEYINPUT47), .ZN(n548) );
  AND2_X1 U465 ( .A1(n562), .A2(n561), .ZN(n574) );
  INV_X1 U466 ( .A(KEYINPUT8), .ZN(n398) );
  XNOR2_X1 U467 ( .A(n399), .B(n398), .ZN(n474) );
  XNOR2_X1 U468 ( .A(n389), .B(n433), .ZN(n390) );
  XNOR2_X1 U469 ( .A(n567), .B(n386), .ZN(n684) );
  INV_X1 U470 ( .A(KEYINPUT63), .ZN(n602) );
  XOR2_X1 U471 ( .A(KEYINPUT73), .B(G137), .Z(n389) );
  XNOR2_X1 U472 ( .A(n388), .B(KEYINPUT4), .ZN(n433) );
  XOR2_X1 U473 ( .A(G131), .B(G140), .Z(n464) );
  XOR2_X1 U474 ( .A(G107), .B(n464), .Z(n392) );
  NAND2_X1 U475 ( .A1(G227), .A2(n724), .ZN(n391) );
  XNOR2_X1 U476 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U477 ( .A(n430), .B(n393), .ZN(n394) );
  XNOR2_X1 U478 ( .A(n425), .B(n394), .ZN(n697) );
  NAND2_X1 U479 ( .A1(n697), .A2(n441), .ZN(n396) );
  INV_X1 U480 ( .A(G469), .ZN(n395) );
  XNOR2_X1 U481 ( .A(KEYINPUT68), .B(KEYINPUT1), .ZN(n397) );
  INV_X1 U482 ( .A(G953), .ZN(n428) );
  NAND2_X1 U483 ( .A1(n428), .A2(G234), .ZN(n399) );
  NAND2_X1 U484 ( .A1(G221), .A2(n474), .ZN(n401) );
  XNOR2_X1 U485 ( .A(KEYINPUT10), .B(KEYINPUT72), .ZN(n400) );
  XNOR2_X1 U486 ( .A(n400), .B(n432), .ZN(n463) );
  XOR2_X1 U487 ( .A(n401), .B(n463), .Z(n409) );
  XOR2_X1 U488 ( .A(G140), .B(G110), .Z(n403) );
  XNOR2_X1 U489 ( .A(G128), .B(G119), .ZN(n402) );
  XNOR2_X1 U490 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U491 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n405) );
  XNOR2_X1 U492 ( .A(G137), .B(KEYINPUT94), .ZN(n404) );
  XNOR2_X1 U493 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U494 ( .A(n407), .B(n406), .Z(n408) );
  XNOR2_X1 U495 ( .A(n409), .B(n408), .ZN(n606) );
  NOR2_X1 U496 ( .A1(n606), .A2(G902), .ZN(n413) );
  NAND2_X1 U497 ( .A1(G234), .A2(n594), .ZN(n410) );
  XNOR2_X1 U498 ( .A(KEYINPUT20), .B(n410), .ZN(n414) );
  NAND2_X1 U499 ( .A1(G217), .A2(n414), .ZN(n411) );
  XNOR2_X2 U500 ( .A(n413), .B(n412), .ZN(n527) );
  AND2_X1 U501 ( .A1(n414), .A2(G221), .ZN(n415) );
  XNOR2_X1 U502 ( .A(n415), .B(KEYINPUT21), .ZN(n487) );
  NAND2_X1 U503 ( .A1(n527), .A2(n487), .ZN(n674) );
  NOR2_X1 U504 ( .A1(n673), .A2(n674), .ZN(n416) );
  INV_X1 U505 ( .A(n416), .ZN(n499) );
  XNOR2_X1 U506 ( .A(n417), .B(G119), .ZN(n437) );
  INV_X1 U507 ( .A(n437), .ZN(n420) );
  XOR2_X1 U508 ( .A(KEYINPUT95), .B(n421), .Z(n422) );
  XNOR2_X1 U509 ( .A(n423), .B(KEYINPUT80), .ZN(n458) );
  NAND2_X1 U510 ( .A1(G210), .A2(n458), .ZN(n424) );
  NAND2_X1 U511 ( .A1(n597), .A2(n441), .ZN(n529) );
  INV_X1 U512 ( .A(G472), .ZN(n528) );
  XNOR2_X2 U513 ( .A(n529), .B(n528), .ZN(n498) );
  XOR2_X1 U514 ( .A(KEYINPUT6), .B(n498), .Z(n551) );
  NOR2_X1 U515 ( .A1(n499), .A2(n551), .ZN(n427) );
  XNOR2_X1 U516 ( .A(KEYINPUT92), .B(KEYINPUT33), .ZN(n426) );
  XNOR2_X1 U517 ( .A(KEYINPUT81), .B(KEYINPUT17), .ZN(n431) );
  XNOR2_X1 U518 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U519 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U520 ( .A(n436), .B(G107), .ZN(n473) );
  XNOR2_X1 U521 ( .A(n437), .B(n473), .ZN(n439) );
  XOR2_X1 U522 ( .A(KEYINPUT77), .B(KEYINPUT16), .Z(n438) );
  INV_X1 U523 ( .A(G237), .ZN(n440) );
  NAND2_X1 U524 ( .A1(n441), .A2(n440), .ZN(n445) );
  NAND2_X1 U525 ( .A1(n445), .A2(G210), .ZN(n444) );
  INV_X1 U526 ( .A(KEYINPUT84), .ZN(n442) );
  XNOR2_X1 U527 ( .A(n442), .B(KEYINPUT93), .ZN(n443) );
  NAND2_X1 U528 ( .A1(n445), .A2(G214), .ZN(n659) );
  NAND2_X1 U529 ( .A1(n537), .A2(n659), .ZN(n447) );
  INV_X1 U530 ( .A(KEYINPUT19), .ZN(n446) );
  XNOR2_X1 U531 ( .A(n447), .B(n446), .ZN(n545) );
  NAND2_X1 U532 ( .A1(G234), .A2(G237), .ZN(n448) );
  XNOR2_X1 U533 ( .A(n448), .B(KEYINPUT14), .ZN(n690) );
  NOR2_X1 U534 ( .A1(G902), .A2(n724), .ZN(n450) );
  NOR2_X1 U535 ( .A1(n355), .A2(G952), .ZN(n449) );
  NOR2_X1 U536 ( .A1(n450), .A2(n449), .ZN(n451) );
  NAND2_X1 U537 ( .A1(n690), .A2(n451), .ZN(n524) );
  AND2_X1 U538 ( .A1(n355), .A2(G898), .ZN(n452) );
  OR2_X1 U539 ( .A1(n524), .A2(n452), .ZN(n453) );
  NOR2_X2 U540 ( .A1(n545), .A2(n453), .ZN(n454) );
  XNOR2_X1 U541 ( .A(n454), .B(KEYINPUT0), .ZN(n488) );
  INV_X1 U542 ( .A(n503), .ZN(n500) );
  XNOR2_X1 U543 ( .A(KEYINPUT34), .B(n455), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n360), .B(n456), .ZN(n457) );
  XOR2_X1 U545 ( .A(n457), .B(KEYINPUT11), .Z(n462) );
  NAND2_X1 U546 ( .A1(n458), .A2(G214), .ZN(n460) );
  XNOR2_X1 U547 ( .A(G143), .B(KEYINPUT97), .ZN(n459) );
  XNOR2_X1 U548 ( .A(n464), .B(n463), .ZN(n721) );
  NOR2_X1 U549 ( .A1(n615), .A2(G902), .ZN(n469) );
  XOR2_X1 U550 ( .A(KEYINPUT99), .B(KEYINPUT13), .Z(n468) );
  XNOR2_X1 U551 ( .A(KEYINPUT98), .B(G475), .ZN(n467) );
  XNOR2_X1 U552 ( .A(KEYINPUT102), .B(G478), .ZN(n480) );
  XOR2_X1 U553 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n471) );
  XNOR2_X1 U554 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n470) );
  XNOR2_X1 U555 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U556 ( .A(n473), .B(n472), .Z(n478) );
  NAND2_X1 U557 ( .A1(G217), .A2(n474), .ZN(n475) );
  XNOR2_X1 U558 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U559 ( .A(n478), .B(n477), .Z(n610) );
  NOR2_X1 U560 ( .A1(G902), .A2(n610), .ZN(n479) );
  NOR2_X1 U561 ( .A1(n494), .A2(n497), .ZN(n536) );
  XNOR2_X1 U562 ( .A(n536), .B(KEYINPUT82), .ZN(n481) );
  NAND2_X1 U563 ( .A1(n482), .A2(n481), .ZN(n485) );
  INV_X1 U564 ( .A(KEYINPUT35), .ZN(n483) );
  XNOR2_X2 U565 ( .A(n485), .B(n484), .ZN(n735) );
  NAND2_X1 U566 ( .A1(n735), .A2(KEYINPUT44), .ZN(n509) );
  AND2_X1 U567 ( .A1(n494), .A2(n497), .ZN(n486) );
  XNOR2_X1 U568 ( .A(n486), .B(KEYINPUT105), .ZN(n662) );
  INV_X1 U569 ( .A(n487), .ZN(n671) );
  NOR2_X1 U570 ( .A1(n662), .A2(n671), .ZN(n489) );
  NAND2_X1 U571 ( .A1(n489), .A2(n488), .ZN(n490) );
  INV_X1 U572 ( .A(n673), .ZN(n558) );
  NAND2_X1 U573 ( .A1(n361), .A2(n551), .ZN(n491) );
  XOR2_X1 U574 ( .A(KEYINPUT89), .B(n491), .Z(n493) );
  INV_X1 U575 ( .A(KEYINPUT106), .ZN(n492) );
  XNOR2_X1 U576 ( .A(n527), .B(n492), .ZN(n670) );
  NOR2_X1 U577 ( .A1(n493), .A2(n670), .ZN(n628) );
  INV_X1 U578 ( .A(n494), .ZN(n496) );
  NAND2_X1 U579 ( .A1(n497), .A2(n496), .ZN(n495) );
  XNOR2_X1 U580 ( .A(KEYINPUT103), .B(n495), .ZN(n643) );
  NOR2_X1 U581 ( .A1(n497), .A2(n496), .ZN(n645) );
  INV_X1 U582 ( .A(n645), .ZN(n636) );
  XOR2_X1 U583 ( .A(KEYINPUT104), .B(n636), .Z(n584) );
  NOR2_X1 U584 ( .A1(n643), .A2(n584), .ZN(n664) );
  OR2_X1 U585 ( .A1(n498), .A2(n499), .ZN(n682) );
  NOR2_X1 U586 ( .A1(n500), .A2(n682), .ZN(n501) );
  XOR2_X1 U587 ( .A(KEYINPUT31), .B(n501), .Z(n646) );
  INV_X1 U588 ( .A(n502), .ZN(n534) );
  INV_X1 U589 ( .A(n534), .ZN(n544) );
  INV_X1 U590 ( .A(n498), .ZN(n677) );
  NOR2_X1 U591 ( .A1(n677), .A2(n674), .ZN(n504) );
  NAND2_X1 U592 ( .A1(n504), .A2(n503), .ZN(n505) );
  NOR2_X1 U593 ( .A1(n544), .A2(n505), .ZN(n630) );
  NOR2_X1 U594 ( .A1(n646), .A2(n630), .ZN(n506) );
  NOR2_X1 U595 ( .A1(n664), .A2(n506), .ZN(n507) );
  NOR2_X1 U596 ( .A1(n628), .A2(n507), .ZN(n508) );
  AND2_X1 U597 ( .A1(n509), .A2(n508), .ZN(n519) );
  NOR2_X1 U598 ( .A1(n677), .A2(n527), .ZN(n510) );
  INV_X1 U599 ( .A(n670), .ZN(n512) );
  NOR2_X1 U600 ( .A1(n673), .A2(n512), .ZN(n513) );
  XNOR2_X1 U601 ( .A(n514), .B(KEYINPUT32), .ZN(n605) );
  NAND2_X1 U602 ( .A1(n520), .A2(KEYINPUT44), .ZN(n517) );
  XNOR2_X1 U603 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U604 ( .A(n521), .B(KEYINPUT71), .ZN(n522) );
  XNOR2_X1 U605 ( .A(KEYINPUT86), .B(KEYINPUT45), .ZN(n523) );
  NOR2_X1 U606 ( .A1(n671), .A2(n524), .ZN(n526) );
  NAND2_X1 U607 ( .A1(n355), .A2(G900), .ZN(n525) );
  NAND2_X1 U608 ( .A1(n526), .A2(n525), .ZN(n539) );
  INV_X1 U609 ( .A(n527), .ZN(n540) );
  OR2_X1 U610 ( .A1(n539), .A2(n540), .ZN(n533) );
  XOR2_X1 U611 ( .A(n529), .B(n528), .Z(n530) );
  NAND2_X1 U612 ( .A1(n530), .A2(n659), .ZN(n531) );
  XNOR2_X1 U613 ( .A(n531), .B(KEYINPUT30), .ZN(n532) );
  NOR2_X1 U614 ( .A1(n533), .A2(n532), .ZN(n535) );
  AND2_X1 U615 ( .A1(n535), .A2(n534), .ZN(n564) );
  NAND2_X1 U616 ( .A1(n564), .A2(n536), .ZN(n538) );
  BUF_X1 U617 ( .A(n537), .Z(n555) );
  INV_X1 U618 ( .A(n555), .ZN(n579) );
  NOR2_X1 U619 ( .A1(n538), .A2(n579), .ZN(n639) );
  XNOR2_X1 U620 ( .A(n539), .B(KEYINPUT75), .ZN(n541) );
  NAND2_X1 U621 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U622 ( .A(n542), .B(KEYINPUT74), .ZN(n552) );
  NOR2_X1 U623 ( .A1(n552), .A2(n498), .ZN(n543) );
  OR2_X2 U624 ( .A1(n385), .A2(n544), .ZN(n568) );
  BUF_X1 U625 ( .A(n545), .Z(n546) );
  NOR2_X2 U626 ( .A1(n568), .A2(n546), .ZN(n547) );
  NOR2_X1 U627 ( .A1(n664), .A2(n635), .ZN(n549) );
  XNOR2_X1 U628 ( .A(n549), .B(n548), .ZN(n550) );
  NOR2_X1 U629 ( .A1(n639), .A2(n550), .ZN(n562) );
  INV_X1 U630 ( .A(n643), .ZN(n641) );
  NOR2_X1 U631 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U632 ( .A1(n553), .A2(n659), .ZN(n554) );
  NOR2_X1 U633 ( .A1(n641), .A2(n554), .ZN(n577) );
  NAND2_X1 U634 ( .A1(n577), .A2(n555), .ZN(n557) );
  XOR2_X1 U635 ( .A(KEYINPUT110), .B(KEYINPUT36), .Z(n556) );
  XNOR2_X1 U636 ( .A(n557), .B(n556), .ZN(n559) );
  NAND2_X1 U637 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U638 ( .A(n560), .B(KEYINPUT111), .ZN(n732) );
  INV_X1 U639 ( .A(n732), .ZN(n561) );
  XNOR2_X1 U640 ( .A(KEYINPUT78), .B(KEYINPUT38), .ZN(n563) );
  XNOR2_X1 U641 ( .A(n579), .B(n563), .ZN(n660) );
  XOR2_X1 U642 ( .A(n565), .B(KEYINPUT39), .Z(n583) );
  NAND2_X1 U643 ( .A1(n583), .A2(n643), .ZN(n566) );
  NAND2_X1 U644 ( .A1(n660), .A2(n659), .ZN(n663) );
  NOR2_X1 U645 ( .A1(n662), .A2(n663), .ZN(n567) );
  XNOR2_X1 U646 ( .A(n569), .B(KEYINPUT42), .ZN(n737) );
  NAND2_X1 U647 ( .A1(n738), .A2(n737), .ZN(n572) );
  XOR2_X1 U648 ( .A(KEYINPUT46), .B(KEYINPUT88), .Z(n570) );
  XNOR2_X1 U649 ( .A(KEYINPUT64), .B(n570), .ZN(n571) );
  XNOR2_X1 U650 ( .A(n572), .B(n571), .ZN(n573) );
  NAND2_X1 U651 ( .A1(n577), .A2(n673), .ZN(n578) );
  XNOR2_X1 U652 ( .A(KEYINPUT43), .B(n578), .ZN(n580) );
  AND2_X1 U653 ( .A1(n580), .A2(n579), .ZN(n582) );
  INV_X1 U654 ( .A(KEYINPUT108), .ZN(n581) );
  XNOR2_X1 U655 ( .A(n582), .B(n581), .ZN(n736) );
  AND2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n649) );
  INV_X1 U657 ( .A(n723), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n710), .A2(n589), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n587), .A2(KEYINPUT2), .ZN(n652) );
  NOR2_X1 U660 ( .A1(KEYINPUT2), .A2(KEYINPUT79), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n723), .A2(KEYINPUT79), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n592), .A2(n710), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n652), .A2(n593), .ZN(n596) );
  INV_X1 U666 ( .A(n594), .ZN(n595) );
  AND2_X2 U667 ( .A1(n596), .A2(n595), .ZN(n621) );
  NAND2_X1 U668 ( .A1(n621), .A2(G472), .ZN(n599) );
  XOR2_X1 U669 ( .A(n597), .B(KEYINPUT62), .Z(n598) );
  XNOR2_X1 U670 ( .A(n599), .B(n598), .ZN(n601) );
  INV_X1 U671 ( .A(G952), .ZN(n600) );
  AND2_X1 U672 ( .A1(n600), .A2(n355), .ZN(n704) );
  XNOR2_X1 U673 ( .A(n603), .B(n602), .ZN(G57) );
  XOR2_X1 U674 ( .A(n604), .B(G110), .Z(G12) );
  XOR2_X1 U675 ( .A(n605), .B(G119), .Z(G21) );
  NAND2_X1 U676 ( .A1(n696), .A2(G217), .ZN(n608) );
  XOR2_X1 U677 ( .A(KEYINPUT123), .B(n606), .Z(n607) );
  XNOR2_X1 U678 ( .A(n608), .B(n607), .ZN(n609) );
  NOR2_X1 U679 ( .A1(n609), .A2(n704), .ZN(G66) );
  NAND2_X1 U680 ( .A1(n696), .A2(G478), .ZN(n612) );
  XNOR2_X1 U681 ( .A(n610), .B(KEYINPUT122), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n612), .B(n611), .ZN(n613) );
  NOR2_X1 U683 ( .A1(n613), .A2(n704), .ZN(G63) );
  NAND2_X1 U684 ( .A1(n621), .A2(G475), .ZN(n617) );
  XNOR2_X1 U685 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n618) );
  XOR2_X1 U688 ( .A(KEYINPUT69), .B(KEYINPUT60), .Z(n619) );
  XNOR2_X1 U689 ( .A(n620), .B(n619), .ZN(G60) );
  NAND2_X1 U690 ( .A1(n621), .A2(G210), .ZN(n625) );
  XNOR2_X1 U691 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n357), .B(n623), .ZN(n624) );
  XNOR2_X1 U693 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U694 ( .A(n627), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U695 ( .A(G101), .B(n628), .Z(G3) );
  NAND2_X1 U696 ( .A1(n630), .A2(n643), .ZN(n629) );
  XNOR2_X1 U697 ( .A(n629), .B(G104), .ZN(G6) );
  XNOR2_X1 U698 ( .A(G107), .B(KEYINPUT27), .ZN(n634) );
  XOR2_X1 U699 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n632) );
  NAND2_X1 U700 ( .A1(n630), .A2(n645), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(G9) );
  NOR2_X1 U703 ( .A1(n636), .A2(n635), .ZN(n638) );
  XNOR2_X1 U704 ( .A(G128), .B(KEYINPUT29), .ZN(n637) );
  XNOR2_X1 U705 ( .A(n638), .B(n637), .ZN(G30) );
  XNOR2_X1 U706 ( .A(n639), .B(G143), .ZN(n640) );
  XNOR2_X1 U707 ( .A(n640), .B(KEYINPUT113), .ZN(G45) );
  NOR2_X1 U708 ( .A1(n641), .A2(n635), .ZN(n642) );
  XOR2_X1 U709 ( .A(G146), .B(n642), .Z(G48) );
  NAND2_X1 U710 ( .A1(n646), .A2(n643), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n644), .B(G113), .ZN(G15) );
  NAND2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U713 ( .A(n647), .B(KEYINPUT114), .ZN(n648) );
  XNOR2_X1 U714 ( .A(G116), .B(n648), .ZN(G18) );
  XOR2_X1 U715 ( .A(G134), .B(n649), .Z(G36) );
  NOR2_X1 U716 ( .A1(n669), .A2(n684), .ZN(n650) );
  NOR2_X1 U717 ( .A1(n355), .A2(n650), .ZN(n658) );
  INV_X1 U718 ( .A(KEYINPUT2), .ZN(n653) );
  NAND2_X1 U719 ( .A1(n723), .A2(n653), .ZN(n651) );
  XOR2_X1 U720 ( .A(KEYINPUT85), .B(n651), .Z(n656) );
  NAND2_X1 U721 ( .A1(n710), .A2(n653), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n652), .A2(n654), .ZN(n655) );
  NAND2_X1 U723 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U724 ( .A1(n658), .A2(n657), .ZN(n694) );
  NOR2_X1 U725 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U726 ( .A1(n662), .A2(n661), .ZN(n667) );
  NOR2_X1 U727 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U728 ( .A(KEYINPUT117), .B(n665), .Z(n666) );
  NOR2_X1 U729 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U730 ( .A1(n669), .A2(n668), .ZN(n687) );
  NAND2_X1 U731 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U732 ( .A(KEYINPUT49), .B(n672), .Z(n680) );
  XOR2_X1 U733 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n676) );
  NAND2_X1 U734 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U735 ( .A(n676), .B(n675), .ZN(n678) );
  NOR2_X1 U736 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U737 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U738 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U739 ( .A(KEYINPUT51), .B(n683), .ZN(n685) );
  NOR2_X1 U740 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U741 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U742 ( .A(n688), .B(KEYINPUT52), .ZN(n689) );
  XNOR2_X1 U743 ( .A(n689), .B(KEYINPUT118), .ZN(n692) );
  NAND2_X1 U744 ( .A1(n690), .A2(G952), .ZN(n691) );
  NOR2_X1 U745 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U746 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U747 ( .A(KEYINPUT53), .B(n695), .ZN(G75) );
  NAND2_X1 U748 ( .A1(n696), .A2(G469), .ZN(n702) );
  XOR2_X1 U749 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n699) );
  XNOR2_X1 U750 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n698) );
  XNOR2_X1 U751 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U752 ( .A(n697), .B(n700), .ZN(n701) );
  XNOR2_X1 U753 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U754 ( .A1(n704), .A2(n703), .ZN(G54) );
  XNOR2_X1 U755 ( .A(n705), .B(G101), .ZN(n706) );
  XNOR2_X1 U756 ( .A(n707), .B(n706), .ZN(n709) );
  NOR2_X1 U757 ( .A1(G898), .A2(n724), .ZN(n708) );
  NOR2_X1 U758 ( .A1(n709), .A2(n708), .ZN(n720) );
  INV_X1 U759 ( .A(n710), .ZN(n711) );
  NOR2_X1 U760 ( .A1(n711), .A2(n355), .ZN(n717) );
  NAND2_X1 U761 ( .A1(G224), .A2(n355), .ZN(n712) );
  XNOR2_X1 U762 ( .A(n712), .B(KEYINPUT61), .ZN(n713) );
  XNOR2_X1 U763 ( .A(KEYINPUT124), .B(n713), .ZN(n714) );
  NAND2_X1 U764 ( .A1(n714), .A2(G898), .ZN(n715) );
  XNOR2_X1 U765 ( .A(n715), .B(KEYINPUT125), .ZN(n716) );
  NOR2_X1 U766 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U767 ( .A(n718), .B(KEYINPUT126), .Z(n719) );
  XNOR2_X1 U768 ( .A(n720), .B(n719), .ZN(G69) );
  XNOR2_X1 U769 ( .A(n722), .B(n721), .ZN(n726) );
  XOR2_X1 U770 ( .A(n723), .B(n726), .Z(n725) );
  NAND2_X1 U771 ( .A1(n725), .A2(n724), .ZN(n731) );
  XNOR2_X1 U772 ( .A(n726), .B(G227), .ZN(n727) );
  XNOR2_X1 U773 ( .A(n727), .B(KEYINPUT127), .ZN(n728) );
  NAND2_X1 U774 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U775 ( .A1(n355), .A2(n729), .ZN(n730) );
  NAND2_X1 U776 ( .A1(n731), .A2(n730), .ZN(G72) );
  XOR2_X1 U777 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n734) );
  XNOR2_X1 U778 ( .A(G125), .B(n732), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n734), .B(n733), .ZN(G27) );
  XOR2_X1 U780 ( .A(G122), .B(n735), .Z(G24) );
  XNOR2_X1 U781 ( .A(G140), .B(n736), .ZN(G42) );
  XNOR2_X1 U782 ( .A(G137), .B(n737), .ZN(G39) );
  XNOR2_X1 U783 ( .A(G131), .B(n738), .ZN(G33) );
endmodule

