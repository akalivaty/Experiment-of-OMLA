//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0006(.A(G250), .ZN(new_n207));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n207), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n215), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n214), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n232), .A2(G1), .A3(G13), .ZN(new_n233));
  INV_X1    g0033(.A(G68), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n202), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g0037(.A(new_n237), .B1(new_n216), .B2(KEYINPUT0), .ZN(new_n238));
  NAND3_X1  g0038(.A1(new_n217), .A2(new_n228), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g0039(.A(new_n239), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n224), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT16), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT7), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT65), .B(G20), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR4_X1   g0062(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT7), .A4(G20), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n262), .A2(new_n263), .A3(new_n234), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G58), .A2(G68), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT69), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G58), .A3(G68), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(new_n268), .A3(new_n235), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(G159), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n209), .A2(new_n272), .A3(KEYINPUT66), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT66), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(G20), .B2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n270), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n256), .B1(new_n264), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n260), .A2(new_n261), .A3(new_n257), .ZN(new_n283));
  OR2_X1    g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n209), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT7), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n283), .A2(new_n287), .A3(G68), .ZN(new_n288));
  AOI22_X1  g0088(.A1(G20), .A2(new_n269), .B1(new_n276), .B2(G159), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(KEYINPUT16), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n279), .A2(new_n282), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n209), .A2(G1), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n294), .A2(KEYINPUT70), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(new_n281), .A3(new_n280), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n294), .B2(KEYINPUT70), .ZN(new_n298));
  INV_X1    g0098(.A(new_n296), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n295), .A2(new_n298), .B1(new_n299), .B2(new_n292), .ZN(new_n300));
  INV_X1    g0100(.A(G41), .ZN(new_n301));
  OAI211_X1 g0101(.A(G1), .B(G13), .C1(new_n272), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G45), .ZN(new_n303));
  AOI21_X1  g0103(.A(G1), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(G274), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n307), .B2(new_n224), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(G226), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G87), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G1698), .ZN(new_n313));
  OAI211_X1 g0113(.A(G223), .B(new_n313), .C1(new_n258), .C2(new_n259), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT71), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT3), .B(G33), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n317), .A2(KEYINPUT71), .A3(G223), .A4(new_n313), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n312), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n309), .B(G190), .C1(new_n319), .C2(new_n302), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n316), .A2(new_n318), .ZN(new_n321));
  INV_X1    g0121(.A(new_n312), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n302), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(G200), .B1(new_n323), .B2(new_n308), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n291), .A2(new_n300), .A3(new_n320), .A4(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT17), .ZN(new_n326));
  OAI21_X1  g0126(.A(G169), .B1(new_n323), .B2(new_n308), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n309), .B(G179), .C1(new_n319), .C2(new_n302), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n290), .A2(new_n282), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n260), .A2(new_n257), .A3(new_n209), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n232), .A2(new_n317), .ZN(new_n332));
  OAI211_X1 g0132(.A(G68), .B(new_n331), .C1(new_n332), .C2(new_n257), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT16), .B1(new_n333), .B2(new_n289), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n300), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT18), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n329), .A2(new_n335), .A3(KEYINPUT18), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n326), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n317), .A2(G223), .A3(G1698), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n317), .A2(new_n313), .ZN(new_n344));
  INV_X1    g0144(.A(G222), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n343), .B1(new_n219), .B2(new_n317), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n281), .B1(G33), .B2(G41), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n305), .ZN(new_n349));
  INV_X1    g0149(.A(new_n307), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(G226), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n261), .A2(G33), .ZN(new_n356));
  INV_X1    g0156(.A(G150), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n355), .B1(new_n356), .B2(new_n292), .C1(new_n357), .C2(new_n277), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n282), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n297), .A2(new_n201), .A3(new_n293), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n201), .B2(new_n299), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n354), .B(new_n362), .C1(G179), .C2(new_n352), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n362), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(KEYINPUT9), .B1(new_n352), .B2(G200), .ZN(new_n366));
  INV_X1    g0166(.A(new_n352), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT9), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n367), .A2(G190), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT10), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT10), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n366), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n364), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n317), .A2(G232), .A3(G1698), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n317), .A2(G226), .A3(new_n313), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n375), .B(new_n376), .C1(new_n272), .C2(new_n225), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n347), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT13), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n349), .B1(G238), .B2(new_n350), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n379), .B1(new_n378), .B2(new_n380), .ZN(new_n382));
  OAI21_X1  g0182(.A(G200), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n378), .A2(new_n380), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT13), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n378), .A2(new_n380), .A3(new_n379), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(G190), .A3(new_n386), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n356), .A2(new_n219), .B1(new_n209), .B2(G68), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n277), .A2(new_n201), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n282), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT11), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n297), .A2(new_n234), .A3(new_n293), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT12), .B1(new_n296), .B2(G68), .ZN(new_n394));
  OR3_X1    g0194(.A1(new_n296), .A2(KEYINPUT12), .A3(G68), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n390), .B2(new_n391), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n383), .A2(new_n387), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(G169), .B1(new_n381), .B2(new_n382), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT14), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n385), .A2(new_n386), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT14), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(G169), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n385), .A2(G179), .A3(new_n386), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n398), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n400), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n277), .A2(new_n292), .B1(new_n219), .B2(new_n261), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT15), .B(G87), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n356), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n282), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(G77), .B1(new_n209), .B2(G1), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n297), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n219), .B2(new_n299), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n317), .A2(G232), .A3(new_n313), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n317), .A2(G238), .A3(G1698), .ZN(new_n419));
  AND2_X1   g0219(.A1(KEYINPUT68), .A2(G107), .ZN(new_n420));
  NOR2_X1   g0220(.A1(KEYINPUT68), .A2(G107), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n418), .B(new_n419), .C1(new_n317), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n347), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n305), .B1(new_n307), .B2(new_n220), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT67), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT67), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n305), .B(new_n427), .C1(new_n307), .C2(new_n220), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n417), .B1(new_n429), .B2(G190), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G200), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n353), .ZN(new_n434));
  INV_X1    g0234(.A(G179), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n424), .A2(new_n435), .A3(new_n426), .A4(new_n428), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n436), .A3(new_n417), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n342), .A2(new_n374), .A3(new_n409), .A4(new_n438), .ZN(new_n439));
  OR2_X1    g0239(.A1(G238), .A2(G1698), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n220), .A2(G1698), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n440), .B(new_n441), .C1(new_n258), .C2(new_n259), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G116), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n347), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT73), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n208), .A2(G45), .A3(G274), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n347), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n303), .A2(G1), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n302), .A2(KEYINPUT73), .A3(G274), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(G250), .B1(new_n303), .B2(G1), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n347), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n445), .A2(new_n451), .A3(new_n435), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT74), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n229), .A2(new_n231), .A3(G33), .A4(G97), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT19), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n229), .A2(new_n231), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n221), .ZN(new_n463));
  NOR2_X1   g0263(.A1(G87), .A2(G97), .ZN(new_n464));
  NAND2_X1  g0264(.A1(KEYINPUT68), .A2(G107), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n261), .A2(new_n317), .A3(G68), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n459), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n282), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n411), .A2(new_n299), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n297), .B1(new_n208), .B2(G33), .ZN(new_n472));
  INV_X1    g0272(.A(new_n411), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n470), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n445), .A2(new_n451), .A3(new_n454), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n353), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n453), .B1(new_n444), .B2(new_n347), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT74), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(new_n435), .A4(new_n451), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n456), .A2(new_n475), .A3(new_n477), .A4(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT75), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n476), .A2(G200), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n469), .A2(new_n282), .B1(new_n299), .B2(new_n411), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n472), .A2(G87), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n478), .A2(G190), .A3(new_n451), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n483), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n481), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT6), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n490), .A2(G97), .A3(G107), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n225), .A2(KEYINPUT6), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n221), .A2(KEYINPUT72), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n221), .A2(KEYINPUT72), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n491), .A2(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT72), .B(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n225), .A2(new_n221), .A3(KEYINPUT6), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n490), .A2(G97), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n499), .A3(new_n232), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n276), .A2(G77), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n262), .A2(new_n263), .A3(new_n422), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n282), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n296), .A2(G97), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n282), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n507), .B(new_n296), .C1(G1), .C2(new_n272), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n508), .B2(new_n225), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(G1698), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(G244), .C1(new_n259), .C2(new_n258), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n220), .B1(new_n284), .B2(new_n285), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n515), .C1(new_n516), .C2(KEYINPUT4), .ZN(new_n517));
  OAI21_X1  g0317(.A(G250), .B1(new_n258), .B2(new_n259), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n313), .B1(new_n518), .B2(KEYINPUT4), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n347), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g0320(.A(KEYINPUT5), .B(G41), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n347), .B1(new_n449), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n347), .A2(new_n447), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n522), .A2(G257), .B1(new_n523), .B2(new_n521), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n353), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(new_n435), .A3(new_n524), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n511), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n525), .A2(G200), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n463), .A2(new_n465), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n331), .B(new_n530), .C1(new_n332), .C2(new_n257), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(new_n501), .A3(new_n500), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n509), .B1(new_n532), .B2(new_n282), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n520), .A2(G190), .A3(new_n524), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n529), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n482), .B1(new_n481), .B2(new_n487), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n489), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT21), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n317), .A2(G264), .A3(G1698), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n317), .A2(G257), .A3(new_n313), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n260), .A2(G303), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n543), .A2(new_n347), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n522), .A2(G270), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n523), .A2(new_n521), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(G169), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n296), .A2(G116), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G116), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n508), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n280), .A2(new_n281), .B1(G20), .B2(new_n551), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n515), .B1(new_n225), .B2(G33), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n232), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT20), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n552), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n539), .B1(new_n548), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n557), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n549), .B1(new_n472), .B2(G116), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n543), .A2(new_n347), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n546), .A3(new_n545), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n563), .A2(KEYINPUT21), .A3(G169), .A4(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n544), .A2(new_n547), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(new_n563), .A3(G179), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n560), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(G190), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n559), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n565), .A2(G200), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(KEYINPUT76), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n563), .B1(new_n567), .B2(G190), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT76), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n572), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n569), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  XOR2_X1   g0378(.A(KEYINPUT78), .B(KEYINPUT25), .Z(new_n579));
  NOR2_X1   g0379(.A1(new_n296), .A2(G107), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n579), .B1(KEYINPUT79), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT79), .B1(new_n299), .B2(new_n221), .ZN(new_n582));
  XOR2_X1   g0382(.A(new_n581), .B(new_n582), .Z(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(G107), .B2(new_n472), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT77), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT22), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n229), .B(new_n231), .C1(new_n258), .C2(new_n259), .ZN(new_n587));
  INV_X1    g0387(.A(G87), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n261), .A2(new_n317), .A3(KEYINPUT22), .A4(G87), .ZN(new_n590));
  OAI21_X1  g0390(.A(KEYINPUT23), .B1(new_n530), .B2(new_n209), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n443), .A2(G20), .ZN(new_n592));
  NOR2_X1   g0392(.A1(KEYINPUT23), .A2(G107), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n592), .B1(new_n232), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n589), .A2(new_n590), .A3(new_n591), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT24), .ZN(new_n596));
  INV_X1    g0396(.A(new_n593), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n261), .A2(new_n597), .B1(G20), .B2(new_n443), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT23), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n422), .B2(G20), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT24), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(new_n590), .A4(new_n589), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n596), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n585), .B1(new_n604), .B2(new_n282), .ZN(new_n605));
  AOI211_X1 g0405(.A(KEYINPUT77), .B(new_n507), .C1(new_n596), .C2(new_n603), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n584), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n317), .A2(G257), .A3(G1698), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G33), .A2(G294), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n608), .B(new_n609), .C1(new_n344), .C2(new_n207), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n347), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n522), .A2(G264), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n546), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(G179), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n353), .B2(new_n613), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G200), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n611), .A2(new_n570), .A3(new_n546), .A4(new_n612), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n584), .B(new_n620), .C1(new_n605), .C2(new_n606), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n538), .A2(new_n578), .A3(new_n616), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n439), .A2(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n439), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n528), .A2(new_n535), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n475), .A2(new_n477), .A3(new_n455), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n487), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n621), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT80), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n569), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n560), .A2(new_n566), .A3(KEYINPUT80), .A4(new_n568), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n629), .B1(new_n616), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n626), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n627), .A2(new_n528), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n489), .A2(new_n537), .A3(new_n528), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(new_n637), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n624), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT81), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n329), .A2(new_n335), .A3(KEYINPUT18), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT18), .B1(new_n329), .B2(new_n335), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n338), .A2(KEYINPUT81), .A3(new_n339), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n437), .B(KEYINPUT82), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n408), .B2(new_n407), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n326), .A2(new_n399), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n646), .B(new_n647), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n371), .A2(new_n373), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n364), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n642), .A2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(KEYINPUT84), .ZN(new_n655));
  INV_X1    g0455(.A(G13), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(G1), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n261), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n261), .A2(new_n660), .A3(new_n657), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n659), .A2(G213), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n559), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n633), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n574), .A2(new_n577), .ZN(new_n666));
  INV_X1    g0466(.A(new_n569), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(KEYINPUT83), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT83), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n578), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n655), .B(new_n665), .C1(new_n672), .C2(new_n664), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n668), .A2(KEYINPUT83), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n578), .A2(new_n670), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n664), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n665), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT84), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n663), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n607), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n616), .A2(new_n681), .A3(new_n621), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n607), .A2(new_n615), .A3(new_n680), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n679), .A2(G330), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n569), .A2(new_n663), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n616), .A3(new_n621), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n607), .A2(new_n615), .A3(new_n663), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(G399));
  NOR2_X1   g0492(.A1(new_n213), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G1), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n422), .A2(new_n551), .A3(new_n464), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n695), .A2(new_n696), .B1(new_n236), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n565), .A2(new_n435), .ZN(new_n699));
  AND4_X1   g0499(.A1(new_n612), .A2(new_n611), .A3(new_n451), .A4(new_n478), .ZN(new_n700));
  INV_X1    g0500(.A(new_n525), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n699), .A2(new_n700), .A3(KEYINPUT30), .A4(new_n701), .ZN(new_n705));
  AOI21_X1  g0505(.A(G179), .B1(new_n478), .B2(new_n451), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n613), .A2(new_n525), .A3(new_n565), .A4(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n708), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT31), .B1(new_n708), .B2(new_n680), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n622), .B2(new_n680), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n616), .A2(new_n667), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n621), .A2(new_n628), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT85), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n528), .A2(new_n535), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n717), .B1(new_n528), .B2(new_n535), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n715), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n481), .A2(new_n487), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT75), .ZN(new_n723));
  INV_X1    g0523(.A(new_n528), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n637), .A3(new_n488), .A4(new_n724), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n504), .A2(new_n510), .B1(new_n525), .B2(new_n353), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(new_n487), .A3(new_n626), .A4(new_n527), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n635), .B1(new_n727), .B2(KEYINPUT26), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(KEYINPUT86), .B(new_n680), .C1(new_n721), .C2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT86), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n536), .A2(KEYINPUT85), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n528), .A2(new_n535), .A3(new_n717), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(new_n621), .A3(new_n628), .A4(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n569), .B1(new_n607), .B2(new_n615), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n725), .B(new_n728), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n731), .B1(new_n736), .B2(new_n663), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT29), .B1(new_n730), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n641), .A2(new_n663), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT29), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n714), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n698), .B1(new_n742), .B2(G1), .ZN(G364));
  NOR2_X1   g0543(.A1(new_n213), .A2(new_n260), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n744), .A2(G355), .B1(new_n551), .B2(new_n213), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n213), .A2(new_n317), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G45), .B2(new_n236), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n251), .A2(new_n303), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(G20), .B1(KEYINPUT88), .B2(G169), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(KEYINPUT88), .A2(G169), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n281), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n749), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n232), .A2(new_n656), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G45), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n694), .A2(G1), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT87), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n435), .A2(new_n617), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT89), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n261), .B1(new_n765), .B2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(KEYINPUT91), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT91), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n768), .B(new_n261), .C1(new_n765), .C2(G190), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT92), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n767), .A2(new_n769), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT92), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n225), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n261), .A2(G190), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n617), .A2(G179), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT90), .Z(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G107), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n779), .A2(G20), .A3(G190), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n435), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n778), .A2(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n317), .B1(new_n588), .B2(new_n783), .C1(new_n785), .C2(new_n219), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n765), .A2(new_n778), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G159), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n786), .B1(KEYINPUT32), .B2(new_n789), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(KEYINPUT32), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n435), .A2(new_n617), .ZN(new_n792));
  AND3_X1   g0592(.A1(new_n232), .A2(G190), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n778), .A2(new_n792), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n794), .A2(new_n201), .B1(new_n795), .B2(new_n234), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n232), .A2(G190), .A3(new_n784), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(G58), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n782), .A2(new_n790), .A3(new_n791), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n777), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(KEYINPUT93), .ZN(new_n803));
  INV_X1    g0603(.A(G329), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n787), .A2(new_n804), .B1(new_n785), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G322), .A2(new_n798), .B1(new_n793), .B2(G326), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n783), .B(KEYINPUT94), .Z(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G303), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n260), .B(new_n807), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n795), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT33), .B(G317), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n806), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G283), .ZN(new_n815));
  INV_X1    g0615(.A(new_n781), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n814), .B1(new_n815), .B2(new_n816), .C1(new_n817), .C2(new_n773), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n802), .A2(KEYINPUT93), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n803), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n758), .B(new_n763), .C1(new_n820), .C2(new_n753), .ZN(new_n821));
  INV_X1    g0621(.A(new_n756), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n679), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G330), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n673), .A2(new_n678), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n679), .A2(G330), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n826), .A3(new_n763), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NAND2_X1  g0629(.A1(new_n680), .A2(new_n417), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n648), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT96), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n437), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n434), .A2(KEYINPUT96), .A3(new_n417), .A4(new_n436), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n433), .A2(new_n830), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT97), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n831), .B1(new_n430), .B2(new_n432), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT97), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n839), .A2(new_n834), .A3(new_n840), .A4(new_n835), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n832), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n739), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n842), .B(new_n663), .C1(new_n634), .C2(new_n640), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n762), .B1(new_n846), .B2(new_n713), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n713), .B2(new_n846), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n753), .A2(new_n754), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n762), .B1(G77), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n812), .A2(KEYINPUT95), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n812), .A2(KEYINPUT95), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(G283), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n317), .B1(new_n793), .B2(G303), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n809), .A2(new_n221), .B1(new_n551), .B2(new_n785), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n787), .A2(new_n805), .B1(new_n817), .B2(new_n797), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n781), .A2(G87), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n856), .A2(new_n857), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n812), .A2(G150), .B1(G137), .B2(new_n793), .ZN(new_n863));
  INV_X1    g0663(.A(G143), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n863), .B1(new_n864), .B2(new_n797), .C1(new_n271), .C2(new_n785), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT34), .Z(new_n866));
  OAI21_X1  g0666(.A(new_n317), .B1(new_n809), .B2(new_n201), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(G132), .B2(new_n788), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n781), .A2(G68), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n868), .B(new_n869), .C1(new_n202), .C2(new_n773), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n777), .A2(new_n862), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n851), .B1(new_n871), .B2(new_n753), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n842), .B2(new_n755), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n848), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(G384));
  NOR2_X1   g0675(.A1(new_n233), .A2(new_n551), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n495), .A2(new_n499), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT35), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  NAND2_X1  g0681(.A1(new_n266), .A2(new_n268), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n235), .A2(G50), .A3(G77), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n882), .A2(new_n883), .B1(G50), .B2(new_n234), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(G1), .A3(new_n656), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT98), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n738), .A2(new_n741), .A3(new_n624), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n653), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n662), .B(KEYINPUT99), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n646), .B2(new_n647), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n406), .B1(new_n401), .B2(KEYINPUT14), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n404), .B1(new_n403), .B2(G169), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n408), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n408), .A2(new_n680), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n399), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n408), .B(new_n680), .C1(new_n407), .C2(new_n400), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n836), .A2(new_n663), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n899), .B1(new_n845), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT16), .B1(new_n288), .B2(new_n289), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n300), .B1(new_n330), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n662), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n341), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n335), .A2(new_n890), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n325), .A2(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n291), .A2(new_n300), .B1(new_n327), .B2(new_n328), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n903), .B1(new_n329), .B2(new_n662), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(KEYINPUT37), .A3(new_n325), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n906), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n904), .B1(new_n326), .B2(new_n340), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n917), .B1(new_n918), .B2(new_n914), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n891), .B1(new_n901), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n407), .A2(new_n408), .A3(new_n663), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n916), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n326), .A2(new_n646), .A3(new_n647), .ZN(new_n925));
  INV_X1    g0725(.A(new_n908), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n325), .A2(new_n908), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n325), .A2(new_n908), .A3(new_n643), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n336), .A2(new_n928), .B1(new_n929), .B2(KEYINPUT37), .ZN(new_n930));
  NOR4_X1   g0730(.A1(new_n909), .A2(new_n643), .A3(new_n910), .A4(new_n907), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT38), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n918), .A2(new_n914), .A3(new_n917), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n923), .B(new_n924), .C1(new_n935), .C2(KEYINPUT39), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n921), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n889), .B(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n622), .A2(new_n680), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n708), .A2(new_n680), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT31), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n708), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n842), .B(new_n898), .C1(new_n939), .C2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT40), .B1(new_n935), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n898), .A2(new_n842), .ZN(new_n947));
  INV_X1    g0747(.A(new_n939), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n947), .B1(new_n948), .B2(new_n711), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT40), .B1(new_n916), .B2(new_n919), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n439), .B1(new_n948), .B2(new_n711), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n824), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n938), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n208), .B2(new_n759), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n938), .A2(new_n955), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n887), .B1(new_n957), .B2(new_n958), .ZN(G367));
  NAND2_X1  g0759(.A1(new_n760), .A2(G1), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n679), .A2(G330), .A3(new_n684), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n533), .A2(new_n663), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n720), .A2(new_n963), .B1(new_n724), .B2(new_n680), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n690), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n690), .A2(new_n964), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n961), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n685), .A2(new_n966), .A3(new_n969), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n688), .B1(new_n684), .B2(new_n687), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n826), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n679), .A2(G330), .A3(new_n974), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n742), .B1(new_n973), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n693), .B(KEYINPUT41), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n960), .B1(new_n981), .B2(KEYINPUT103), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT103), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n979), .A2(new_n983), .A3(new_n980), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n663), .B1(new_n484), .B2(new_n485), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n626), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n628), .B2(new_n986), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT100), .Z(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n964), .A2(new_n688), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT42), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n720), .A2(new_n963), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n528), .B1(new_n993), .B2(new_n616), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n663), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n991), .A2(KEYINPUT42), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n992), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT101), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(KEYINPUT101), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n990), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(KEYINPUT102), .B1(new_n685), .B2(new_n964), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT102), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n964), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n961), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n989), .B(KEYINPUT43), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n998), .A2(new_n1006), .A3(new_n999), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1001), .A2(new_n1002), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1005), .A2(new_n1002), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1007), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n1010), .B2(new_n1000), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n985), .A2(new_n1013), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n746), .A2(new_n247), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n757), .B1(new_n212), .B2(new_n411), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n762), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n780), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(G97), .ZN(new_n1019));
  INV_X1    g0819(.A(G317), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(KEYINPUT104), .B(G311), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n787), .A2(new_n1020), .B1(new_n794), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n785), .A2(new_n815), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n783), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT46), .B1(new_n1024), .B2(G116), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1022), .A2(new_n317), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n808), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n798), .A2(G303), .ZN(new_n1028));
  AND4_X1   g0828(.A1(new_n1019), .A2(new_n1026), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n817), .B2(new_n854), .C1(new_n422), .C2(new_n773), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n785), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n855), .A2(G159), .B1(G50), .B2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT105), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(KEYINPUT105), .ZN(new_n1034));
  INV_X1    g0834(.A(G137), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n787), .A2(new_n1035), .B1(new_n780), .B2(new_n219), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n317), .B1(new_n202), .B2(new_n783), .C1(new_n794), .C2(new_n864), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(G150), .C2(new_n798), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1033), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n776), .A2(new_n234), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1030), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT47), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1017), .B1(new_n1042), .B2(new_n753), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n822), .B2(new_n989), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1014), .A2(new_n1044), .ZN(G387));
  NAND2_X1  g0845(.A1(new_n976), .A2(new_n977), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n694), .B1(new_n1046), .B2(new_n742), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n742), .B2(new_n1046), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n960), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n753), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n317), .B1(new_n219), .B2(new_n783), .C1(new_n787), .C2(new_n357), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n781), .B2(G97), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT106), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n775), .A2(new_n473), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1031), .A2(G68), .B1(G50), .B2(new_n798), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n292), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n812), .A2(new_n1056), .B1(G159), .B2(new_n793), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n317), .B1(new_n788), .B2(G326), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G317), .A2(new_n798), .B1(new_n793), .B2(G322), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n810), .B2(new_n785), .C1(new_n854), .C2(new_n1021), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n770), .A2(G283), .B1(G294), .B2(new_n1024), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT49), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1059), .B1(new_n551), .B2(new_n780), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1058), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1050), .B1(new_n1070), .B2(KEYINPUT107), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(KEYINPUT107), .B2(new_n1070), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n746), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n244), .B2(G45), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n696), .B2(new_n744), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1056), .A2(new_n201), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT50), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n303), .B1(new_n234), .B2(new_n219), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1077), .A2(new_n696), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1075), .A2(new_n1079), .B1(G107), .B2(new_n212), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n763), .B1(new_n1080), .B2(new_n757), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1072), .B(new_n1081), .C1(new_n684), .C2(new_n822), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1049), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT108), .B1(new_n1048), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1048), .A2(new_n1083), .A3(KEYINPUT108), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(G393));
  NOR2_X1   g0887(.A1(new_n1073), .A2(new_n254), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n757), .B1(new_n225), .B2(new_n212), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G311), .A2(new_n798), .B1(new_n793), .B2(G317), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n260), .B1(new_n783), .B2(new_n815), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n785), .A2(new_n817), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(G322), .C2(new_n788), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1094), .B(new_n782), .C1(new_n810), .C2(new_n854), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1091), .B(new_n1095), .C1(G116), .C2(new_n770), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n775), .A2(G77), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1097), .B1(new_n201), .B2(new_n854), .C1(new_n292), .C2(new_n785), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT110), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n260), .B1(new_n1024), .B2(G68), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n861), .B(new_n1100), .C1(new_n864), .C2(new_n787), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G159), .A2(new_n798), .B1(new_n793), .B2(G150), .ZN(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n1103));
  XNOR2_X1  g0903(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1096), .B1(new_n1099), .B2(new_n1105), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n762), .B1(new_n1088), .B2(new_n1089), .C1(new_n1106), .C2(new_n1050), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT111), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n964), .A2(new_n756), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n971), .A2(new_n972), .A3(new_n960), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT112), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1112), .A2(KEYINPUT112), .A3(new_n1113), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n742), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n978), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n973), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n694), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n973), .B1(new_n978), .B2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1118), .A2(new_n1124), .ZN(G390));
  NAND2_X1  g0925(.A1(new_n927), .A2(new_n932), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n917), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT39), .B1(new_n1127), .B2(new_n916), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n924), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n1128), .A2(new_n1129), .B1(new_n901), .B2(new_n923), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n842), .B1(new_n730), .B2(new_n737), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n899), .B1(new_n1131), .B2(new_n900), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n922), .B1(new_n933), .B2(new_n934), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(G330), .B(new_n842), .C1(new_n939), .C2(new_n944), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(new_n899), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n712), .A2(G330), .A3(new_n842), .A4(new_n898), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1130), .B(new_n1138), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT113), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n714), .A2(new_n624), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n888), .A2(new_n653), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1135), .A2(new_n899), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1138), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n845), .A2(new_n900), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1144), .A2(new_n1131), .A3(new_n1138), .A4(new_n900), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1140), .B(new_n1141), .C1(new_n1143), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1140), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1141), .B1(new_n1149), .B2(new_n1143), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1150), .A2(new_n693), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n754), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n762), .B1(new_n1056), .B2(new_n850), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n776), .A2(new_n271), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n855), .A2(G137), .ZN(new_n1158));
  INV_X1    g0958(.A(G125), .ZN(new_n1159));
  INV_X1    g0959(.A(G128), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1159), .A2(new_n787), .B1(new_n794), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G50), .B2(new_n1018), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT53), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1024), .B2(G150), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n783), .A2(KEYINPUT53), .A3(new_n357), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1164), .A2(new_n260), .A3(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT54), .B(G143), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT114), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1031), .A2(new_n1168), .B1(G132), .B2(new_n798), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1158), .A2(new_n1162), .A3(new_n1166), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1097), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n855), .A2(new_n530), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n785), .A2(new_n225), .B1(new_n551), .B2(new_n797), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n794), .A2(new_n815), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(G87), .C2(new_n808), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n317), .B1(new_n788), .B2(G294), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1172), .A2(new_n1175), .A3(new_n869), .A4(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1157), .A2(new_n1170), .B1(new_n1171), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1156), .B1(new_n1178), .B2(new_n753), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT115), .Z(new_n1180));
  AOI22_X1  g0980(.A1(new_n1151), .A2(new_n960), .B1(new_n1155), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1154), .A2(new_n1181), .ZN(G378));
  INV_X1    g0982(.A(new_n960), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n947), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1184), .B(new_n712), .C1(new_n934), .C2(new_n933), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1185), .A2(KEYINPUT40), .B1(new_n949), .B2(new_n950), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n662), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n365), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n374), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n374), .A2(new_n1189), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OR3_X1    g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1194), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n1186), .A2(new_n1197), .A3(new_n824), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n952), .B2(G330), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n937), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1197), .B1(new_n1186), .B2(new_n824), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n952), .A2(G330), .A3(new_n1199), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n937), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1183), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n317), .A2(G41), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n780), .A2(new_n202), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT116), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1207), .B1(new_n219), .B2(new_n783), .C1(new_n797), .C2(new_n221), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n225), .A2(new_n795), .B1(new_n785), .B2(new_n411), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G283), .C2(new_n788), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1040), .B1(G116), .B2(new_n793), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT117), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(KEYINPUT117), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1211), .B(new_n1214), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT58), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1209), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1219), .B2(new_n1218), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n785), .A2(new_n1035), .B1(new_n1160), .B2(new_n797), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1168), .A2(new_n1024), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1159), .B2(new_n794), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(G132), .C2(new_n812), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n776), .B2(new_n357), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT119), .ZN(new_n1227));
  XOR2_X1   g1027(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1228));
  XNOR2_X1  g1028(.A(new_n1227), .B(new_n1228), .ZN(new_n1229));
  AOI211_X1 g1029(.A(G33), .B(G41), .C1(new_n788), .C2(G124), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n271), .B2(new_n780), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n753), .B1(new_n1221), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1197), .A2(new_n754), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n763), .B1(new_n201), .B2(new_n849), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1206), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1137), .A2(new_n1139), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1143), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT120), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1240), .A2(KEYINPUT120), .A3(new_n1241), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT57), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT57), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1240), .A2(KEYINPUT120), .A3(new_n1241), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT120), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1250), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n693), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1238), .B1(new_n1248), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT121), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1238), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n694), .B1(new_n1246), .B2(new_n1250), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1247), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1249), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1258), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT121), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1257), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(G375));
  OAI21_X1  g1065(.A(new_n762), .B1(G68), .B2(new_n850), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n776), .A2(new_n201), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n855), .A2(new_n1168), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n260), .B1(new_n793), .B2(G132), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n785), .A2(new_n357), .B1(new_n1035), .B2(new_n797), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n787), .A2(new_n1160), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1270), .B(new_n1271), .C1(G159), .C2(new_n808), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1268), .A2(new_n1211), .A3(new_n1269), .A4(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1054), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n855), .A2(G116), .B1(G77), .B2(new_n781), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n317), .B1(new_n793), .B2(G294), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n808), .A2(G97), .B1(G283), .B2(new_n798), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n788), .A2(G303), .B1(new_n1031), .B2(new_n530), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n1267), .A2(new_n1273), .B1(new_n1274), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1266), .B1(new_n1280), .B2(new_n753), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n898), .B2(new_n755), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1149), .B2(new_n1183), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n980), .B1(new_n1149), .B2(new_n1143), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1149), .A2(new_n1143), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1284), .B1(new_n1285), .B2(new_n1287), .ZN(G381));
  AOI21_X1  g1088(.A(new_n1012), .B1(new_n982), .B2(new_n984), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1044), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1289), .A2(G390), .A3(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1085), .A2(new_n828), .A3(new_n1086), .ZN(new_n1292));
  NOR4_X1   g1092(.A1(G378), .A2(new_n1292), .A3(G384), .A4(G381), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1264), .A2(new_n1291), .A3(new_n1293), .ZN(G407));
  INV_X1    g1094(.A(G378), .ZN(new_n1295));
  INV_X1    g1095(.A(G343), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(G213), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1297), .B(KEYINPUT122), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1264), .A2(new_n1295), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(G407), .A2(new_n1299), .A3(G213), .ZN(G409));
  OAI21_X1  g1100(.A(G390), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n1116), .A2(new_n1117), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n984), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n983), .B1(new_n979), .B2(new_n980), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n960), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1044), .B(new_n1302), .C1(new_n1305), .C2(new_n1012), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1086), .ZN(new_n1307));
  OAI21_X1  g1107(.A(G396), .B1(new_n1307), .B2(new_n1084), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1292), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1301), .A2(new_n1306), .A3(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1309), .B1(new_n1301), .B2(new_n1306), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G378), .B(new_n1238), .C1(new_n1248), .C2(new_n1254), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT123), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1206), .A2(new_n1315), .A3(new_n1237), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1204), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n960), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT123), .B1(new_n1319), .B2(new_n1236), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1316), .A2(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n980), .B(new_n1247), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1295), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1314), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1298), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1143), .A2(new_n1147), .A3(KEYINPUT60), .A4(new_n1148), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n693), .ZN(new_n1328));
  OAI21_X1  g1128(.A(KEYINPUT60), .B1(new_n1149), .B2(new_n1143), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1286), .B2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n874), .B1(new_n1330), .B2(new_n1283), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT124), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT124), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1333), .B(new_n874), .C1(new_n1330), .C2(new_n1283), .ZN(new_n1334));
  OR3_X1    g1134(.A1(new_n1330), .A2(new_n874), .A3(new_n1283), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1332), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1325), .A2(new_n1326), .A3(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT125), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1325), .A2(KEYINPUT125), .A3(new_n1326), .A4(new_n1337), .ZN(new_n1341));
  AOI21_X1  g1141(.A(KEYINPUT62), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1298), .A2(G2897), .ZN(new_n1343));
  NOR3_X1   g1143(.A1(new_n1330), .A2(new_n874), .A3(new_n1283), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1344), .B1(KEYINPUT124), .B2(new_n1331), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1343), .B1(new_n1345), .B2(new_n1334), .ZN(new_n1346));
  AND4_X1   g1146(.A1(new_n1334), .A2(new_n1332), .A3(new_n1335), .A4(new_n1343), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(G378), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1349), .B1(new_n1262), .B2(G378), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1348), .B1(new_n1350), .B2(new_n1298), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT61), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT62), .ZN(new_n1353));
  AOI211_X1 g1153(.A(new_n1298), .B(new_n1336), .C1(new_n1314), .C2(new_n1324), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1351), .B(new_n1352), .C1(new_n1353), .C2(new_n1354), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1313), .B1(new_n1342), .B2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT63), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1340), .A2(new_n1357), .A3(new_n1341), .ZN(new_n1358));
  AND2_X1   g1158(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1354), .A2(KEYINPUT63), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1358), .A2(new_n1359), .A3(new_n1312), .A4(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1356), .A2(new_n1361), .ZN(G405));
  NAND3_X1  g1162(.A1(new_n1257), .A2(new_n1263), .A3(new_n1295), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT126), .ZN(new_n1364));
  AOI22_X1  g1164(.A1(new_n1364), .A2(new_n1337), .B1(new_n1262), .B2(G378), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1363), .A2(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1366), .A2(KEYINPUT127), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1336), .A2(KEYINPUT126), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1368), .ZN(new_n1369));
  OAI21_X1  g1169(.A(new_n1369), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1301), .A2(new_n1306), .ZN(new_n1371));
  INV_X1    g1171(.A(new_n1309), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1301), .A2(new_n1306), .A3(new_n1309), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1373), .A2(new_n1374), .A3(new_n1368), .ZN(new_n1375));
  AND2_X1   g1175(.A1(new_n1370), .A2(new_n1375), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT127), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1363), .A2(new_n1365), .A3(new_n1377), .ZN(new_n1378));
  AND3_X1   g1178(.A1(new_n1367), .A2(new_n1376), .A3(new_n1378), .ZN(new_n1379));
  AOI21_X1  g1179(.A(new_n1376), .B1(new_n1367), .B2(new_n1378), .ZN(new_n1380));
  NOR2_X1   g1180(.A1(new_n1379), .A2(new_n1380), .ZN(G402));
endmodule


