//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n639,
    new_n640, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G235), .A3(G237), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT72), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT71), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n462), .B(new_n468), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(G101), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT73), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n465), .A2(KEYINPUT3), .A3(new_n466), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n476), .A2(new_n480), .A3(G137), .A4(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n474), .A2(new_n475), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G101), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT72), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(new_n487), .B2(new_n472), .ZN(new_n488));
  AND4_X1   g063(.A1(G137), .A2(new_n476), .A3(new_n480), .A4(new_n482), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT73), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n480), .ZN(new_n492));
  NAND2_X1  g067(.A1(G113), .A2(G2104), .ZN(new_n493));
  INV_X1    g068(.A(G125), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n481), .A2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n482), .A2(new_n499), .A3(KEYINPUT69), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n493), .B1(new_n501), .B2(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  AOI211_X1 g078(.A(new_n503), .B(new_n494), .C1(new_n498), .C2(new_n500), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n492), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n491), .A2(new_n505), .ZN(G160));
  AND2_X1   g081(.A1(new_n476), .A2(new_n482), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(new_n468), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n476), .A2(new_n482), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT74), .B1(new_n510), .B2(G2105), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G136), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT75), .ZN(new_n514));
  OAI221_X1 g089(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n480), .C2(G112), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(new_n492), .ZN(new_n516));
  INV_X1    g091(.A(G124), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n514), .A2(new_n518), .ZN(G162));
  NAND2_X1  g094(.A1(G126), .A2(G2105), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n468), .A2(G114), .ZN(new_n521));
  OAI21_X1  g096(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n510), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G138), .ZN(new_n524));
  NOR3_X1   g099(.A1(new_n478), .A2(new_n479), .A3(new_n524), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n526));
  AND3_X1   g101(.A1(new_n482), .A2(new_n499), .A3(KEYINPUT69), .ZN(new_n527));
  AOI21_X1  g102(.A(KEYINPUT69), .B1(new_n482), .B2(new_n499), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n525), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n525), .A2(new_n482), .A3(new_n476), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n529), .A2(KEYINPUT77), .B1(KEYINPUT4), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n498), .A2(new_n500), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n532), .A2(new_n533), .A3(new_n525), .A4(new_n526), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n523), .B1(new_n531), .B2(new_n534), .ZN(G164));
  XNOR2_X1  g110(.A(KEYINPUT5), .B(G543), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n536), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT6), .B(G651), .Z(new_n538));
  OAI21_X1  g113(.A(KEYINPUT78), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n536), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR3_X1   g117(.A1(new_n537), .A2(KEYINPUT78), .A3(new_n538), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(new_n543), .ZN(G303));
  INV_X1    g119(.A(G303), .ZN(G166));
  INV_X1    g120(.A(KEYINPUT80), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g122(.A(KEYINPUT6), .B(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT80), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n547), .A2(G543), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G51), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT81), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n536), .B(KEYINPUT79), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n553), .A2(G63), .A3(G651), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n536), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n538), .ZN(new_n557));
  NAND3_X1  g132(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT7), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n558), .A2(KEYINPUT7), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n557), .A2(G89), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n552), .B1(new_n551), .B2(new_n554), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT82), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n563), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT82), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n565), .A2(new_n566), .A3(new_n555), .A4(new_n561), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G168));
  NAND2_X1  g143(.A1(new_n553), .A2(G64), .ZN(new_n569));
  NAND2_X1  g144(.A1(G77), .A2(G543), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n540), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n557), .A2(G90), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n547), .A2(G543), .A3(new_n549), .ZN(new_n573));
  INV_X1    g148(.A(G52), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n571), .A2(new_n575), .ZN(G171));
  NAND2_X1  g151(.A1(G68), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n536), .B(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(G56), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  XNOR2_X1  g157(.A(KEYINPUT83), .B(G81), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n550), .A2(G43), .B1(new_n557), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G860), .ZN(G153));
  NAND4_X1  g162(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g163(.A1(G1), .A2(G3), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT8), .ZN(new_n590));
  NAND4_X1  g165(.A1(G319), .A2(G483), .A3(G661), .A4(new_n590), .ZN(G188));
  NAND4_X1  g166(.A1(new_n547), .A2(G53), .A3(G543), .A4(new_n549), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(KEYINPUT9), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(KEYINPUT9), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G78), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G65), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n556), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n557), .A2(G91), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n595), .A2(new_n602), .ZN(G299));
  INV_X1    g178(.A(G171), .ZN(G301));
  AND2_X1   g179(.A1(new_n564), .A2(new_n567), .ZN(G286));
  OAI21_X1  g180(.A(G651), .B1(new_n553), .B2(G74), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(KEYINPUT84), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n550), .A2(G49), .B1(G87), .B2(new_n557), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n609), .B(G651), .C1(new_n553), .C2(G74), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(G288));
  AOI22_X1  g186(.A1(new_n536), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(new_n540), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n536), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(new_n538), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT85), .ZN(G305));
  NAND2_X1  g192(.A1(G72), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G60), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n579), .B2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n540), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n621), .B2(new_n620), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n550), .A2(G47), .B1(G85), .B2(new_n557), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(G290));
  AND3_X1   g200(.A1(new_n536), .A2(new_n548), .A3(G92), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT10), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n550), .A2(G54), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n536), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(new_n540), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G868), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(G171), .ZN(G284));
  OAI21_X1  g209(.A(new_n633), .B1(new_n632), .B2(G171), .ZN(G321));
  NOR2_X1   g210(.A1(G299), .A2(G868), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g212(.A(new_n636), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g213(.A(new_n631), .ZN(new_n639));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G860), .ZN(G148));
  NAND2_X1  g216(.A1(new_n585), .A2(new_n632), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n631), .A2(G559), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(new_n632), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g220(.A1(new_n487), .A2(new_n472), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(new_n532), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT12), .Z(new_n648));
  XOR2_X1   g223(.A(KEYINPUT87), .B(KEYINPUT13), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(G2100), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(G2100), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n512), .A2(G135), .ZN(new_n653));
  OAI221_X1 g228(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n480), .C2(G111), .ZN(new_n654));
  INV_X1    g229(.A(G123), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n516), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n652), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT88), .ZN(G156));
  XNOR2_X1  g235(.A(G2427), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(KEYINPUT14), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2451), .B(G2454), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  OR2_X1    g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(G14), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n670), .B2(new_n673), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(G401));
  INV_X1    g252(.A(KEYINPUT18), .ZN(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(KEYINPUT17), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G2072), .B(G2078), .Z(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n681), .B2(KEYINPUT18), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT90), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(G227));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT19), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n697), .A2(new_n698), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n696), .A2(new_n699), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n696), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G1981), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n708), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n693), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n713), .A2(new_n709), .A3(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT91), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n712), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n712), .B2(new_n714), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n692), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n712), .A2(new_n714), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(new_n716), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n712), .A2(new_n714), .A3(new_n717), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n722), .A2(new_n723), .A3(new_n691), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(new_n724), .ZN(G229));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G24), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n623), .A2(new_n624), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n726), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G1986), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n693), .B(new_n727), .C1(new_n728), .C2(new_n726), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G25), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n512), .A2(G131), .ZN(new_n734));
  INV_X1    g309(.A(new_n516), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G119), .ZN(new_n736));
  OAI221_X1 g311(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n480), .C2(G107), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(new_n732), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n740), .A2(new_n742), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n730), .A2(new_n731), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n726), .A2(G23), .ZN(new_n746));
  INV_X1    g321(.A(G288), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(new_n726), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT33), .B(G1976), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT32), .B(G1981), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT85), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n616), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G16), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G6), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n751), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n751), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n754), .B(new_n758), .C1(G6), .C2(G16), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n726), .A2(G22), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G303), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1971), .ZN(new_n763));
  AND3_X1   g338(.A1(new_n750), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n745), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT36), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n750), .A2(new_n760), .A3(new_n763), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n770));
  INV_X1    g345(.A(new_n765), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n766), .B(new_n768), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  AND3_X1   g350(.A1(new_n730), .A2(new_n743), .A3(new_n744), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n776), .B(new_n731), .C1(new_n769), .C2(new_n771), .ZN(new_n777));
  INV_X1    g352(.A(new_n774), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(new_n772), .ZN(new_n779));
  INV_X1    g354(.A(new_n768), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n775), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(G16), .A2(G21), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G286), .B2(new_n726), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT101), .B(G1966), .Z(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n732), .A2(G26), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT28), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n512), .A2(G140), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n480), .A2(G116), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n735), .A2(G128), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(G29), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2067), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n785), .A2(new_n786), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n787), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n732), .A2(G32), .ZN(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT26), .Z(new_n804));
  INV_X1    g379(.A(G129), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n516), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G141), .B2(new_n512), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n646), .A2(G105), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT99), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n802), .B1(new_n811), .B2(new_n732), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT27), .B(G1996), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT25), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n532), .A2(G127), .ZN(new_n818));
  INV_X1    g393(.A(G115), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n464), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n817), .B1(new_n820), .B2(new_n492), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n512), .A2(G139), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G29), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n732), .A2(G33), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n815), .B1(G2072), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(G160), .A2(G29), .ZN(new_n828));
  INV_X1    g403(.A(G34), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(KEYINPUT24), .ZN(new_n830));
  AOI21_X1  g405(.A(G29), .B1(new_n829), .B2(KEYINPUT24), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(KEYINPUT98), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(KEYINPUT98), .B2(new_n831), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n828), .A2(G2084), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n827), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n826), .A2(G2072), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT97), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n801), .B1(new_n838), .B2(KEYINPUT100), .ZN(new_n839));
  NOR2_X1   g414(.A1(G171), .A2(new_n726), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G5), .B2(new_n726), .ZN(new_n841));
  INV_X1    g416(.A(G1961), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(G2084), .B1(new_n828), .B2(new_n833), .ZN(new_n844));
  NOR2_X1   g419(.A1(G4), .A2(G16), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n639), .B2(G16), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(G1348), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n846), .A2(G1348), .ZN(new_n848));
  NOR4_X1   g423(.A1(new_n843), .A2(new_n844), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G11), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT31), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(KEYINPUT31), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT30), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n853), .A2(G28), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n732), .B1(new_n853), .B2(G28), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n851), .B(new_n852), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n657), .B2(G29), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n585), .A2(G16), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n726), .A2(G19), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT95), .Z(new_n860));
  AND3_X1   g435(.A1(new_n858), .A2(G1341), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(G1341), .B1(new_n858), .B2(new_n860), .ZN(new_n862));
  OAI221_X1 g437(.A(new_n857), .B1(new_n861), .B2(new_n862), .C1(new_n841), .C2(new_n842), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT102), .B(KEYINPUT23), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n726), .A2(G20), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(G299), .B2(G16), .ZN(new_n868));
  INV_X1    g443(.A(G1956), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n812), .B2(new_n814), .ZN(new_n871));
  NOR2_X1   g446(.A1(G27), .A2(G29), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(G164), .B2(G29), .ZN(new_n873));
  INV_X1    g448(.A(G2078), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n849), .A2(new_n864), .A3(new_n871), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n732), .A2(G35), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(G162), .B2(new_n732), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT29), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(G2090), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(G2090), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n835), .B2(new_n837), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n839), .A2(new_n881), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n783), .A2(new_n885), .ZN(G311));
  OAI21_X1  g461(.A(KEYINPUT103), .B1(new_n783), .B2(new_n885), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n836), .B(KEYINPUT97), .Z(new_n888));
  NAND4_X1  g463(.A1(new_n888), .A2(KEYINPUT100), .A3(new_n834), .A4(new_n827), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n787), .A2(new_n800), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n884), .A2(new_n889), .A3(new_n890), .A4(new_n799), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n879), .A2(G2090), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n849), .A2(new_n871), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n864), .A2(new_n875), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n882), .A4(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n766), .B1(new_n773), .B2(new_n774), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(new_n780), .A3(new_n781), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n896), .A2(new_n897), .A3(new_n899), .A4(new_n775), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n887), .A2(new_n900), .ZN(G150));
  NAND2_X1  g476(.A1(new_n553), .A2(G67), .ZN(new_n902));
  NAND2_X1  g477(.A1(G80), .A2(G543), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G651), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n557), .A2(G93), .ZN(new_n906));
  INV_X1    g481(.A(G55), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n906), .B1(new_n573), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n909), .A3(KEYINPUT104), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n540), .B1(new_n902), .B2(new_n903), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n911), .B1(new_n912), .B2(new_n908), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n585), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n585), .A2(new_n912), .A3(new_n908), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n631), .A2(new_n640), .ZN(new_n919));
  XOR2_X1   g494(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n920));
  XNOR2_X1  g495(.A(new_n919), .B(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n918), .B(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT39), .ZN(new_n923));
  AOI21_X1  g498(.A(G860), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(KEYINPUT106), .Z(new_n926));
  NAND2_X1  g501(.A1(new_n914), .A2(G860), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT37), .Z(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(G145));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n930), .B(new_n523), .C1(new_n531), .C2(new_n534), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n529), .A2(KEYINPUT77), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n530), .A2(KEYINPUT4), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n534), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n523), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT107), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n797), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n739), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n930), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n934), .A2(KEYINPUT107), .A3(new_n935), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n797), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n738), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n810), .B(new_n823), .ZN(new_n947));
  OAI21_X1  g522(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n948), .B(KEYINPUT109), .Z(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n480), .A2(G118), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n512), .A2(G142), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n735), .A2(G130), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(new_n648), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n947), .B(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n946), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(G160), .B(new_n657), .Z(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(G162), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n939), .A2(new_n958), .A3(new_n945), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT110), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n960), .A2(new_n966), .A3(new_n962), .A4(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n962), .B1(new_n960), .B2(new_n963), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(G37), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n968), .A2(KEYINPUT40), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT40), .B1(new_n968), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(G395));
  INV_X1    g548(.A(KEYINPUT114), .ZN(new_n974));
  XNOR2_X1  g549(.A(G290), .B(new_n753), .ZN(new_n975));
  XNOR2_X1  g550(.A(G288), .B(G303), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n976), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n728), .A2(new_n753), .ZN(new_n979));
  NOR2_X1   g554(.A1(G290), .A2(G305), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n977), .A2(KEYINPUT42), .A3(new_n981), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n586), .B1(new_n913), .B2(new_n910), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n643), .B1(new_n987), .B2(new_n916), .ZN(new_n988));
  INV_X1    g563(.A(new_n643), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n915), .A2(new_n989), .A3(new_n917), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(G299), .A2(new_n631), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n601), .B1(new_n593), .B2(new_n594), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n639), .A2(new_n993), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n992), .A2(KEYINPUT41), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT41), .B1(new_n992), .B2(new_n994), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT112), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n991), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G299), .A2(new_n631), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n639), .A2(new_n993), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n988), .A2(new_n990), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT111), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n988), .A2(new_n990), .A3(new_n1007), .A4(new_n1004), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n999), .A2(new_n1001), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n986), .B1(new_n1009), .B2(KEYINPUT113), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n999), .A2(new_n1001), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1011), .B(new_n986), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1016));
  AND4_X1   g591(.A1(new_n974), .A2(new_n1015), .A3(G868), .A4(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n914), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT114), .B1(new_n1018), .B2(G868), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n632), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(new_n1016), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1017), .A2(new_n1021), .ZN(G295));
  NOR2_X1   g597(.A1(new_n1017), .A2(new_n1021), .ZN(G331));
  AND3_X1   g598(.A1(new_n564), .A2(new_n567), .A3(G301), .ZN(new_n1024));
  AOI21_X1  g599(.A(G301), .B1(new_n564), .B2(new_n567), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n918), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G168), .A2(G171), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n987), .A2(new_n916), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n564), .A2(new_n567), .A3(G301), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n997), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1026), .A2(new_n1030), .A3(new_n1004), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(G37), .B1(new_n1034), .B2(new_n982), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n1037));
  INV_X1    g612(.A(new_n982), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1032), .A2(new_n1038), .A3(new_n1033), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1026), .A2(new_n1030), .A3(new_n1004), .ZN(new_n1041));
  INV_X1    g616(.A(new_n997), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(new_n1030), .B2(new_n1026), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n982), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G37), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1044), .A2(new_n1039), .A3(new_n1037), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT115), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1039), .A3(new_n1045), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT43), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1040), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT44), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(KEYINPUT44), .A3(new_n1046), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(G397));
  INV_X1    g629(.A(G1384), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n941), .A2(new_n1055), .A3(new_n942), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT45), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n491), .A2(new_n505), .A3(G40), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(new_n693), .A3(new_n728), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(G1986), .A3(G290), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT116), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n797), .A2(G2067), .ZN(new_n1065));
  INV_X1    g640(.A(G2067), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n792), .A2(new_n1066), .A3(new_n796), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(KEYINPUT117), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1996), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n810), .B(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n738), .B(new_n741), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1068), .A2(new_n1071), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1075), .A2(new_n1060), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1064), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n491), .A2(new_n505), .A3(G40), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1057), .B1(G164), .B2(G1384), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n940), .A2(KEYINPUT45), .A3(new_n1055), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n786), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n940), .A2(new_n1085), .A3(new_n1055), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1078), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1083), .B(G168), .C1(G2084), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G8), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(KEYINPUT122), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(KEYINPUT122), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1088), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1087), .A2(G2084), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1083), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(G8), .A3(G286), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1093), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT62), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1092), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n1097), .A4(new_n1094), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n940), .A2(new_n1055), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1059), .B1(new_n1057), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n941), .A2(KEYINPUT45), .A3(new_n1055), .A4(new_n942), .ZN(new_n1107));
  AOI21_X1  g682(.A(G1971), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1087), .A2(G2090), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G303), .A2(G8), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT55), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(G8), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1078), .A2(new_n1055), .A3(new_n940), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n747), .A2(G1976), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(G8), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT52), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1105), .A2(new_n1059), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(new_n1089), .ZN(new_n1120));
  INV_X1    g695(.A(G1976), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT52), .B1(G288), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1116), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n616), .A2(new_n708), .ZN(new_n1124));
  OAI21_X1  g699(.A(G1981), .B1(new_n613), .B2(new_n615), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1124), .B(new_n1125), .C1(KEYINPUT118), .C2(KEYINPUT49), .ZN(new_n1126));
  AND2_X1   g701(.A1(KEYINPUT118), .A2(KEYINPUT49), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1120), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1118), .A2(new_n1123), .A3(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(G8), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1112), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1114), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1106), .A2(new_n1107), .A3(new_n874), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1135), .A2(G2078), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1137), .A2(new_n1138), .B1(new_n1087), .B2(new_n842), .ZN(new_n1139));
  AOI21_X1  g714(.A(G301), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1100), .A2(new_n1104), .A3(new_n1133), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1114), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1129), .A2(new_n1121), .A3(new_n747), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1124), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1142), .A2(new_n1130), .B1(new_n1120), .B2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1087), .A2(new_n842), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1107), .A2(new_n1078), .A3(new_n1138), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT45), .B1(new_n937), .B2(new_n1055), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(G171), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT123), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1136), .A2(new_n1139), .A3(G301), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1153), .A2(KEYINPUT54), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1058), .A2(new_n1078), .A3(new_n1107), .A4(new_n1138), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1136), .A2(new_n1155), .A3(new_n1147), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(G171), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1152), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1102), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT54), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1156), .A2(G171), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n1162), .B2(new_n1140), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1159), .A2(new_n1133), .A3(new_n1160), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(G1348), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1087), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1119), .A2(new_n1066), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n631), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT56), .B(G2072), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1106), .A2(new_n1107), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1087), .A2(new_n869), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT57), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n993), .A2(KEYINPUT121), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1172), .A2(KEYINPUT121), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1172), .A2(KEYINPUT121), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n993), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1170), .A2(new_n1171), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1168), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1178), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1106), .A2(new_n1107), .A3(new_n1072), .ZN(new_n1185));
  XOR2_X1   g760(.A(KEYINPUT58), .B(G1341), .Z(new_n1186));
  NAND2_X1  g761(.A1(new_n1115), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n586), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT59), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1188), .A2(new_n1191), .A3(new_n586), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1183), .A2(new_n1184), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1166), .A2(KEYINPUT60), .A3(new_n631), .A4(new_n1167), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1166), .A2(KEYINPUT60), .A3(new_n1167), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n639), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT60), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1170), .A2(new_n1177), .A3(new_n1171), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n1199), .A2(new_n1180), .A3(new_n1184), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1182), .B1(new_n1193), .B2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n1141), .B(new_n1145), .C1(new_n1164), .C2(new_n1202), .ZN(new_n1203));
  AOI211_X1 g778(.A(new_n1089), .B(G286), .C1(new_n1095), .C2(new_n1083), .ZN(new_n1204));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n1133), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1114), .A2(KEYINPUT63), .A3(new_n1204), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1131), .A2(KEYINPUT119), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1112), .B1(new_n1131), .B2(KEYINPUT119), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1130), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1206), .B1(new_n1209), .B2(KEYINPUT120), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT120), .ZN(new_n1211));
  OAI211_X1 g786(.A(new_n1211), .B(new_n1130), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1205), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1077), .B1(new_n1203), .B2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n738), .A2(new_n742), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT124), .ZN(new_n1216));
  NAND4_X1  g791(.A1(new_n1071), .A2(new_n1068), .A3(new_n1073), .A4(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1217), .A2(new_n1067), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(new_n1060), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1219), .B(KEYINPUT125), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1071), .A2(new_n811), .A3(new_n1068), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1221), .A2(new_n1060), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1060), .A2(new_n1072), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n1223), .B(KEYINPUT46), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT47), .ZN(new_n1225));
  AND3_X1   g800(.A1(new_n1222), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1225), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1227));
  XNOR2_X1  g802(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1228));
  XNOR2_X1  g803(.A(new_n1061), .B(new_n1228), .ZN(new_n1229));
  OAI22_X1  g804(.A1(new_n1226), .A2(new_n1227), .B1(new_n1076), .B2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1220), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1214), .A2(new_n1231), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g807(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1234));
  NAND3_X1  g808(.A1(new_n720), .A2(new_n724), .A3(new_n1234), .ZN(new_n1235));
  OR2_X1    g809(.A1(new_n1235), .A2(KEYINPUT127), .ZN(new_n1236));
  NAND2_X1  g810(.A1(new_n1235), .A2(KEYINPUT127), .ZN(new_n1237));
  AOI22_X1  g811(.A1(new_n968), .A2(new_n970), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AND2_X1   g812(.A1(new_n1238), .A2(new_n1050), .ZN(G308));
  NAND2_X1  g813(.A1(new_n1238), .A2(new_n1050), .ZN(G225));
endmodule


