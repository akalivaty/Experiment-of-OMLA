//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1272, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AND2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT1), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n211), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n203), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n218), .B(new_n224), .C1(new_n213), .C2(new_n212), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n215), .A2(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G68), .B(G77), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT65), .B(G50), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G41), .ZN(new_n243));
  INV_X1    g0043(.A(G45), .ZN(new_n244));
  AOI21_X1  g0044(.A(G1), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G1), .A3(G13), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n245), .A2(new_n247), .A3(G274), .ZN(new_n248));
  INV_X1    g0048(.A(G244), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n248), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G107), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n255), .B(new_n257), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G232), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT3), .B(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G238), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n259), .B1(new_n262), .B2(new_n263), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n267), .A2(KEYINPUT68), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n247), .B1(new_n267), .B2(KEYINPUT68), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n253), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G179), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n273), .A2(new_n221), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n276), .A2(new_n277), .B1(G20), .B2(G77), .ZN(new_n278));
  XOR2_X1   g0078(.A(KEYINPUT15), .B(G87), .Z(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(new_n222), .A3(G33), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n274), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n250), .A2(G20), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G77), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n283), .A2(new_n285), .B1(G77), .B2(new_n282), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n270), .B2(G169), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n272), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n270), .B2(G190), .ZN(new_n291));
  XOR2_X1   g0091(.A(KEYINPUT69), .B(G200), .Z(new_n292));
  OAI21_X1  g0092(.A(new_n291), .B1(new_n270), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G226), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n248), .B1(new_n294), .B2(new_n252), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n258), .A2(G77), .ZN(new_n296));
  INV_X1    g0096(.A(G222), .ZN(new_n297));
  INV_X1    g0097(.A(G223), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n296), .B1(new_n262), .B2(new_n297), .C1(new_n265), .C2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n271), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n284), .A2(G50), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n283), .A2(new_n303), .B1(G50), .B2(new_n282), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT67), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT67), .ZN(new_n306));
  OAI221_X1 g0106(.A(new_n306), .B1(G50), .B2(new_n282), .C1(new_n283), .C2(new_n303), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n309));
  INV_X1    g0109(.A(G150), .ZN(new_n310));
  INV_X1    g0110(.A(new_n277), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n222), .A2(G33), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n309), .B1(new_n310), .B2(new_n311), .C1(new_n275), .C2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n274), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n302), .B(new_n316), .C1(G169), .C2(new_n301), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n290), .A2(new_n293), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT66), .ZN(new_n319));
  INV_X1    g0119(.A(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n294), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n263), .A2(new_n320), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n264), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G33), .A2(G97), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n247), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n248), .B1(new_n266), .B2(new_n252), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT13), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(G226), .B1(new_n260), .B2(new_n261), .ZN(new_n330));
  INV_X1    g0130(.A(new_n324), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n258), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n326), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n300), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n328), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G190), .ZN(new_n339));
  OR3_X1    g0139(.A1(new_n338), .A2(KEYINPUT71), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT71), .B1(new_n338), .B2(new_n339), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT72), .B1(new_n282), .B2(G68), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT12), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT11), .ZN(new_n345));
  INV_X1    g0145(.A(G50), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n311), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G77), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n312), .A2(new_n348), .B1(new_n222), .B2(G68), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n314), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n344), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n350), .A2(new_n345), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n274), .A2(G68), .A3(new_n282), .A4(new_n284), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(G200), .B2(new_n338), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n342), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(KEYINPUT70), .A2(KEYINPUT10), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n308), .A2(KEYINPUT9), .A3(new_n315), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT9), .B1(new_n308), .B2(new_n315), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT70), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT10), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n301), .A2(new_n292), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n301), .A2(G190), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n358), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n301), .A2(G190), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n369), .B1(new_n363), .B2(new_n364), .C1(new_n292), .C2(new_n301), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT9), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n316), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n359), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n370), .A2(new_n373), .A3(new_n357), .ZN(new_n374));
  NOR4_X1   g0174(.A1(new_n318), .A2(new_n356), .A3(new_n368), .A4(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n248), .B1(new_n263), .B2(new_n252), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n255), .A2(new_n257), .A3(G226), .A4(G1698), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n377), .B(new_n378), .C1(new_n262), .C2(new_n298), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n300), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G200), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(G190), .B2(new_n380), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n264), .B2(G20), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n202), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n277), .A2(G159), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G58), .A2(G68), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT74), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT74), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(G58), .A3(G68), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n390), .A2(new_n392), .A3(new_n203), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n388), .B1(new_n393), .B2(new_n222), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT75), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT16), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT75), .B(new_n397), .C1(new_n387), .C2(new_n394), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n398), .A3(new_n314), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n276), .A2(new_n284), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n400), .A2(new_n283), .B1(new_n282), .B2(new_n276), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n383), .A2(new_n399), .A3(KEYINPUT78), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n274), .B1(new_n395), .B2(KEYINPUT16), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n401), .B1(new_n406), .B2(new_n398), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(KEYINPUT78), .A3(KEYINPUT17), .A4(new_n383), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT77), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n380), .A2(new_n271), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(G169), .B2(new_n380), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n399), .B2(new_n402), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n410), .B1(new_n413), .B2(KEYINPUT18), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  OAI211_X1 g0215(.A(KEYINPUT77), .B(new_n415), .C1(new_n407), .C2(new_n412), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT76), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n413), .B2(KEYINPUT18), .ZN(new_n419));
  NOR4_X1   g0219(.A1(new_n407), .A2(KEYINPUT76), .A3(new_n415), .A4(new_n412), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n409), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n327), .A2(KEYINPUT13), .A3(new_n328), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n336), .B1(new_n334), .B2(new_n335), .ZN(new_n424));
  OAI21_X1  g0224(.A(G169), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n423), .A2(new_n424), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n425), .A2(KEYINPUT14), .B1(new_n426), .B2(G179), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n425), .A2(KEYINPUT73), .A3(KEYINPUT14), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT73), .ZN(new_n429));
  INV_X1    g0229(.A(G169), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n329), .B2(new_n337), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT14), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n427), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n354), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n375), .A2(new_n422), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n255), .A2(new_n257), .A3(new_n222), .A4(G87), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT22), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT22), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n264), .A2(new_n439), .A3(new_n222), .A4(G87), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT24), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G116), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G20), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT23), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n222), .B2(G107), .ZN(new_n446));
  INV_X1    g0246(.A(G107), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(KEYINPUT23), .A3(G20), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n444), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n441), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n442), .B1(new_n441), .B2(new_n449), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n314), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n282), .A2(G107), .ZN(new_n453));
  XOR2_X1   g0253(.A(new_n453), .B(KEYINPUT25), .Z(new_n454));
  INV_X1    g0254(.A(KEYINPUT80), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n250), .A2(G33), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n274), .A2(new_n455), .A3(new_n282), .A4(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n282), .A2(new_n456), .A3(new_n221), .A4(new_n273), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n454), .B1(G107), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n452), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n244), .A2(G1), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  NOR2_X1   g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n466), .A2(G264), .A3(new_n247), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G294), .ZN(new_n468));
  INV_X1    g0268(.A(G257), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(new_n320), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n321), .A2(new_n322), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(G250), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n468), .B1(new_n472), .B2(new_n258), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n467), .B1(new_n473), .B2(new_n300), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(G274), .A3(new_n247), .A4(new_n463), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT86), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(G250), .B1(new_n260), .B2(new_n261), .ZN(new_n478));
  INV_X1    g0278(.A(new_n470), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n258), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n468), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n300), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n467), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT86), .A4(new_n476), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n339), .B1(new_n477), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n482), .A2(new_n483), .A3(new_n476), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n381), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n462), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT86), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(G169), .A3(new_n484), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n474), .A2(G179), .A3(new_n476), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n492), .A2(new_n493), .B1(new_n452), .B2(new_n461), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT85), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n466), .A2(G270), .A3(new_n247), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(G179), .A3(new_n476), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT84), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n469), .B1(new_n321), .B2(new_n322), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G264), .A2(G1698), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n255), .A2(new_n257), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n300), .B1(new_n264), .B2(G303), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n499), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(G257), .B1(new_n260), .B2(new_n261), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(new_n264), .A3(new_n501), .ZN(new_n507));
  INV_X1    g0307(.A(G303), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n247), .B1(new_n258), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT84), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n498), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G116), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n458), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n282), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n512), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n273), .A2(new_n221), .B1(G20), .B2(new_n512), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G283), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n517), .B(new_n222), .C1(G33), .C2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(KEYINPUT20), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT20), .B1(new_n516), .B2(new_n519), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n513), .B(new_n515), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n496), .B1(new_n511), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n511), .A2(new_n496), .A3(new_n523), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n505), .A2(new_n510), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n497), .A2(new_n476), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n522), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n520), .ZN(new_n533));
  MUX2_X1   g0333(.A(new_n282), .B(new_n458), .S(G116), .Z(new_n534));
  AOI21_X1  g0334(.A(new_n430), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(new_n535), .A3(KEYINPUT21), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n529), .B1(new_n505), .B2(new_n510), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G190), .ZN(new_n538));
  INV_X1    g0338(.A(new_n523), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n538), .B(new_n539), .C1(new_n381), .C2(new_n537), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n523), .A2(G169), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(new_n537), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n527), .A2(new_n536), .A3(new_n540), .A4(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT7), .B1(new_n258), .B2(new_n222), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n384), .B(G20), .C1(new_n255), .C2(new_n257), .ZN(new_n546));
  OAI21_X1  g0346(.A(G107), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n311), .A2(new_n348), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT6), .ZN(new_n549));
  AND2_X1   g0349(.A1(G97), .A2(G107), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT79), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n553), .A2(new_n447), .A3(KEYINPUT6), .A4(G97), .ZN(new_n554));
  NAND2_X1  g0354(.A1(KEYINPUT6), .A2(G97), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT79), .B1(new_n555), .B2(G107), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n548), .B1(new_n557), .B2(G20), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n547), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n314), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n562));
  OAI21_X1  g0362(.A(G97), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n514), .A2(G97), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT81), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n518), .B1(new_n457), .B2(new_n459), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT81), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n567), .A2(new_n568), .A3(new_n564), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n560), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n262), .B2(new_n249), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n471), .A2(new_n264), .A3(KEYINPUT4), .A4(G244), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n255), .A2(new_n257), .A3(G250), .A4(G1698), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n572), .A2(new_n517), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n300), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n466), .A2(new_n247), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n476), .B1(new_n577), .B2(new_n469), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n430), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n576), .A2(new_n271), .A3(new_n579), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n570), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n274), .B1(new_n547), .B2(new_n558), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n563), .A2(KEYINPUT81), .A3(new_n565), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n568), .B1(new_n567), .B2(new_n564), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n574), .A2(new_n517), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n262), .A2(new_n249), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(KEYINPUT4), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n247), .B1(new_n590), .B2(new_n572), .ZN(new_n591));
  OAI21_X1  g0391(.A(G200), .B1(new_n591), .B2(new_n578), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n576), .A2(G190), .A3(new_n579), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n587), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n583), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n279), .A2(new_n282), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT19), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n222), .B1(new_n326), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(G87), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n551), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n255), .A2(new_n257), .A3(new_n222), .A4(G68), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n597), .B1(new_n312), .B2(new_n518), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n596), .B1(new_n604), .B2(new_n314), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n457), .A2(new_n459), .A3(new_n279), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n605), .A2(KEYINPUT83), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT83), .B1(new_n605), .B2(new_n606), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n250), .A2(G45), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n610), .A2(G250), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n247), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n247), .A2(G274), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(new_n610), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT82), .B1(new_n262), .B2(new_n266), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT82), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n471), .A2(new_n264), .A3(new_n616), .A4(G238), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n255), .A2(new_n257), .A3(G244), .A4(G1698), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n615), .A2(new_n443), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n614), .B1(new_n619), .B2(new_n300), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n271), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n443), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n471), .A2(new_n264), .A3(G238), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(KEYINPUT82), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n247), .B1(new_n624), .B2(new_n617), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n430), .B1(new_n625), .B2(new_n614), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n609), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n460), .A2(G87), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n628), .A2(new_n605), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n619), .A2(new_n300), .ZN(new_n630));
  INV_X1    g0430(.A(new_n614), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G190), .A3(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n629), .B(new_n632), .C1(new_n292), .C2(new_n620), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n544), .A2(new_n595), .A3(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n436), .A2(new_n495), .A3(new_n635), .ZN(G372));
  INV_X1    g0436(.A(new_n317), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n413), .B(new_n415), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n356), .A2(new_n290), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(new_n354), .B2(new_n434), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n639), .B1(new_n641), .B2(new_n409), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT90), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n374), .B2(new_n368), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n357), .B1(new_n370), .B2(new_n373), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n362), .A2(new_n367), .A3(new_n358), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT90), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n637), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n595), .A2(new_n489), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT88), .B1(new_n620), .B2(new_n292), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT88), .ZN(new_n652));
  INV_X1    g0452(.A(new_n292), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n652), .B(new_n653), .C1(new_n625), .C2(new_n614), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n651), .A2(new_n654), .A3(new_n629), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT89), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT89), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n651), .A2(new_n654), .A3(new_n657), .A4(new_n629), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n632), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n626), .A2(KEYINPUT87), .ZN(new_n660));
  OR3_X1    g0460(.A1(new_n620), .A2(KEYINPUT87), .A3(G169), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n620), .A2(new_n271), .B1(new_n605), .B2(new_n606), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n511), .A2(new_n496), .A3(new_n523), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n536), .B(new_n543), .C1(new_n664), .C2(new_n524), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n492), .A2(new_n493), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n462), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n650), .A2(new_n659), .A3(new_n663), .A4(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  INV_X1    g0471(.A(new_n583), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n659), .A2(new_n671), .A3(new_n672), .A4(new_n663), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT26), .B1(new_n634), .B2(new_n583), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n670), .A2(new_n673), .A3(new_n663), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n436), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n649), .A2(new_n676), .ZN(G369));
  INV_X1    g0477(.A(new_n495), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n250), .A2(new_n222), .A3(G13), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n452), .B2(new_n461), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n678), .A2(new_n686), .B1(new_n668), .B2(new_n685), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n539), .A2(new_n685), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n665), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n544), .B2(new_n688), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n494), .A2(new_n685), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n665), .A2(new_n685), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n495), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n692), .A2(new_n693), .A3(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n216), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n600), .A2(G116), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n219), .B2(new_n700), .ZN(new_n703));
  XOR2_X1   g0503(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n704));
  XNOR2_X1  g0504(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n672), .A2(new_n671), .A3(new_n633), .A4(new_n627), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n670), .A2(new_n663), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n663), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n655), .A2(KEYINPUT89), .B1(G190), .B2(new_n620), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n658), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n671), .B1(new_n710), .B2(new_n672), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n685), .B1(new_n707), .B2(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n675), .A2(new_n685), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n630), .A2(new_n474), .A3(new_n631), .ZN(new_n717));
  INV_X1    g0517(.A(new_n498), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n528), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT92), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n591), .A2(new_n578), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n511), .A2(KEYINPUT92), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n717), .A2(new_n721), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI211_X1 g0526(.A(new_n725), .B(new_n578), .C1(new_n575), .C2(new_n300), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n717), .A2(new_n721), .A3(new_n723), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n537), .A2(G179), .ZN(new_n729));
  INV_X1    g0529(.A(new_n620), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n729), .A2(new_n730), .A3(new_n487), .A4(new_n580), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT31), .B(new_n684), .C1(new_n726), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT93), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n728), .A2(new_n731), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n724), .A2(new_n725), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n685), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT94), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n738), .A2(new_n739), .A3(KEYINPUT31), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n684), .B1(new_n726), .B2(new_n732), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT94), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n735), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  AND4_X1   g0544(.A1(new_n583), .A2(new_n627), .A3(new_n594), .A4(new_n633), .ZN(new_n745));
  INV_X1    g0545(.A(new_n540), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n665), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n495), .A2(new_n745), .A3(new_n747), .A4(new_n685), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT95), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT95), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n635), .A2(new_n750), .A3(new_n495), .A4(new_n685), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n739), .B1(new_n738), .B2(KEYINPUT31), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n741), .A2(KEYINPUT94), .A3(new_n742), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n753), .A2(new_n754), .A3(new_n734), .A4(new_n733), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n744), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n716), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT96), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n705), .B1(new_n760), .B2(G1), .ZN(G364));
  INV_X1    g0561(.A(G13), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n250), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n699), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n264), .A2(G355), .A3(new_n216), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G116), .B2(new_n216), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n238), .A2(G45), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n698), .A2(new_n264), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n244), .B2(new_n220), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n768), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n222), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT98), .Z(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n221), .B1(G20), .B2(new_n430), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n766), .B1(new_n773), .B2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n339), .A2(G179), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n222), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n518), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n222), .A2(G179), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G190), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G159), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n784), .B1(KEYINPUT32), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(KEYINPUT32), .B2(new_n789), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n222), .A2(new_n271), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT100), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT100), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n791), .B1(G50), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n792), .A2(new_n786), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n792), .A2(new_n339), .A3(G200), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n264), .B1(new_n798), .B2(new_n348), .C1(new_n202), .C2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n653), .A2(G190), .A3(new_n785), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n599), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n653), .A2(new_n339), .A3(new_n785), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n800), .B(new_n802), .C1(G107), .C2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n792), .A2(G190), .A3(new_n381), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT99), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n797), .B(new_n805), .C1(new_n201), .C2(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G322), .A2(new_n810), .B1(new_n796), .B2(G326), .ZN(new_n813));
  INV_X1    g0613(.A(new_n801), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G283), .A2(new_n804), .B1(new_n814), .B2(G303), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n258), .B1(new_n798), .B2(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(KEYINPUT33), .B(G317), .Z(new_n818));
  INV_X1    g0618(.A(G329), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n799), .A2(new_n818), .B1(new_n819), .B2(new_n787), .ZN(new_n820));
  INV_X1    g0620(.A(new_n783), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n817), .B(new_n820), .C1(G294), .C2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n813), .A2(new_n815), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n812), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n781), .B1(new_n824), .B2(new_n778), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n690), .B2(new_n776), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n690), .A2(G330), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT97), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n691), .A2(new_n766), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT101), .Z(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  NAND2_X1  g0632(.A1(new_n288), .A2(new_n684), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n293), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n290), .ZN(new_n835));
  OR3_X1    g0635(.A1(new_n272), .A2(new_n289), .A3(new_n684), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n714), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n835), .A2(new_n836), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n675), .A2(new_n685), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n766), .B1(new_n757), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n757), .B2(new_n841), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n258), .B1(new_n788), .B2(G132), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n844), .B1(new_n201), .B2(new_n783), .C1(new_n803), .C2(new_n202), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n810), .A2(G143), .ZN(new_n846));
  INV_X1    g0646(.A(new_n799), .ZN(new_n847));
  INV_X1    g0647(.A(new_n798), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n847), .A2(G150), .B1(new_n848), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(new_n796), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n846), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT34), .Z(new_n853));
  AOI211_X1 g0653(.A(new_n845), .B(new_n853), .C1(G50), .C2(new_n814), .ZN(new_n854));
  INV_X1    g0654(.A(G294), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n811), .A2(new_n855), .B1(new_n850), .B2(new_n508), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n599), .A2(new_n803), .B1(new_n801), .B2(new_n447), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G116), .A2(new_n848), .B1(new_n788), .B2(G311), .ZN(new_n858));
  INV_X1    g0658(.A(G283), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n858), .B(new_n258), .C1(new_n859), .C2(new_n799), .ZN(new_n860));
  NOR4_X1   g0660(.A1(new_n856), .A2(new_n857), .A3(new_n784), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n778), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n837), .A2(new_n774), .ZN(new_n863));
  INV_X1    g0663(.A(new_n766), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n778), .A2(new_n774), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n864), .B1(new_n348), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n862), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n843), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(G384));
  NOR2_X1   g0669(.A1(new_n763), .A2(new_n250), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n733), .A2(KEYINPUT104), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n741), .A2(new_n742), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n741), .A2(KEYINPUT104), .A3(new_n742), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n752), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT103), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n329), .A2(G179), .A3(new_n337), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n431), .B2(new_n432), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT73), .B1(new_n425), .B2(KEYINPUT14), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n431), .A2(new_n429), .A3(new_n432), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n354), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n876), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n434), .A2(KEYINPUT103), .A3(new_n354), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n882), .A2(new_n685), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n342), .B2(new_n355), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(new_n356), .B2(new_n434), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n837), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n399), .A2(new_n402), .ZN(new_n890));
  INV_X1    g0690(.A(new_n682), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n412), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(KEYINPUT18), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT76), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n413), .A2(new_n418), .A3(KEYINPUT18), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n895), .A2(new_n414), .A3(new_n416), .A4(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n409), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n892), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n890), .A2(new_n893), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n407), .A2(new_n383), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n892), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n900), .A2(new_n892), .A3(new_n904), .A4(new_n901), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n899), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n892), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n638), .B2(new_n409), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n903), .A2(new_n905), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n875), .B(new_n889), .C1(new_n908), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n887), .A2(new_n888), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n839), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT104), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n738), .A2(new_n916), .A3(KEYINPUT31), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n872), .B2(new_n871), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n915), .B1(new_n752), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(KEYINPUT38), .B(new_n911), .C1(new_n422), .C2(new_n892), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n907), .B1(new_n899), .B2(new_n906), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT40), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n913), .A2(KEYINPUT40), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT105), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n436), .A2(new_n875), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(G330), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n436), .B1(new_n713), .B2(new_n715), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n649), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n908), .B2(new_n912), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n883), .A2(new_n884), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n933), .A2(new_n684), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT39), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n914), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n840), .B2(new_n836), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n920), .A2(new_n921), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n638), .A2(new_n682), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n936), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n930), .B(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n870), .B1(new_n928), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n928), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n557), .A2(KEYINPUT35), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n557), .A2(KEYINPUT35), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n946), .A2(G116), .A3(new_n223), .A4(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT36), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n220), .A2(G77), .A3(new_n392), .A4(new_n390), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n951), .A2(KEYINPUT102), .B1(new_n346), .B2(G68), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(KEYINPUT102), .B2(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(G1), .A3(new_n762), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n945), .A2(new_n949), .A3(new_n954), .ZN(G367));
  NAND2_X1  g0755(.A1(new_n672), .A2(new_n684), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n583), .B(new_n594), .C1(new_n587), .C2(new_n685), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(new_n495), .A3(new_n695), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(KEYINPUT42), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n959), .A2(KEYINPUT42), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n583), .B1(new_n957), .B2(new_n668), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n960), .B(new_n961), .C1(new_n685), .C2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n629), .A2(new_n685), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n663), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n710), .B2(new_n964), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT106), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n963), .B1(KEYINPUT43), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n958), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n692), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n970), .B(new_n972), .Z(new_n973));
  XNOR2_X1  g0773(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n699), .B(new_n974), .Z(new_n975));
  INV_X1    g0775(.A(KEYINPUT110), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n758), .B(KEYINPUT96), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT109), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n696), .B1(new_n691), .B2(new_n978), .C1(new_n687), .C2(new_n695), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n691), .A2(new_n978), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n976), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n981), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n760), .A2(KEYINPUT110), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n696), .A2(new_n693), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT108), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n985), .A2(new_n971), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n986), .A2(KEYINPUT108), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n988), .B(new_n989), .Z(new_n990));
  NOR2_X1   g0790(.A1(new_n985), .A2(new_n971), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(new_n692), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n982), .A2(new_n984), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n975), .B1(new_n995), .B2(new_n760), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n973), .B1(new_n996), .B2(new_n765), .ZN(new_n997));
  INV_X1    g0797(.A(new_n279), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n779), .B1(new_n216), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n233), .A2(new_n771), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n766), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n847), .A2(G159), .B1(new_n788), .B2(G137), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1002), .B(new_n264), .C1(new_n346), .C2(new_n798), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G68), .B2(new_n821), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G58), .A2(new_n814), .B1(new_n804), .B2(G77), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G150), .A2(new_n810), .B1(new_n796), .B2(G143), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n814), .A2(G116), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT46), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n508), .B2(new_n811), .C1(new_n816), .C2(new_n850), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n804), .A2(G97), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n821), .A2(G107), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n264), .B1(new_n788), .B2(G317), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n847), .A2(G294), .B1(new_n848), .B2(G283), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1007), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n1017));
  XNOR2_X1  g0817(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1001), .B1(new_n1018), .B2(new_n778), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n967), .B2(new_n776), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n997), .A2(new_n1020), .ZN(G387));
  NAND2_X1  g0821(.A1(new_n982), .A2(new_n984), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n699), .B1(new_n760), .B2(new_n983), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G50), .A2(new_n810), .B1(new_n796), .B2(G159), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n998), .A2(new_n783), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n799), .A2(new_n275), .B1(new_n798), .B2(new_n202), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n264), .B1(new_n787), .B2(new_n310), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n814), .A2(G77), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1026), .A2(new_n1011), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n264), .B1(new_n788), .B2(G326), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n796), .A2(G322), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n816), .B2(new_n799), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT113), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(KEYINPUT113), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n810), .A2(G317), .B1(G303), .B2(new_n848), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT48), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n814), .A2(G294), .B1(G283), .B2(new_n821), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1033), .B1(new_n512), .B2(new_n803), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1032), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT114), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n778), .A3(new_n1051), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n687), .A2(new_n776), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n701), .A2(new_n258), .A3(new_n698), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n447), .B2(new_n698), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT112), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n230), .A2(new_n244), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n276), .A2(new_n346), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT50), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n701), .B(new_n244), .C1(new_n202), .C2(new_n348), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n770), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1056), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n864), .B1(new_n1062), .B2(new_n779), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n1052), .A2(new_n1053), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n765), .B2(new_n983), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1025), .A2(new_n1065), .ZN(G393));
  NAND2_X1  g0866(.A1(new_n994), .A2(new_n765), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n958), .A2(new_n776), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT115), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n779), .B1(new_n518), .B2(new_n216), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n241), .A2(new_n770), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n766), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G311), .A2(new_n810), .B1(new_n796), .B2(G317), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT52), .Z(new_n1074));
  AOI22_X1  g0874(.A1(new_n847), .A2(G303), .B1(new_n788), .B2(G322), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n258), .C1(new_n855), .C2(new_n798), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G116), .B2(new_n821), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G107), .A2(new_n804), .B1(new_n814), .B2(G283), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1074), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G159), .A2(new_n810), .B1(new_n796), .B2(G150), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT51), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n847), .A2(G50), .B1(new_n788), .B2(G143), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n258), .B1(new_n848), .B2(new_n276), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(new_n348), .C2(new_n783), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n202), .A2(new_n801), .B1(new_n803), .B2(new_n599), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1079), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1072), .B1(new_n1087), .B2(new_n778), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1069), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n995), .A2(new_n699), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n994), .B1(new_n982), .B2(new_n984), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1067), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(G390));
  AND3_X1   g0892(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT39), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n912), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT39), .B1(new_n1094), .B2(new_n920), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n774), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n802), .B1(G68), .B2(new_n804), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G116), .A2(new_n810), .B1(new_n796), .B2(G283), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n258), .B1(new_n798), .B2(new_n518), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n799), .A2(new_n447), .B1(new_n787), .B2(new_n855), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(G77), .C2(new_n821), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1097), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G132), .A2(new_n810), .B1(new_n796), .B2(G128), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT54), .B(G143), .ZN(new_n1104));
  INV_X1    g0904(.A(G125), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n798), .A2(new_n1104), .B1(new_n787), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n264), .B1(new_n799), .B2(new_n851), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G159), .C2(new_n821), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1103), .B(new_n1108), .C1(new_n346), .C2(new_n803), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n801), .A2(new_n310), .ZN(new_n1110));
  XOR2_X1   g0910(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1111));
  XNOR2_X1  g0911(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1102), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n778), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n864), .B1(new_n275), .B2(new_n865), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1096), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(G330), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n918), .B2(new_n752), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n889), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n840), .A2(new_n836), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n914), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n934), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1122), .A2(new_n1123), .B1(new_n932), .B2(new_n935), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n908), .B2(new_n912), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n685), .B(new_n835), .C1(new_n707), .C2(new_n711), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n836), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1125), .B1(new_n914), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1120), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n1093), .A2(new_n1095), .B1(new_n938), .B2(new_n934), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1125), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1127), .A2(new_n914), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n756), .A2(G330), .A3(new_n839), .A4(new_n914), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1130), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1116), .B1(new_n1136), .B2(new_n764), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1118), .A2(new_n436), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n929), .A2(new_n649), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n756), .A2(G330), .A3(new_n839), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1140), .A2(new_n937), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1121), .B1(new_n1141), .B2(new_n1120), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n875), .A2(G330), .A3(new_n839), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n937), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1127), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n1134), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1139), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1130), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1119), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1150), .A3(KEYINPUT116), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1140), .A2(new_n937), .B1(new_n889), .B2(new_n1118), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1121), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1146), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n929), .A2(new_n1138), .A3(new_n649), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1154), .A2(new_n1129), .A3(new_n1135), .A4(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT116), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1151), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n700), .B1(new_n1160), .B2(new_n1136), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1137), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(G378));
  NAND3_X1  g0963(.A1(new_n644), .A2(new_n317), .A3(new_n647), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n316), .A2(new_n891), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n644), .A2(new_n317), .A3(new_n647), .A4(new_n1165), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n774), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n243), .B(new_n258), .C1(new_n799), .C2(new_n518), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n998), .A2(new_n798), .B1(new_n859), .B2(new_n787), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(G68), .C2(new_n821), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n804), .A2(G58), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G107), .A2(new_n810), .B1(new_n796), .B2(G116), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1176), .A2(new_n1031), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT58), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G50), .B1(new_n254), .B2(new_n243), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n264), .B2(G41), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n847), .A2(G132), .B1(new_n848), .B2(G137), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n310), .B2(new_n783), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1104), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n814), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(G128), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1186), .B1(new_n1105), .B2(new_n850), .C1(new_n1187), .C2(new_n811), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n804), .A2(G159), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G33), .B(G41), .C1(new_n788), .C2(G124), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1180), .B(new_n1182), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT118), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n778), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n864), .B1(new_n346), .B2(new_n865), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1173), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT119), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1172), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n749), .A2(new_n751), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n916), .B1(new_n738), .B2(KEYINPUT31), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n738), .A2(KEYINPUT31), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n874), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n889), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n897), .A2(new_n898), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1209), .A2(new_n909), .B1(new_n903), .B2(new_n905), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n912), .B1(new_n1210), .B2(KEYINPUT38), .ZN(new_n1211));
  OAI21_X1  g1011(.A(KEYINPUT40), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT40), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n939), .A2(new_n1213), .A3(new_n875), .A4(new_n889), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1203), .B1(new_n1215), .B2(G330), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1117), .B(new_n1172), .C1(new_n1212), .C2(new_n1214), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1216), .A2(new_n1217), .A3(new_n942), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n942), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1172), .B1(new_n923), .B2(new_n1117), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1215), .A2(G330), .A3(new_n1203), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1202), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n942), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1220), .A2(new_n1219), .A3(new_n1221), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(KEYINPUT119), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1201), .B1(new_n1227), .B2(new_n765), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT116), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1155), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1227), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1139), .B1(new_n1151), .B2(new_n1158), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT120), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1224), .A2(new_n1234), .A3(new_n1225), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1220), .A2(new_n1221), .A3(new_n1219), .A4(KEYINPUT120), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(KEYINPUT57), .A3(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n699), .B1(new_n1233), .B2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1228), .B1(new_n1232), .B2(new_n1238), .ZN(G375));
  NAND3_X1  g1039(.A1(new_n1142), .A2(new_n1139), .A3(new_n1146), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT121), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1240), .B(new_n1241), .ZN(new_n1242));
  OR3_X1    g1042(.A1(new_n1242), .A2(new_n975), .A3(new_n1147), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1154), .A2(new_n765), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n937), .A2(new_n774), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT122), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G107), .A2(new_n848), .B1(new_n788), .B2(G303), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1247), .B(new_n258), .C1(new_n512), .C2(new_n799), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n348), .A2(new_n803), .B1(new_n801), .B2(new_n518), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1248), .A2(new_n1249), .A3(new_n1027), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1250), .B1(new_n859), .B2(new_n811), .C1(new_n855), .C2(new_n850), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G137), .A2(new_n810), .B1(new_n796), .B2(G132), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n798), .A2(new_n310), .B1(new_n787), .B2(new_n1187), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n264), .B1(new_n799), .B2(new_n1104), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(G50), .C2(new_n821), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n814), .A2(G159), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1252), .A2(new_n1255), .A3(new_n1177), .A4(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1251), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n778), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n864), .B1(new_n202), .B2(new_n865), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1246), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1244), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1243), .A2(new_n1263), .ZN(G381));
  NAND3_X1  g1064(.A1(new_n1025), .A2(new_n831), .A3(new_n1065), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(G384), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT123), .ZN(new_n1267));
  INV_X1    g1067(.A(G390), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1268), .A2(new_n1162), .A3(new_n1263), .A4(new_n1243), .ZN(new_n1269));
  OR4_X1    g1069(.A1(G387), .A2(new_n1267), .A3(G375), .A4(new_n1269), .ZN(G407));
  NAND2_X1  g1070(.A1(new_n683), .A2(G213), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1162), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G407), .B(G213), .C1(G375), .C2(new_n1273), .ZN(G409));
  NAND2_X1  g1074(.A1(new_n1272), .A2(G2897), .ZN(new_n1275));
  XOR2_X1   g1075(.A(new_n1275), .B(KEYINPUT125), .Z(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1240), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n700), .B1(new_n1278), .B2(KEYINPUT60), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1160), .A2(KEYINPUT60), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1242), .B2(new_n1280), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1281), .A2(G384), .A3(new_n1263), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G384), .B1(new_n1281), .B2(new_n1263), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1277), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1263), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n868), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1281), .A2(G384), .A3(new_n1263), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1276), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1284), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1235), .A2(new_n765), .A3(new_n1236), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1200), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT124), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n975), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1231), .A2(new_n1294), .A3(new_n1227), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT124), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1291), .A2(new_n1296), .A3(new_n1200), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1293), .A2(new_n1295), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1162), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G378), .B(new_n1228), .C1(new_n1232), .C2(new_n1238), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1271), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT61), .B1(new_n1290), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1304), .B1(new_n1302), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G390), .B1(new_n997), .B2(new_n1020), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n831), .B1(new_n1025), .B2(new_n1065), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1311), .A2(KEYINPUT126), .A3(new_n1265), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT126), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1025), .A2(new_n831), .A3(new_n1065), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1313), .B1(new_n1314), .B2(new_n1310), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1312), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n997), .A2(new_n1020), .A3(G390), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1309), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1317), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1315), .B1(new_n1319), .B2(new_n1308), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1272), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(KEYINPUT63), .A3(new_n1305), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1303), .A2(new_n1307), .A3(new_n1321), .A4(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT62), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1322), .A2(new_n1325), .A3(new_n1305), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT61), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1327), .B1(new_n1322), .B2(new_n1289), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1325), .B1(new_n1322), .B2(new_n1305), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1326), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1324), .B1(new_n1330), .B2(new_n1321), .ZN(G405));
  NAND2_X1  g1131(.A1(G375), .A2(new_n1162), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1300), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1333), .B(new_n1306), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1334), .B(new_n1321), .ZN(G402));
endmodule


