//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956;
  INV_X1    g000(.A(KEYINPUT1), .ZN(new_n202));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT68), .B(G120gat), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n205), .A2(G120gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n202), .B(new_n203), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n209));
  OR2_X1    g008(.A1(G127gat), .A2(G134gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211));
  NAND2_X1  g010(.A1(G127gat), .A2(G134gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n205), .A2(G120gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n202), .B1(new_n207), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n215), .B1(new_n214), .B2(new_n217), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n208), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G141gat), .B(G148gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(G155gat), .B(G162gat), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(KEYINPUT74), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(KEYINPUT74), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  INV_X1    g026(.A(G162gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT2), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n222), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n223), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n221), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n217), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT67), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n218), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n233), .B1(new_n226), .B2(new_n229), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(new_n208), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G225gat), .A2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT75), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(KEYINPUT5), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n243), .B1(new_n236), .B2(new_n241), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT5), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT75), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n241), .A2(KEYINPUT4), .ZN(new_n251));
  INV_X1    g050(.A(new_n208), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(new_n238), .B2(new_n218), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n240), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n259), .A3(new_n221), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(new_n243), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n247), .A2(new_n250), .A3(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n260), .A2(new_n249), .A3(new_n243), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n256), .A2(KEYINPUT76), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT76), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n251), .A2(new_n265), .A3(new_n255), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268));
  INV_X1    g067(.A(G85gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT0), .B(G57gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n262), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n273), .B1(new_n262), .B2(new_n267), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI211_X1 g077(.A(new_n275), .B(new_n273), .C1(new_n262), .C2(new_n267), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT82), .ZN(new_n281));
  XNOR2_X1  g080(.A(G197gat), .B(G204gat), .ZN(new_n282));
  AND2_X1   g081(.A1(G211gat), .A2(G218gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(KEYINPUT22), .B2(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(G211gat), .B(G218gat), .Z(new_n285));
  OR2_X1    g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n285), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n292));
  NOR2_X1   g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT23), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT25), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301));
  INV_X1    g100(.A(G183gat), .ZN(new_n302));
  INV_X1    g101(.A(G190gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n304), .B(new_n305), .C1(G183gat), .C2(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n298), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n298), .B(new_n306), .C1(new_n299), .C2(KEYINPUT25), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT27), .B(G183gat), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT65), .B1(new_n311), .B2(new_n303), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n312), .A2(KEYINPUT28), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n293), .A2(KEYINPUT26), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n297), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n293), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(KEYINPUT28), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n313), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n292), .B1(new_n310), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n310), .A2(new_n318), .A3(new_n292), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(KEYINPUT70), .B(KEYINPUT29), .Z(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n291), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n318), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n291), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT71), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n329), .A3(new_n291), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n289), .B1(new_n325), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n321), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n291), .B1(new_n333), .B2(new_n319), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n291), .B1(new_n326), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n322), .A2(KEYINPUT72), .A3(new_n291), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n288), .ZN(new_n340));
  XOR2_X1   g139(.A(G64gat), .B(G92gat), .Z(new_n341));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n332), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT37), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n332), .A2(new_n340), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n288), .B1(new_n325), .B2(new_n331), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n338), .A2(new_n339), .A3(new_n289), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT37), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT38), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n343), .B(KEYINPUT73), .Z(new_n351));
  NAND4_X1  g150(.A1(new_n346), .A2(new_n349), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n280), .A2(new_n281), .A3(new_n344), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n332), .A2(new_n340), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n343), .B1(new_n354), .B2(KEYINPUT37), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n355), .A2(KEYINPUT83), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n346), .B1(new_n355), .B2(KEYINPUT83), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT38), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n262), .A2(new_n267), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n272), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n275), .A3(new_n274), .ZN(new_n361));
  INV_X1    g160(.A(new_n279), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n361), .A2(new_n352), .A3(new_n362), .A4(new_n344), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT82), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n353), .A2(new_n358), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n288), .B1(new_n259), .B2(new_n324), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n288), .A2(KEYINPUT79), .A3(new_n336), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n258), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT79), .B1(new_n288), .B2(new_n336), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n235), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n367), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n240), .B1(KEYINPUT77), .B2(new_n289), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n287), .A2(KEYINPUT77), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n324), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n377), .A2(new_n378), .A3(new_n257), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n377), .B2(new_n257), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n379), .A2(new_n380), .A3(new_n366), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n374), .B1(new_n381), .B2(new_n373), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G22gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n384));
  INV_X1    g183(.A(G22gat), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n385), .B(new_n374), .C1(new_n381), .C2(new_n373), .ZN(new_n386));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT31), .B(G50gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n383), .A2(new_n384), .A3(new_n386), .A4(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(KEYINPUT80), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n392), .A2(new_n389), .B1(new_n383), .B2(new_n386), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT30), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n344), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n354), .A2(new_n351), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT30), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n399), .B2(new_n344), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n264), .A2(new_n260), .A3(new_n266), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n244), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n236), .A2(new_n241), .A3(new_n243), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n404), .A2(KEYINPUT81), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(KEYINPUT81), .ZN(new_n406));
  AND4_X1   g205(.A1(KEYINPUT39), .A2(new_n403), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT40), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n273), .B1(new_n403), .B2(KEYINPUT39), .ZN(new_n409));
  OR3_X1    g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n407), .B2(new_n409), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n401), .A2(new_n360), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n365), .A2(new_n395), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n326), .A2(new_n221), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n253), .A2(new_n310), .A3(new_n318), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G227gat), .ZN(new_n417));
  INV_X1    g216(.A(G233gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT32), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT33), .B1(new_n416), .B2(new_n419), .ZN(new_n423));
  XNOR2_X1  g222(.A(G15gat), .B(G43gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(G71gat), .B(G99gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT34), .B1(new_n416), .B2(new_n419), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT34), .ZN(new_n429));
  INV_X1    g228(.A(new_n419), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n428), .B(new_n431), .C1(new_n423), .C2(new_n426), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n422), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n422), .A3(new_n434), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT36), .ZN(new_n439));
  INV_X1    g238(.A(new_n280), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n400), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n439), .B1(new_n441), .B2(new_n394), .ZN(new_n442));
  INV_X1    g241(.A(new_n438), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n391), .B2(new_n393), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT35), .B1(new_n444), .B2(new_n441), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n392), .A2(new_n389), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n383), .A2(new_n386), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n438), .B1(new_n448), .B2(new_n390), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT35), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n440), .A4(new_n400), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n413), .A2(new_n442), .B1(new_n445), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G231gat), .A2(G233gat), .ZN(new_n453));
  INV_X1    g252(.A(G211gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G8gat), .ZN(new_n456));
  OR2_X1    g255(.A1(G15gat), .A2(G22gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(G15gat), .A2(G22gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT87), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(G1gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(KEYINPUT87), .A3(new_n458), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n461), .A2(new_n463), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT16), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT88), .B1(new_n466), .B2(G1gat), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(new_n462), .A3(KEYINPUT16), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n456), .B(new_n464), .C1(new_n465), .C2(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n461), .B2(new_n463), .ZN(new_n473));
  OAI21_X1  g272(.A(G8gat), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(G71gat), .B(G78gat), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G64gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G57gat), .ZN(new_n480));
  INV_X1    g279(.A(G57gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G64gat), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n480), .A2(new_n482), .A3(KEYINPUT91), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT91), .B1(new_n480), .B2(new_n482), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n478), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n486), .B(KEYINPUT92), .ZN(new_n490));
  INV_X1    g289(.A(new_n480), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT93), .B(G57gat), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(G64gat), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n490), .A2(new_n493), .A3(new_n477), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT21), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n476), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G183gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n476), .A2(new_n496), .A3(new_n302), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n500), .B1(new_n498), .B2(new_n499), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n455), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n503), .ZN(new_n505));
  INV_X1    g304(.A(new_n455), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n495), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(G127gat), .B(G155gat), .Z(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n504), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n504), .B2(new_n507), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G50gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G43gat), .ZN(new_n516));
  INV_X1    g315(.A(G43gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G50gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n518), .A3(KEYINPUT15), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  INV_X1    g319(.A(G36gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT14), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n520), .A3(new_n521), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n519), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT85), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n530), .B1(new_n525), .B2(new_n526), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n525), .A2(new_n530), .A3(new_n526), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n518), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT15), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(new_n523), .A3(new_n519), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n534), .A2(new_n538), .A3(KEYINPUT86), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT86), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n516), .A2(new_n518), .A3(KEYINPUT15), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT15), .B1(new_n516), .B2(new_n518), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n541), .A2(new_n542), .A3(new_n522), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n525), .A2(new_n530), .A3(new_n526), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(new_n531), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n540), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n529), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT17), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT86), .B1(new_n534), .B2(new_n538), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n543), .A2(new_n545), .A3(new_n540), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n552), .A3(new_n529), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(G92gat), .ZN(new_n556));
  INV_X1    g355(.A(G92gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(KEYINPUT97), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n269), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G85gat), .A2(G92gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(KEYINPUT96), .A3(KEYINPUT7), .ZN(new_n561));
  NAND2_X1  g360(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(G85gat), .A3(G92gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT8), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(G99gat), .B2(G106gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n559), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT98), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n572), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT98), .B1(new_n574), .B2(new_n569), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n568), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n557), .A2(KEYINPUT97), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n555), .A2(G92gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n566), .B1(new_n580), .B2(new_n269), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n581), .A2(new_n564), .B1(new_n575), .B2(new_n573), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n554), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT99), .ZN(new_n586));
  XOR2_X1   g385(.A(G190gat), .B(G218gat), .Z(new_n587));
  AND2_X1   g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n547), .A2(new_n583), .B1(KEYINPUT41), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n554), .A2(new_n590), .A3(new_n584), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n586), .A2(new_n587), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n592), .A2(KEYINPUT100), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n588), .A2(KEYINPUT41), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(new_n228), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT95), .B(G134gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n586), .A2(new_n589), .A3(new_n591), .ZN(new_n598));
  INV_X1    g397(.A(new_n587), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n593), .A2(new_n597), .B1(new_n600), .B2(new_n592), .ZN(new_n601));
  AND4_X1   g400(.A1(KEYINPUT100), .A2(new_n600), .A3(new_n592), .A4(new_n597), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n551), .A2(new_n529), .B1(new_n474), .B2(new_n471), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n554), .B2(new_n476), .ZN(new_n605));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT18), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT89), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n552), .B1(new_n551), .B2(new_n529), .ZN(new_n610));
  AOI211_X1 g409(.A(KEYINPUT17), .B(new_n528), .C1(new_n549), .C2(new_n550), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n476), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n547), .A2(new_n475), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n612), .A2(KEYINPUT18), .A3(new_n606), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n606), .B(KEYINPUT13), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n547), .A2(new_n475), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n616), .B1(new_n617), .B2(new_n604), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT90), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g419(.A(KEYINPUT90), .B(new_n616), .C1(new_n617), .C2(new_n604), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n614), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n612), .A2(new_n606), .A3(new_n613), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT89), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G113gat), .B(G141gat), .ZN(new_n628));
  INV_X1    g427(.A(G197gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT11), .B(G169gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT84), .Z(new_n634));
  NAND3_X1  g433(.A1(new_n614), .A2(new_n620), .A3(new_n621), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(new_n607), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n627), .A2(new_n634), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OAI22_X1  g437(.A1(new_n489), .A2(new_n494), .B1(new_n577), .B2(new_n582), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n480), .A2(new_n482), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT91), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n480), .A2(new_n482), .A3(KEYINPUT91), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n477), .B1(new_n645), .B2(new_n490), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT93), .B(G57gat), .Z(new_n647));
  OAI21_X1  g446(.A(new_n480), .B1(new_n647), .B2(new_n479), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n478), .A3(new_n488), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n568), .A2(new_n576), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n581), .A2(new_n575), .A3(new_n573), .A4(new_n564), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n646), .A2(new_n649), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n639), .A2(new_n640), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n495), .A2(KEYINPUT10), .A3(new_n583), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n639), .A2(KEYINPUT101), .A3(new_n652), .A4(new_n640), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G230gat), .A2(G233gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n639), .B2(new_n652), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n661), .B1(new_n658), .B2(new_n659), .ZN(new_n669));
  INV_X1    g468(.A(new_n666), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n663), .A2(new_n668), .A3(new_n666), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n638), .A2(new_n674), .ZN(new_n675));
  NOR4_X1   g474(.A1(new_n452), .A2(new_n514), .A3(new_n603), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n280), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT103), .B(G1gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1324gat));
  AND2_X1   g478(.A1(new_n676), .A2(new_n401), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT42), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n456), .B2(new_n680), .ZN(G1325gat));
  AOI21_X1  g483(.A(G15gat), .B1(new_n676), .B2(new_n443), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n676), .A2(G15gat), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n439), .B2(new_n686), .ZN(G1326gat));
  NAND2_X1  g486(.A1(new_n676), .A2(new_n394), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  AND2_X1   g489(.A1(new_n600), .A2(new_n592), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(KEYINPUT100), .A3(new_n597), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n593), .A2(new_n597), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(new_n691), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n452), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n514), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n675), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n520), .A3(new_n280), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n413), .A2(new_n442), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n445), .A2(new_n451), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n603), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT44), .B1(new_n452), .B2(new_n694), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n707), .A2(new_n697), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n708), .A2(new_n280), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n700), .B1(new_n520), .B2(new_n709), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n698), .A2(new_n521), .A3(new_n401), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT46), .Z(new_n712));
  AND2_X1   g511(.A1(new_n708), .A2(new_n401), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n521), .B2(new_n713), .ZN(G1329gat));
  AOI21_X1  g513(.A(G43gat), .B1(new_n698), .B2(new_n443), .ZN(new_n715));
  INV_X1    g514(.A(new_n439), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n517), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n715), .B1(new_n708), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1330gat));
  NAND3_X1  g519(.A1(new_n698), .A2(new_n515), .A3(new_n394), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n707), .A2(new_n394), .A3(new_n697), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G50gat), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n722), .A2(new_n723), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT48), .B(new_n721), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n722), .A2(G50gat), .ZN(new_n729));
  INV_X1    g528(.A(new_n721), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n731), .ZN(G1331gat));
  NOR2_X1   g531(.A1(new_n669), .A2(new_n670), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n671), .B(new_n733), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n694), .A2(new_n696), .A3(new_n637), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT105), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n452), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n280), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n647), .ZN(G1332gat));
  OR2_X1    g538(.A1(new_n737), .A2(KEYINPUT106), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(KEYINPUT106), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n400), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n737), .A2(new_n747), .A3(new_n443), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n716), .B1(new_n740), .B2(new_n741), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(new_n747), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1334gat));
  AOI21_X1  g551(.A(new_n395), .B1(new_n740), .B2(new_n741), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g553(.A1(new_n514), .A2(new_n637), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n695), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT51), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n695), .A2(new_n759), .A3(new_n756), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(new_n734), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n269), .A3(new_n280), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n755), .A2(new_n674), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n707), .A2(new_n280), .A3(new_n764), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(KEYINPUT108), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(G85gat), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n763), .A2(new_n768), .ZN(G1336gat));
  NAND3_X1  g568(.A1(new_n707), .A2(new_n401), .A3(new_n764), .ZN(new_n770));
  INV_X1    g569(.A(new_n580), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n400), .A2(G92gat), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n734), .A3(new_n760), .A4(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n759), .A2(KEYINPUT109), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n695), .B2(new_n756), .ZN(new_n778));
  AND4_X1   g577(.A1(new_n703), .A2(new_n603), .A3(new_n756), .A4(new_n777), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(new_n674), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n781), .A2(new_n773), .B1(new_n771), .B2(new_n770), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n776), .B1(new_n782), .B2(new_n775), .ZN(G1337gat));
  XOR2_X1   g582(.A(KEYINPUT111), .B(G99gat), .Z(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n762), .A2(new_n443), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n707), .A2(new_n439), .A3(new_n764), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n787), .A2(KEYINPUT110), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(KEYINPUT110), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(G1338gat));
  NOR3_X1   g590(.A1(new_n395), .A2(G106gat), .A3(new_n674), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT112), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n761), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n704), .B1(new_n703), .B2(new_n603), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n452), .A2(KEYINPUT44), .A3(new_n694), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n394), .B(new_n764), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G106gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n794), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n793), .B1(new_n778), .B2(new_n779), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT113), .B1(new_n802), .B2(KEYINPUT53), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n804), .B(new_n795), .C1(new_n799), .C2(new_n801), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n800), .B1(new_n803), .B2(new_n805), .ZN(G1339gat));
  NOR4_X1   g605(.A1(new_n603), .A2(new_n638), .A3(new_n514), .A4(new_n734), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n666), .B1(new_n660), .B2(KEYINPUT54), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n659), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n655), .A2(new_n810), .A3(new_n656), .A4(new_n657), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n660), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n660), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n808), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n669), .A2(new_n670), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n813), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n622), .A2(new_n633), .A3(new_n625), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n551), .A2(new_n474), .A3(new_n471), .A4(new_n529), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n613), .A2(new_n820), .A3(new_n615), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n613), .A2(new_n820), .A3(KEYINPUT114), .A4(new_n615), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n606), .B1(new_n612), .B2(new_n613), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT115), .B(new_n632), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n823), .B(new_n824), .C1(new_n605), .C2(new_n606), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT115), .B1(new_n829), .B2(new_n632), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n819), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n637), .A2(new_n818), .B1(new_n831), .B2(new_n674), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n694), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n632), .B1(new_n825), .B2(new_n826), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n836), .A2(new_n827), .B1(new_n636), .B2(new_n633), .ZN(new_n837));
  INV_X1    g636(.A(new_n818), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n603), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n807), .B1(new_n840), .B2(new_n514), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n444), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n440), .A2(new_n401), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n637), .ZN(new_n845));
  XOR2_X1   g644(.A(KEYINPUT116), .B(G113gat), .Z(new_n846));
  XNOR2_X1  g645(.A(new_n845), .B(new_n846), .ZN(G1340gat));
  NAND3_X1  g646(.A1(new_n842), .A2(new_n734), .A3(new_n843), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G120gat), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n204), .B2(new_n848), .ZN(G1341gat));
  NOR2_X1   g649(.A1(new_n844), .A2(new_n514), .ZN(new_n851));
  XOR2_X1   g650(.A(KEYINPUT117), .B(G127gat), .Z(new_n852));
  XNOR2_X1  g651(.A(new_n851), .B(new_n852), .ZN(G1342gat));
  NAND3_X1  g652(.A1(new_n842), .A2(new_n603), .A3(new_n843), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(G134gat), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(KEYINPUT56), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(KEYINPUT56), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(G134gat), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n856), .A2(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT119), .ZN(G1343gat));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n831), .B2(new_n674), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n734), .A2(new_n837), .A3(KEYINPUT120), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT121), .B(new_n814), .C1(new_n815), .C2(new_n808), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n809), .A2(new_n812), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n814), .A2(KEYINPUT121), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n868), .B(new_n817), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n637), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n694), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n696), .B1(new_n873), .B2(new_n839), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n394), .B1(new_n874), .B2(new_n807), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(KEYINPUT57), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n696), .B1(new_n833), .B2(new_n839), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n394), .B1(new_n877), .B2(new_n807), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n716), .A2(new_n843), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(G141gat), .A3(new_n638), .ZN(new_n882));
  INV_X1    g681(.A(G141gat), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n878), .A2(new_n880), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n885), .B2(new_n637), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n863), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n887), .B(new_n888), .ZN(G1344gat));
  INV_X1    g688(.A(G148gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n884), .A2(new_n890), .A3(new_n734), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n893), .B(new_n394), .C1(new_n874), .C2(new_n807), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n674), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n716), .A3(new_n843), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n892), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  AOI211_X1 g699(.A(KEYINPUT59), .B(new_n890), .C1(new_n881), .C2(new_n734), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n891), .B1(new_n900), .B2(new_n901), .ZN(G1345gat));
  AOI21_X1  g701(.A(G155gat), .B1(new_n884), .B2(new_n696), .ZN(new_n903));
  INV_X1    g702(.A(new_n881), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(new_n514), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n905), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g705(.A(G162gat), .B1(new_n884), .B2(new_n603), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n904), .A2(new_n228), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n603), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n280), .A2(new_n400), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n842), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n638), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(G169gat), .ZN(G1348gat));
  AOI22_X1  g713(.A1(new_n912), .A2(new_n734), .B1(KEYINPUT123), .B2(G176gat), .ZN(new_n915));
  NOR2_X1   g714(.A1(KEYINPUT123), .A2(G176gat), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n915), .B(new_n916), .Z(G1349gat));
  NAND2_X1  g716(.A1(new_n912), .A2(new_n696), .ZN(new_n918));
  MUX2_X1   g717(.A(new_n311), .B(G183gat), .S(new_n918), .Z(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g719(.A1(new_n912), .A2(new_n603), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G190gat), .ZN(new_n922));
  XOR2_X1   g721(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(G190gat), .B2(new_n921), .ZN(G1351gat));
  NAND2_X1  g724(.A1(new_n716), .A2(new_n910), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n897), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G197gat), .B1(new_n928), .B2(new_n637), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n878), .A2(new_n926), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n629), .A3(new_n638), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1352gat));
  INV_X1    g731(.A(new_n926), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n898), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G204gat), .ZN(new_n935));
  INV_X1    g734(.A(new_n930), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n936), .A2(G204gat), .A3(new_n674), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT62), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n938), .ZN(G1353gat));
  NAND4_X1  g738(.A1(new_n896), .A2(KEYINPUT126), .A3(new_n696), .A4(new_n933), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n894), .A2(new_n895), .A3(new_n696), .A4(new_n933), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n940), .A2(G211gat), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT63), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT63), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n940), .A2(new_n946), .A3(G211gat), .A4(new_n943), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n454), .A3(new_n696), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT125), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT127), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n945), .A2(new_n952), .A3(new_n947), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1354gat));
  OAI21_X1  g753(.A(G218gat), .B1(new_n928), .B2(new_n694), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n694), .A2(G218gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n936), .B2(new_n956), .ZN(G1355gat));
endmodule


