//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G128), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n191), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n199), .A3(KEYINPUT64), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n190), .A2(new_n192), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT88), .ZN(new_n203));
  INV_X1    g017(.A(G224), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G953), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n205), .B(KEYINPUT87), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n202), .A2(new_n203), .B1(KEYINPUT7), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT1), .B1(new_n195), .B2(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n197), .A2(G128), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n194), .B(new_n196), .C1(KEYINPUT1), .C2(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n202), .B1(G125), .B2(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n207), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G110), .B(G122), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT80), .A3(G104), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n220), .A2(new_n216), .A3(KEYINPUT80), .A4(G104), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G107), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n218), .A2(new_n219), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n223), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n222), .A2(G107), .ZN(new_n226));
  OAI21_X1  g040(.A(G101), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT5), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G116), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(G113), .B(new_n231), .C1(new_n233), .C2(new_n229), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n232), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n218), .A2(new_n221), .A3(new_n223), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G101), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT4), .A3(new_n224), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n242), .A3(G101), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n233), .A2(new_n235), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n237), .A3(KEYINPUT68), .ZN(new_n246));
  OR3_X1    g060(.A1(new_n236), .A2(KEYINPUT68), .A3(new_n232), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI221_X1 g062(.A(new_n215), .B1(new_n228), .B2(new_n238), .C1(new_n244), .C2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n215), .B(KEYINPUT8), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n238), .A2(new_n228), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n238), .A2(new_n228), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n207), .A2(new_n213), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n214), .A2(new_n249), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G902), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n215), .ZN(new_n258));
  AND4_X1   g072(.A1(new_n247), .A2(new_n241), .A3(new_n246), .A4(new_n243), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n252), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n260), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n249), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT86), .A2(KEYINPUT6), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n258), .B(new_n262), .C1(new_n259), .C2(new_n252), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n213), .B(new_n206), .Z(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(G210), .B1(G237), .B2(G902), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n257), .A2(new_n267), .A3(new_n265), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(KEYINPUT89), .A3(new_n270), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n270), .A2(KEYINPUT89), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G214), .B1(G237), .B2(G902), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n274), .B(KEYINPUT85), .Z(new_n275));
  OAI21_X1  g089(.A(KEYINPUT90), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT90), .ZN(new_n277));
  INV_X1    g091(.A(new_n275), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n271), .A2(new_n272), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(KEYINPUT74), .A2(G125), .ZN(new_n281));
  INV_X1    g095(.A(G140), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(KEYINPUT74), .A2(G125), .A3(G140), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(KEYINPUT16), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT16), .ZN(new_n286));
  INV_X1    g100(.A(G125), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(G140), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n193), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n283), .A2(new_n284), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n292));
  XNOR2_X1  g106(.A(G125), .B(G140), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n291), .A2(KEYINPUT19), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n289), .B1(new_n294), .B2(new_n193), .ZN(new_n295));
  INV_X1    g109(.A(G237), .ZN(new_n296));
  INV_X1    g110(.A(G953), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(G214), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(new_n195), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G131), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n300), .B(KEYINPUT91), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n299), .A2(G131), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(G113), .B(G122), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n304), .B(new_n222), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n299), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT18), .ZN(new_n308));
  INV_X1    g122(.A(G131), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n299), .A2(KEYINPUT18), .A3(G131), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n293), .A2(new_n193), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(new_n290), .B2(new_n193), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n303), .A2(new_n306), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(G475), .A2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n314), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT91), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n300), .B(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT17), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n319), .B(new_n320), .C1(G131), .C2(new_n299), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n285), .A2(new_n288), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G146), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n285), .A2(new_n193), .A3(new_n288), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n301), .B2(KEYINPUT17), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n317), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n315), .B(new_n316), .C1(new_n327), .C2(new_n306), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT20), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n321), .A2(new_n326), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n305), .B1(new_n330), .B2(new_n317), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT20), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n315), .A4(new_n316), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n305), .A2(KEYINPUT93), .ZN(new_n334));
  AOI21_X1  g148(.A(G902), .B1(new_n327), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n327), .B2(new_n334), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n329), .A2(new_n333), .B1(new_n336), .B2(G475), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n210), .A2(G143), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT13), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n339), .B(KEYINPUT94), .C1(G128), .C2(new_n195), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n338), .A2(KEYINPUT13), .ZN(new_n341));
  OAI221_X1 g155(.A(G134), .B1(KEYINPUT94), .B2(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(G116), .B(G122), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(new_n216), .ZN(new_n344));
  XNOR2_X1  g158(.A(G128), .B(G143), .ZN(new_n345));
  INV_X1    g159(.A(G134), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n342), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n216), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT95), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n345), .B(new_n346), .ZN(new_n351));
  INV_X1    g165(.A(G116), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT14), .A3(G122), .ZN(new_n353));
  INV_X1    g167(.A(new_n343), .ZN(new_n354));
  OAI211_X1 g168(.A(G107), .B(new_n353), .C1(new_n354), .C2(KEYINPUT14), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n348), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT9), .B(G234), .ZN(new_n358));
  INV_X1    g172(.A(G217), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n358), .A2(new_n359), .A3(G953), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n357), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  XOR2_X1   g176(.A(KEYINPUT72), .B(G902), .Z(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G478), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT96), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(KEYINPUT15), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(KEYINPUT15), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n363), .ZN(new_n372));
  OR3_X1    g186(.A1(new_n361), .A2(new_n372), .A3(new_n370), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n337), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n297), .A2(G952), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(G234), .B2(G237), .ZN(new_n378));
  AOI211_X1 g192(.A(new_n297), .B(new_n363), .C1(G234), .C2(G237), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT21), .B(G898), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G221), .B1(new_n358), .B2(G902), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G469), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT11), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n346), .B2(G137), .ZN(new_n387));
  INV_X1    g201(.A(G137), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT11), .A3(G134), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n346), .A2(G137), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT65), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n387), .A2(new_n389), .A3(KEYINPUT65), .A4(new_n390), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(G131), .A3(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n387), .A2(new_n389), .A3(new_n309), .A4(new_n390), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n396), .A2(KEYINPUT66), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT66), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n393), .A2(new_n399), .A3(G131), .A4(new_n394), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT81), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n212), .A2(new_n403), .A3(new_n224), .A4(new_n227), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n209), .A2(new_n211), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT81), .B1(new_n228), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n228), .A2(new_n405), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT10), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n404), .A2(new_n406), .A3(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n212), .A2(KEYINPUT10), .A3(new_n224), .A4(new_n227), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n190), .A2(new_n192), .A3(new_n200), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n241), .A2(new_n415), .A3(new_n243), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n413), .A2(new_n401), .A3(new_n414), .A4(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n416), .A2(new_n414), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n420), .A2(KEYINPUT82), .A3(new_n401), .A4(new_n413), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n411), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n297), .A2(G227), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n428));
  INV_X1    g242(.A(new_n426), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n422), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n420), .A2(new_n413), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n402), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n426), .B1(new_n419), .B2(new_n421), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(new_n428), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n427), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n385), .B1(new_n436), .B2(new_n256), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n411), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n434), .A2(KEYINPUT84), .A3(new_n411), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n422), .A2(new_n432), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n426), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n385), .A3(new_n363), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n384), .B1(new_n438), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n280), .A2(new_n382), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(G472), .A2(G902), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n246), .A2(new_n247), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n398), .A2(new_n415), .A3(new_n400), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT30), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n388), .A2(G134), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n309), .B1(new_n453), .B2(new_n390), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n396), .A3(new_n212), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n451), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n452), .B1(new_n451), .B2(new_n456), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n450), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n451), .A2(new_n456), .A3(new_n248), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n296), .A2(new_n297), .A3(G210), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n461), .B(KEYINPUT27), .Z(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT26), .B(G101), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n462), .B(new_n463), .Z(new_n464));
  NAND3_X1  g278(.A1(new_n459), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT31), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT31), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n459), .A2(new_n467), .A3(new_n460), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT28), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n248), .B1(new_n451), .B2(new_n456), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT69), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n451), .A2(new_n456), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n450), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n460), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n473), .B1(new_n476), .B2(new_n472), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n460), .A2(new_n470), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n464), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT32), .B(new_n449), .C1(new_n469), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT73), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n459), .A2(new_n460), .ZN(new_n483));
  INV_X1    g297(.A(new_n464), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n477), .A2(new_n478), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n486), .B2(new_n484), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n478), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n476), .B2(KEYINPUT28), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT29), .A3(new_n464), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT71), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n491), .A2(new_n494), .A3(KEYINPUT29), .A4(new_n464), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n372), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G472), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n449), .B1(new_n469), .B2(new_n479), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT70), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT32), .ZN(new_n502));
  OAI211_X1 g316(.A(KEYINPUT70), .B(new_n449), .C1(new_n469), .C2(new_n479), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n482), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n359), .B1(new_n363), .B2(G234), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n297), .A2(G221), .A3(G234), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT78), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT22), .B(G137), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT79), .ZN(new_n512));
  INV_X1    g326(.A(G110), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT24), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT24), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G110), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(G119), .B(G128), .ZN(new_n518));
  OR3_X1    g332(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT77), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT77), .B1(new_n517), .B2(new_n518), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n230), .A2(G128), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n230), .A2(G128), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(KEYINPUT23), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT76), .B(G110), .Z(new_n525));
  OAI211_X1 g339(.A(new_n519), .B(new_n520), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n289), .B1(new_n193), .B2(new_n293), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n524), .A2(G110), .B1(new_n518), .B2(new_n517), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n285), .A2(new_n193), .A3(new_n288), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n528), .B1(new_n529), .B2(new_n289), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n528), .B(KEYINPUT75), .C1(new_n529), .C2(new_n289), .ZN(new_n533));
  AOI221_X4 g347(.A(new_n512), .B1(new_n526), .B2(new_n527), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n526), .A2(new_n527), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT79), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n511), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n532), .A2(new_n533), .B1(new_n526), .B2(new_n527), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n511), .B1(new_n539), .B2(KEYINPUT79), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n363), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n538), .A2(KEYINPUT25), .A3(new_n541), .A4(new_n363), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n507), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n506), .A2(G902), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT75), .B1(new_n325), .B2(new_n528), .ZN(new_n548));
  INV_X1    g362(.A(new_n533), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n536), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n512), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n539), .A2(KEYINPUT79), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n540), .B1(new_n553), .B2(new_n511), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n546), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n505), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n448), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(G101), .ZN(G3));
  OAI21_X1  g372(.A(new_n363), .B1(new_n469), .B2(new_n479), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G472), .ZN(new_n560));
  AND4_X1   g374(.A1(new_n555), .A2(new_n501), .A3(new_n503), .A4(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n275), .B1(new_n269), .B2(new_n270), .ZN(new_n562));
  INV_X1    g376(.A(new_n381), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n333), .A2(new_n329), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n336), .A2(G475), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n361), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n361), .B1(new_n570), .B2(new_n568), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n569), .A2(G478), .A3(new_n363), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n364), .A2(new_n365), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n564), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n561), .A2(new_n447), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT34), .B(G104), .Z(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G6));
  OR2_X1    g393(.A1(new_n329), .A2(KEYINPUT98), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n333), .A2(KEYINPUT98), .A3(new_n329), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n374), .A2(new_n566), .ZN(new_n583));
  AND4_X1   g397(.A1(new_n563), .A2(new_n582), .A3(new_n562), .A4(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n447), .A3(new_n561), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G107), .Z(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(G9));
  AOI21_X1  g401(.A(KEYINPUT25), .B1(new_n554), .B2(new_n363), .ZN(new_n588));
  INV_X1    g402(.A(new_n545), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n506), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT36), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n511), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n550), .B(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n547), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n590), .A2(KEYINPUT99), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n546), .B2(new_n595), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n382), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n501), .A2(new_n560), .A3(new_n503), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n601), .A2(new_n280), .A3(new_n447), .A4(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT37), .B(G110), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G12));
  AND2_X1   g420(.A1(new_n505), .A2(new_n447), .ZN(new_n607));
  INV_X1    g421(.A(new_n600), .ZN(new_n608));
  INV_X1    g422(.A(new_n562), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(G900), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n379), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT100), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n378), .B(KEYINPUT101), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT102), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n582), .A2(new_n583), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n607), .A2(new_n610), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G128), .ZN(G30));
  NAND2_X1  g434(.A1(new_n567), .A2(new_n374), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n275), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n608), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n273), .B(KEYINPUT38), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n446), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n383), .B1(new_n626), .B2(new_n437), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n616), .B(KEYINPUT39), .Z(new_n628));
  OR3_X1    g442(.A1(new_n627), .A2(KEYINPUT40), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT40), .B1(new_n627), .B2(new_n628), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n483), .A2(new_n484), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n256), .B1(new_n476), .B2(new_n464), .ZN(new_n632));
  OAI21_X1  g446(.A(G472), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n633), .B(KEYINPUT103), .Z(new_n634));
  NAND3_X1  g448(.A1(new_n482), .A2(new_n634), .A3(new_n504), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n625), .A2(new_n629), .A3(new_n630), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G143), .ZN(G45));
  NAND3_X1  g451(.A1(new_n567), .A2(new_n574), .A3(new_n616), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n607), .A2(new_n610), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G146), .ZN(G48));
  NAND2_X1  g455(.A1(new_n445), .A2(new_n363), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(G469), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n446), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n384), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n645), .A2(new_n576), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n556), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT41), .B(G113), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT104), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(G15));
  NAND4_X1  g464(.A1(new_n505), .A2(new_n645), .A3(new_n555), .A4(new_n584), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G116), .ZN(G18));
  NAND4_X1  g466(.A1(new_n643), .A2(new_n383), .A3(new_n446), .A4(new_n562), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n601), .A2(new_n505), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G119), .ZN(G21));
  OAI211_X1 g470(.A(new_n466), .B(new_n468), .C1(new_n464), .C2(new_n491), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n449), .B(KEYINPUT105), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n559), .A2(G472), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n659), .A2(new_n555), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n621), .A2(new_n609), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n645), .A2(new_n660), .A3(new_n563), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G122), .ZN(G24));
  AND2_X1   g477(.A1(new_n600), .A2(new_n659), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n654), .A2(new_n664), .A3(KEYINPUT106), .A4(new_n639), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n639), .A2(new_n600), .A3(new_n659), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n666), .B1(new_n667), .B2(new_n653), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G125), .ZN(G27));
  NAND2_X1  g484(.A1(new_n499), .A2(new_n502), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n498), .A2(new_n480), .A3(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n672), .A2(new_n555), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n275), .B1(new_n271), .B2(new_n272), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n674), .B(new_n383), .C1(new_n626), .C2(new_n437), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n673), .A2(KEYINPUT42), .A3(new_n639), .A4(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n676), .A2(new_n505), .A3(new_n555), .A4(new_n639), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n678), .A2(KEYINPUT107), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT107), .B1(new_n678), .B2(new_n679), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G131), .ZN(G33));
  NAND3_X1  g497(.A1(new_n556), .A2(new_n618), .A3(new_n676), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT108), .B(G134), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G36));
  INV_X1    g500(.A(new_n628), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n385), .A2(new_n256), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n385), .B1(new_n436), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n434), .A2(new_n428), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n434), .A2(new_n428), .B1(new_n402), .B2(new_n431), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n691), .A2(new_n692), .B1(new_n426), .B2(new_n423), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT45), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n688), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n446), .B1(new_n695), .B2(KEYINPUT46), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n697), .B(new_n688), .C1(new_n690), .C2(new_n694), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n383), .B(new_n687), .C1(new_n696), .C2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n693), .B2(KEYINPUT45), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n436), .A2(new_n689), .ZN(new_n703));
  OAI22_X1  g517(.A1(new_n702), .A2(new_n703), .B1(new_n385), .B2(new_n256), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n697), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n695), .A2(KEYINPUT46), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n446), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(KEYINPUT109), .A3(new_n383), .A4(new_n687), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n337), .A2(new_n574), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n602), .A2(new_n713), .A3(new_n600), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n713), .B1(new_n602), .B2(new_n600), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g532(.A(KEYINPUT44), .B(new_n712), .C1(new_n714), .C2(new_n715), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n719), .A2(KEYINPUT111), .A3(new_n674), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT111), .B1(new_n719), .B2(new_n674), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n709), .B(new_n718), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G137), .ZN(G39));
  NAND2_X1  g537(.A1(new_n707), .A2(new_n383), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT47), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n707), .A2(new_n726), .A3(new_n383), .ZN(new_n727));
  INV_X1    g541(.A(new_n674), .ZN(new_n728));
  NOR4_X1   g542(.A1(new_n505), .A2(new_n555), .A3(new_n638), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n725), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G140), .ZN(G42));
  NOR3_X1   g545(.A1(new_n710), .A2(new_n384), .A3(new_n275), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n624), .A2(new_n555), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(KEYINPUT49), .B2(new_n644), .ZN(new_n734));
  INV_X1    g548(.A(new_n635), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n734), .B(new_n735), .C1(KEYINPUT49), .C2(new_n644), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT53), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n619), .A2(new_n640), .A3(new_n669), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n546), .A2(new_n595), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n447), .A2(new_n661), .A3(new_n740), .A4(new_n616), .ZN(new_n741));
  OR3_X1    g555(.A1(new_n735), .A2(new_n741), .A3(KEYINPUT112), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT112), .B1(new_n735), .B2(new_n741), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n738), .A2(new_n739), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n619), .A2(new_n640), .A3(new_n669), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT52), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n375), .A2(new_n566), .A3(new_n616), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n505), .A2(new_n582), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n639), .A2(new_n659), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n600), .A3(new_n676), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n567), .A2(new_n573), .A3(new_n572), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n563), .A3(new_n376), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n280), .A2(new_n755), .A3(new_n447), .A4(new_n561), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n604), .A2(new_n756), .A3(new_n662), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n651), .A2(new_n655), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n556), .B1(new_n448), .B2(new_n646), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n752), .A2(new_n757), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n744), .A2(new_n747), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n682), .A2(new_n684), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n737), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n745), .A2(new_n746), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n760), .B1(new_n766), .B2(new_n739), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n739), .B1(new_n619), .B2(new_n669), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n737), .ZN(new_n769));
  INV_X1    g583(.A(new_n763), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n767), .A2(new_n769), .A3(new_n770), .A4(new_n747), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n764), .A2(new_n765), .A3(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n744), .A2(new_n747), .A3(new_n761), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT53), .B1(new_n773), .B2(new_n770), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n768), .A2(KEYINPUT53), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n762), .A2(new_n763), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n772), .B1(new_n777), .B2(new_n765), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n779));
  INV_X1    g593(.A(new_n614), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n712), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(new_n660), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n377), .B1(new_n782), .B2(new_n654), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n644), .A2(new_n728), .A3(new_n384), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n673), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n735), .A2(new_n784), .A3(new_n555), .A4(new_n378), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(new_n575), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n785), .A2(new_n786), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n788), .A2(new_n789), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n783), .A3(new_n787), .A4(new_n791), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT115), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n782), .A2(new_n674), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n725), .A2(new_n727), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n644), .A2(new_n383), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n797), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n624), .A2(new_n275), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n782), .A2(new_n645), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n782), .A2(KEYINPUT50), .A3(new_n645), .A4(new_n802), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n337), .A2(new_n573), .A3(new_n572), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n790), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n781), .A2(new_n784), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n809), .B1(new_n664), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n807), .A2(KEYINPUT51), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n796), .B1(new_n801), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n807), .A2(new_n811), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n799), .B(KEYINPUT113), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n797), .B1(new_n798), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n779), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n812), .A2(new_n801), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(KEYINPUT116), .A3(new_n818), .A4(new_n796), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n778), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(G952), .A2(G953), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n736), .B1(new_n824), .B2(new_n825), .ZN(G75));
  NOR2_X1   g640(.A1(new_n297), .A2(G952), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n363), .B1(new_n764), .B2(new_n771), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT56), .B1(new_n829), .B2(new_n268), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n261), .A2(new_n263), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(new_n264), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT55), .Z(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n828), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n830), .B2(new_n834), .ZN(G51));
  XNOR2_X1  g650(.A(new_n688), .B(KEYINPUT57), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n764), .A2(new_n771), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(KEYINPUT54), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n765), .B1(new_n764), .B2(new_n771), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n445), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n829), .A2(new_n694), .A3(new_n690), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n827), .B1(new_n842), .B2(new_n843), .ZN(G54));
  NAND2_X1  g658(.A1(new_n331), .A2(new_n315), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(KEYINPUT58), .A2(G475), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n829), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n846), .B1(new_n829), .B2(new_n847), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n848), .A2(new_n849), .A3(new_n827), .ZN(G60));
  AND2_X1   g664(.A1(new_n569), .A2(new_n571), .ZN(new_n851));
  NAND2_X1  g665(.A1(G478), .A2(G902), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT59), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n851), .B1(new_n778), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n851), .A2(new_n853), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n839), .B2(new_n840), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n828), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n854), .A2(new_n857), .ZN(G63));
  NAND2_X1  g672(.A1(G217), .A2(G902), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT60), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n764), .B2(new_n771), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(new_n554), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n593), .B(KEYINPUT117), .Z(new_n863));
  AOI21_X1  g677(.A(new_n827), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n861), .A2(new_n863), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT61), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT118), .B1(new_n861), .B2(new_n863), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n862), .B(new_n864), .C1(new_n870), .C2(KEYINPUT61), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(G66));
  OAI21_X1  g686(.A(G953), .B1(new_n380), .B2(new_n204), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n874), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n873), .B1(new_n876), .B2(G953), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n831), .B1(G898), .B2(new_n297), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n877), .B(new_n878), .ZN(G69));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n722), .A2(new_n880), .A3(new_n738), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n722), .B2(new_n738), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n709), .A2(new_n661), .A3(new_n673), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n682), .A2(new_n884), .A3(new_n684), .A4(new_n730), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n297), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n457), .A2(new_n458), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(new_n294), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n611), .B2(new_n297), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n889), .A2(KEYINPUT122), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n297), .B1(G227), .B2(G900), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n753), .A2(new_n376), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n556), .A2(new_n687), .A3(new_n676), .A4(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n730), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n636), .A2(new_n619), .A3(new_n640), .A4(new_n669), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT62), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n899), .A2(KEYINPUT62), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n901), .A2(new_n902), .A3(new_n722), .A4(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n722), .A3(new_n900), .A4(new_n898), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT120), .ZN(new_n906));
  AOI21_X1  g720(.A(G953), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n892), .B(new_n895), .C1(new_n907), .C2(new_n889), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n890), .B1(new_n886), .B2(new_n297), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n889), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n893), .B(new_n894), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n908), .A2(new_n911), .ZN(G72));
  NAND3_X1  g726(.A1(new_n904), .A2(new_n906), .A3(new_n876), .ZN(new_n913));
  NAND2_X1  g727(.A1(G472), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT124), .ZN(new_n915));
  XOR2_X1   g729(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n631), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n485), .A3(new_n917), .ZN(new_n920));
  OAI22_X1  g734(.A1(new_n918), .A2(new_n919), .B1(new_n777), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n876), .B(new_n885), .C1(new_n881), .C2(new_n882), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n923), .A3(new_n917), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n485), .B(KEYINPUT126), .Z(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n923), .B1(new_n922), .B2(new_n917), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n828), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(KEYINPUT127), .B(new_n828), .C1(new_n926), .C2(new_n927), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n921), .B1(new_n930), .B2(new_n931), .ZN(G57));
endmodule


