//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971;
  XOR2_X1   g000(.A(G183gat), .B(G211gat), .Z(new_n202));
  OR2_X1    g001(.A1(G57gat), .A2(G64gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G57gat), .A2(G64gat), .ZN(new_n204));
  AND2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206));
  INV_X1    g005(.A(G71gat), .ZN(new_n207));
  INV_X1    g006(.A(G78gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G71gat), .B(G78gat), .Z(new_n210));
  OAI211_X1 g009(.A(new_n205), .B(new_n209), .C1(new_n210), .C2(KEYINPUT96), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n203), .A3(new_n204), .ZN(new_n212));
  XNOR2_X1  g011(.A(G71gat), .B(G78gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n203), .A2(KEYINPUT96), .A3(new_n204), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n216), .A2(KEYINPUT21), .ZN(new_n217));
  NAND2_X1  g016(.A1(G231gat), .A2(G233gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G127gat), .B(G155gat), .ZN(new_n220));
  XOR2_X1   g019(.A(new_n220), .B(KEYINPUT97), .Z(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n219), .A2(new_n222), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n202), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n225), .ZN(new_n227));
  INV_X1    g026(.A(new_n202), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT16), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n230), .B1(new_n234), .B2(KEYINPUT93), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(G1gat), .B2(new_n231), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI221_X1 g036(.A(new_n234), .B1(KEYINPUT93), .B2(new_n230), .C1(G1gat), .C2(new_n231), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(KEYINPUT21), .B2(new_n216), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n226), .A2(new_n229), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(new_n226), .B2(new_n229), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(G43gat), .A2(G50gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(G43gat), .A2(G50gat), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT15), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G43gat), .ZN(new_n250));
  INV_X1    g049(.A(G50gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT15), .ZN(new_n253));
  NAND2_X1  g052(.A1(G43gat), .A2(G50gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G29gat), .ZN(new_n257));
  INV_X1    g056(.A(G36gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT14), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT14), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(G29gat), .B2(G36gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(G29gat), .A2(G36gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT91), .B1(new_n256), .B2(new_n263), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT91), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n249), .A4(new_n255), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT90), .B1(new_n265), .B2(new_n249), .ZN(new_n269));
  INV_X1    g068(.A(new_n249), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT90), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(new_n263), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(KEYINPUT17), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G85gat), .A2(G92gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT7), .ZN(new_n276));
  NAND2_X1  g075(.A1(G99gat), .A2(G106gat), .ZN(new_n277));
  INV_X1    g076(.A(G85gat), .ZN(new_n278));
  INV_X1    g077(.A(G92gat), .ZN(new_n279));
  AOI22_X1  g078(.A1(KEYINPUT8), .A2(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(G99gat), .A2(G106gat), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT98), .B1(new_n282), .B2(new_n277), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(KEYINPUT98), .A3(new_n277), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n285), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n276), .B(new_n280), .C1(new_n287), .C2(new_n283), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT92), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n264), .A2(new_n267), .B1(new_n269), .B2(new_n272), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(KEYINPUT17), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n268), .A2(new_n273), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT17), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT92), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n290), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G190gat), .B(G218gat), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n289), .ZN(new_n301));
  NAND2_X1  g100(.A1(G232gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n294), .A2(new_n301), .B1(KEYINPUT41), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n298), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n304), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n299), .B1(new_n297), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n303), .A2(KEYINPUT41), .ZN(new_n308));
  XNOR2_X1  g107(.A(G134gat), .B(G162gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n305), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n310), .B1(new_n305), .B2(new_n307), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n246), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G120gat), .B(G148gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(G176gat), .B(G204gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(KEYINPUT99), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n284), .A2(new_n318), .A3(new_n285), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n216), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n289), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n216), .A2(new_n286), .A3(new_n288), .A4(new_n319), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G230gat), .A2(G233gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n317), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n324), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT10), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(new_n327), .A3(new_n322), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n301), .A2(KEYINPUT10), .A3(new_n216), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n323), .A2(new_n324), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n324), .B(KEYINPUT100), .Z(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n328), .B2(new_n329), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n332), .B1(new_n336), .B2(new_n317), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n314), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT95), .ZN(new_n340));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT0), .ZN(new_n342));
  XNOR2_X1  g141(.A(G57gat), .B(G85gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  INV_X1    g143(.A(KEYINPUT2), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n345), .B1(G155gat), .B2(G162gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT81), .ZN(new_n347));
  INV_X1    g146(.A(G148gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G141gat), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT79), .B(G141gat), .Z(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n348), .ZN(new_n351));
  XNOR2_X1  g150(.A(G155gat), .B(G162gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n352), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT80), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n347), .A2(new_n351), .A3(new_n354), .A4(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G141gat), .B(G148gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n355), .B1(new_n358), .B2(new_n346), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT3), .ZN(new_n361));
  INV_X1    g160(.A(G113gat), .ZN(new_n362));
  INV_X1    g161(.A(G120gat), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT1), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(new_n362), .B2(new_n363), .ZN(new_n365));
  XNOR2_X1  g164(.A(G127gat), .B(G134gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT69), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n365), .A2(KEYINPUT69), .A3(new_n367), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT70), .B(G120gat), .ZN(new_n372));
  OR2_X1    g171(.A1(new_n372), .A2(new_n362), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n366), .A2(new_n364), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n370), .A2(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n357), .A2(new_n377), .A3(new_n359), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n376), .B2(new_n360), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n357), .A2(new_n359), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n375), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n379), .B(new_n381), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT5), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n384), .B1(new_n376), .B2(new_n360), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n382), .A2(new_n375), .A3(KEYINPUT4), .ZN(new_n389));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(new_n386), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n388), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n379), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n360), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT83), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n383), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n376), .A2(KEYINPUT83), .A3(new_n360), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n390), .B1(new_n400), .B2(KEYINPUT5), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n344), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(KEYINPUT5), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n391), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n386), .A2(new_n385), .B1(new_n393), .B2(new_n379), .ZN(new_n405));
  INV_X1    g204(.A(new_n344), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT6), .A4(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT27), .B(G183gat), .ZN(new_n412));
  INV_X1    g211(.A(G190gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT28), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(G169gat), .A2(G176gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(KEYINPUT67), .A3(KEYINPUT26), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n418), .A2(KEYINPUT67), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT26), .ZN(new_n421));
  INV_X1    g220(.A(G169gat), .ZN(new_n422));
  INV_X1    g221(.A(G176gat), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n417), .B(new_n419), .C1(new_n420), .C2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n416), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT66), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n417), .B1(new_n431), .B2(KEYINPUT24), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT24), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(KEYINPUT66), .ZN(new_n434));
  OAI221_X1 g233(.A(new_n430), .B1(G183gat), .B2(G190gat), .C1(new_n432), .C2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT23), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(G169gat), .B2(G176gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT65), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n422), .A2(new_n423), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(KEYINPUT23), .B2(new_n418), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n435), .A2(new_n439), .A3(KEYINPUT25), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n417), .A2(new_n433), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n443), .B(new_n430), .C1(G183gat), .C2(G190gat), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n439), .A2(new_n444), .A3(new_n441), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n445), .B2(KEYINPUT25), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n416), .A2(KEYINPUT68), .A3(new_n426), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT74), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n429), .A2(new_n446), .A3(KEYINPUT74), .A4(new_n447), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT29), .B1(new_n446), .B2(new_n427), .ZN(new_n455));
  OR3_X1    g254(.A1(new_n455), .A2(KEYINPUT76), .A3(new_n452), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT73), .B(G197gat), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n457), .A2(G204gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(G204gat), .ZN(new_n459));
  INV_X1    g258(.A(G211gat), .ZN(new_n460));
  INV_X1    g259(.A(G218gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI22_X1  g261(.A1(new_n458), .A2(new_n459), .B1(KEYINPUT22), .B2(new_n462), .ZN(new_n463));
  XOR2_X1   g262(.A(G211gat), .B(G218gat), .Z(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT76), .B1(new_n455), .B2(new_n452), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n454), .A2(new_n456), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(G8gat), .B(G36gat), .Z(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT77), .ZN(new_n469));
  XNOR2_X1  g268(.A(G64gat), .B(G92gat), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n469), .B(new_n470), .Z(new_n471));
  XOR2_X1   g270(.A(KEYINPUT75), .B(KEYINPUT29), .Z(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(new_n452), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n450), .A2(new_n453), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n465), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n446), .A2(new_n452), .A3(new_n427), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n467), .A2(new_n471), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT78), .ZN(new_n480));
  INV_X1    g279(.A(new_n471), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n467), .A2(new_n478), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n480), .A2(KEYINPUT30), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT30), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(KEYINPUT78), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n411), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G78gat), .B(G106gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(new_n251), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G22gat), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n377), .B1(new_n476), .B2(new_n473), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n360), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n465), .B1(new_n378), .B2(new_n472), .ZN(new_n493));
  NAND2_X1  g292(.A1(G228gat), .A2(G233gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n465), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n382), .B1(new_n499), .B2(new_n377), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n495), .B1(new_n500), .B2(new_n493), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n497), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n503), .B1(new_n497), .B2(new_n501), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n490), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n506), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(new_n489), .A3(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n486), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n448), .A2(new_n375), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n429), .A2(new_n376), .A3(new_n446), .A4(new_n447), .ZN(new_n514));
  NAND2_X1  g313(.A1(G227gat), .A2(G233gat), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n515), .B(KEYINPUT64), .Z(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT32), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT33), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G15gat), .B(G43gat), .Z(new_n521));
  XNOR2_X1  g320(.A(G71gat), .B(G99gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n518), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n523), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n517), .B(KEYINPUT32), .C1(new_n519), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT71), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n516), .A2(KEYINPUT34), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n513), .B2(new_n514), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n514), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n515), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n532), .B2(KEYINPUT34), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n527), .A2(KEYINPUT71), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(KEYINPUT36), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n524), .A2(new_n533), .A3(new_n526), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n533), .B1(new_n524), .B2(new_n526), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n512), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n385), .A2(new_n391), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(KEYINPUT39), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(new_n406), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT85), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n400), .B2(new_n390), .ZN(new_n549));
  AOI211_X1 g348(.A(KEYINPUT85), .B(new_n391), .C1(new_n398), .C2(new_n399), .ZN(new_n550));
  OAI211_X1 g349(.A(KEYINPUT39), .B(new_n545), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT40), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n407), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n547), .A2(new_n551), .A3(KEYINPUT40), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n483), .A2(new_n485), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n511), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n454), .A2(new_n456), .A3(new_n466), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n476), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT86), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n476), .B1(new_n475), .B2(new_n477), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n561), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT37), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT38), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n482), .A2(new_n481), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT37), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(new_n471), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n409), .A2(new_n410), .A3(new_n479), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT87), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT87), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n567), .B(new_n481), .C1(new_n482), .C2(KEYINPUT37), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n562), .A2(new_n561), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(new_n564), .A3(new_n560), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n575), .B1(new_n577), .B2(KEYINPUT37), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n409), .A2(new_n410), .A3(new_n479), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n574), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n482), .A2(KEYINPUT37), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n567), .B1(new_n570), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n573), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n544), .B1(new_n558), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n536), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n535), .B1(new_n527), .B2(KEYINPUT71), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n480), .A2(KEYINPUT30), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n589), .A2(new_n568), .A3(new_n485), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n588), .A2(new_n590), .A3(new_n411), .A4(new_n510), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT35), .B1(new_n507), .B2(new_n509), .ZN(new_n592));
  INV_X1    g391(.A(new_n541), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(KEYINPUT88), .A3(new_n539), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT88), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(new_n540), .B2(new_n541), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n592), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n486), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n591), .A2(KEYINPUT35), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n585), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT94), .ZN(new_n601));
  INV_X1    g400(.A(new_n239), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n292), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n294), .A2(new_n239), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT13), .Z(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G197gat), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT11), .B(G169gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n602), .A2(new_n274), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n293), .B2(new_n296), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n604), .A2(KEYINPUT18), .A3(new_n606), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n608), .B(new_n613), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n239), .B1(new_n292), .B2(KEYINPUT17), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT92), .B1(new_n294), .B2(new_n295), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n292), .A2(new_n291), .A3(KEYINPUT17), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT18), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n601), .B1(new_n617), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT18), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n615), .B2(new_n622), .ZN(new_n627));
  INV_X1    g426(.A(new_n616), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n612), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n607), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n632), .B1(new_n603), .B2(new_n604), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n627), .A2(KEYINPUT94), .A3(new_n629), .A4(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n627), .A2(new_n629), .A3(new_n608), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n631), .B(KEYINPUT89), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n625), .A2(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n340), .B1(new_n600), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n625), .A2(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g441(.A(KEYINPUT95), .B(new_n642), .C1(new_n585), .C2(new_n599), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n339), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n411), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g446(.A(new_n230), .B1(new_n644), .B2(new_n557), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  NAND3_X1  g448(.A1(new_n644), .A2(new_n557), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n644), .A2(KEYINPUT42), .A3(new_n557), .A4(new_n649), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n653), .A2(KEYINPUT102), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(KEYINPUT102), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(G1325gat));
  INV_X1    g455(.A(new_n594), .ZN(new_n657));
  INV_X1    g456(.A(new_n596), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(G15gat), .B1(new_n644), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n543), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n537), .A2(KEYINPUT103), .A3(new_n542), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(G15gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT104), .Z(new_n666));
  AOI21_X1  g465(.A(new_n660), .B1(new_n644), .B2(new_n666), .ZN(G1326gat));
  NAND2_X1  g466(.A1(new_n644), .A2(new_n511), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT43), .B(G22gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  NAND2_X1  g469(.A1(new_n639), .A2(new_n643), .ZN(new_n671));
  INV_X1    g470(.A(new_n313), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n245), .A2(new_n672), .A3(new_n337), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n257), .A3(new_n645), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT45), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n674), .A2(KEYINPUT45), .A3(new_n257), .A4(new_n645), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n591), .A2(KEYINPUT35), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n597), .A2(new_n598), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n554), .A2(new_n555), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n510), .B1(new_n682), .B2(new_n590), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n571), .A2(new_n572), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n582), .B1(new_n684), .B2(new_n574), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n683), .B1(new_n685), .B2(new_n573), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n662), .A2(new_n512), .A3(new_n663), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n681), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n313), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n681), .B1(new_n686), .B2(new_n544), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n672), .A2(new_n690), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n689), .A2(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n246), .A2(new_n642), .A3(new_n338), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n645), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G29gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n677), .A2(new_n678), .A3(new_n697), .ZN(G1328gat));
  NOR2_X1   g497(.A1(new_n590), .A2(G36gat), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT95), .B1(new_n691), .B2(new_n642), .ZN(new_n700));
  INV_X1    g499(.A(new_n643), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n673), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT46), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n671), .A2(new_n704), .A3(new_n673), .A4(new_n699), .ZN(new_n705));
  INV_X1    g504(.A(new_n663), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT103), .B1(new_n537), .B2(new_n542), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n510), .B1(new_n590), .B2(new_n411), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n558), .A2(new_n584), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n599), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n690), .B1(new_n711), .B2(new_n672), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n691), .A2(new_n692), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n712), .A2(new_n713), .A3(new_n557), .A4(new_n695), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G36gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n703), .A2(new_n705), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT105), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n715), .A3(new_n705), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(G1329gat));
  NAND4_X1  g519(.A1(new_n712), .A2(new_n713), .A3(new_n664), .A4(new_n695), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(G43gat), .ZN(new_n722));
  INV_X1    g521(.A(new_n659), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(G43gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n671), .A2(new_n673), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT47), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  AOI211_X1 g528(.A(KEYINPUT106), .B(new_n729), .C1(new_n722), .C2(new_n725), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(new_n730), .ZN(G1330gat));
  XOR2_X1   g530(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n732));
  NOR2_X1   g531(.A1(new_n510), .A2(G50gat), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n673), .B(new_n733), .C1(new_n700), .C2(new_n701), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n712), .A2(new_n713), .A3(new_n511), .A4(new_n695), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G50gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n732), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(KEYINPUT48), .A3(new_n734), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(G1331gat));
  NAND4_X1  g541(.A1(new_n314), .A2(new_n640), .A3(new_n641), .A4(new_n337), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n711), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n645), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT109), .B(G57gat), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1332gat));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n557), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT49), .B(G64gat), .Z(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(G1333gat));
  NAND3_X1  g550(.A1(new_n744), .A2(new_n207), .A3(new_n659), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n744), .A2(new_n664), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n207), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n744), .A2(new_n511), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT112), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT111), .B(G78gat), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1335gat));
  NOR3_X1   g559(.A1(new_n245), .A2(new_n642), .A3(new_n338), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n693), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n645), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G85gat), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n245), .A2(new_n642), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n688), .A2(new_n313), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  OR3_X1    g568(.A1(new_n768), .A2(new_n769), .A3(KEYINPUT113), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT113), .B1(new_n768), .B2(new_n769), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n337), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n645), .A2(new_n278), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n764), .B1(new_n772), .B2(new_n773), .ZN(G1336gat));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n590), .A2(G92gat), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n337), .B(new_n776), .C1(new_n768), .C2(new_n769), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n712), .A2(new_n713), .A3(new_n557), .A4(new_n761), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n775), .B(new_n777), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(G92gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT52), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(G1337gat));
  NAND2_X1  g585(.A1(new_n762), .A2(new_n664), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G99gat), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n723), .A2(G99gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n772), .B2(new_n789), .ZN(G1338gat));
  NAND4_X1  g589(.A1(new_n712), .A2(new_n713), .A3(new_n511), .A4(new_n761), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n791), .A2(G106gat), .B1(KEYINPUT115), .B2(KEYINPUT53), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n510), .A2(G106gat), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n337), .B(new_n793), .C1(new_n768), .C2(new_n769), .ZN(new_n794));
  OR2_X1    g593(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n792), .B2(new_n794), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(G1339gat));
  NAND2_X1  g597(.A1(new_n640), .A2(new_n337), .ZN(new_n799));
  INV_X1    g598(.A(new_n612), .ZN(new_n800));
  INV_X1    g599(.A(new_n606), .ZN(new_n801));
  INV_X1    g600(.A(new_n604), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n615), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n603), .A2(new_n604), .A3(new_n632), .ZN(new_n804));
  AOI211_X1 g603(.A(KEYINPUT116), .B(new_n800), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n293), .A2(new_n296), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n802), .B1(new_n807), .B2(new_n618), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n804), .B1(new_n808), .B2(new_n606), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n806), .B1(new_n809), .B2(new_n612), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n328), .A2(new_n334), .A3(new_n329), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n813), .A2(new_n330), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n328), .A2(new_n329), .ZN(new_n816));
  INV_X1    g615(.A(new_n334), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n317), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n812), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n816), .A2(new_n324), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n328), .A2(new_n329), .A3(new_n334), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n317), .B1(new_n335), .B2(new_n814), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(new_n332), .A3(new_n826), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n799), .A2(new_n811), .B1(new_n638), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n672), .ZN(new_n829));
  INV_X1    g628(.A(new_n811), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n821), .A2(new_n332), .A3(new_n826), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n830), .A2(new_n640), .A3(new_n313), .A4(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n245), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NOR4_X1   g632(.A1(new_n246), .A2(new_n642), .A3(new_n313), .A4(new_n337), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT117), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n642), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n640), .B(new_n337), .C1(new_n810), .C2(new_n805), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n313), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n313), .A2(new_n640), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n839), .A2(new_n811), .A3(new_n827), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n246), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n314), .A2(new_n638), .A3(new_n338), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n835), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n511), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n846), .A2(new_n645), .A3(new_n590), .A4(new_n659), .ZN(new_n847));
  OAI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n638), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n835), .A2(new_n844), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n588), .A2(new_n510), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n557), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n645), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT118), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n642), .A2(new_n362), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n848), .B1(new_n853), .B2(new_n854), .ZN(G1340gat));
  OAI21_X1  g654(.A(G120gat), .B1(new_n847), .B2(new_n338), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n337), .A2(new_n372), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n853), .B2(new_n857), .ZN(G1341gat));
  OAI21_X1  g657(.A(G127gat), .B1(new_n847), .B2(new_n246), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n246), .A2(G127gat), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n852), .B2(new_n860), .ZN(G1342gat));
  OR2_X1    g660(.A1(new_n672), .A2(G134gat), .ZN(new_n862));
  OR3_X1    g661(.A1(new_n852), .A2(KEYINPUT119), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT119), .B1(new_n852), .B2(new_n862), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n863), .A2(new_n865), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT56), .ZN(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n847), .B2(new_n672), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n868), .A2(new_n869), .A3(new_n871), .A4(new_n872), .ZN(G1343gat));
  NOR2_X1   g672(.A1(new_n845), .A2(new_n411), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n662), .A2(new_n511), .A3(new_n663), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n557), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n877), .A2(G141gat), .A3(new_n638), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n664), .A2(new_n411), .A3(new_n557), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n511), .B1(new_n833), .B2(new_n834), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT57), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n849), .A2(new_n511), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n879), .B(new_n881), .C1(new_n882), .C2(KEYINPUT57), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n638), .ZN(new_n884));
  INV_X1    g683(.A(new_n350), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n878), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT58), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n878), .B(new_n888), .C1(new_n885), .C2(new_n884), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(G1344gat));
  INV_X1    g689(.A(new_n877), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n348), .A3(new_n337), .ZN(new_n892));
  XNOR2_X1  g691(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n849), .A2(KEYINPUT57), .A3(new_n511), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n337), .A3(new_n879), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n893), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  INV_X1    g699(.A(new_n883), .ZN(new_n901));
  AOI211_X1 g700(.A(KEYINPUT59), .B(new_n348), .C1(new_n901), .C2(new_n337), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n892), .B1(new_n900), .B2(new_n902), .ZN(G1345gat));
  OAI21_X1  g702(.A(G155gat), .B1(new_n883), .B2(new_n246), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n246), .A2(G155gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n877), .B2(new_n905), .ZN(G1346gat));
  AOI21_X1  g705(.A(G162gat), .B1(new_n891), .B2(new_n313), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n313), .A2(G162gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n901), .B2(new_n908), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n590), .A2(new_n645), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n723), .A2(new_n911), .ZN(new_n912));
  AND4_X1   g711(.A1(G169gat), .A2(new_n846), .A3(new_n642), .A4(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n849), .B2(new_n411), .ZN(new_n915));
  AOI211_X1 g714(.A(KEYINPUT122), .B(new_n645), .C1(new_n835), .C2(new_n844), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n850), .A2(new_n590), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n642), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n913), .B1(new_n919), .B2(new_n422), .ZN(G1348gat));
  NAND4_X1  g719(.A1(new_n846), .A2(G176gat), .A3(new_n337), .A4(new_n912), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n337), .B(new_n918), .C1(new_n915), .C2(new_n916), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n922), .A2(new_n923), .A3(new_n423), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n922), .B2(new_n423), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g727(.A(KEYINPUT124), .B(new_n921), .C1(new_n924), .C2(new_n925), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1349gat));
  NAND3_X1  g729(.A1(new_n846), .A2(new_n245), .A3(new_n912), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  AOI22_X1  g731(.A1(new_n931), .A2(G183gat), .B1(new_n932), .B2(KEYINPUT60), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n245), .A2(new_n412), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n846), .A2(new_n313), .A3(new_n912), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(G190gat), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n939), .B2(G190gat), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n313), .A2(new_n413), .ZN(new_n944));
  OAI22_X1  g743(.A1(new_n942), .A2(new_n943), .B1(new_n934), .B2(new_n944), .ZN(G1351gat));
  XNOR2_X1  g744(.A(new_n897), .B(KEYINPUT126), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n664), .A2(new_n911), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(G197gat), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n948), .A2(new_n949), .A3(new_n638), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n875), .A2(new_n590), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n917), .A2(new_n642), .A3(new_n951), .ZN(new_n952));
  AOI22_X1  g751(.A1(new_n946), .A2(new_n950), .B1(new_n949), .B2(new_n952), .ZN(G1352gat));
  AND2_X1   g752(.A1(new_n897), .A2(KEYINPUT126), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n897), .A2(KEYINPUT126), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n337), .B(new_n947), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G204gat), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n338), .A2(G204gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n917), .A2(new_n951), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n957), .A2(new_n960), .A3(new_n961), .ZN(G1353gat));
  NAND4_X1  g761(.A1(new_n917), .A2(new_n460), .A3(new_n245), .A4(new_n951), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n898), .A2(new_n245), .A3(new_n947), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  AND2_X1   g766(.A1(new_n946), .A2(new_n947), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n313), .A2(G218gat), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT127), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n917), .A2(new_n313), .A3(new_n951), .ZN(new_n971));
  AOI22_X1  g770(.A1(new_n968), .A2(new_n970), .B1(new_n461), .B2(new_n971), .ZN(G1355gat));
endmodule


