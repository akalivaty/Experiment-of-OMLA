//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n188));
  INV_X1    g002(.A(G113), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n187), .A2(new_n188), .A3(new_n189), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n191));
  AOI22_X1  g005(.A1(new_n190), .A2(new_n191), .B1(KEYINPUT2), .B2(G113), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT69), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G116), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n193), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n192), .B(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT30), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g020(.A1(KEYINPUT66), .A2(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT66), .A2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(G143), .B2(new_n202), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n206), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n203), .A3(new_n205), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G137), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G137), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G134), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(KEYINPUT65), .A3(G137), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n212), .A2(new_n215), .B1(new_n223), .B2(G131), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n220), .A2(G134), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT11), .B1(new_n216), .B2(G137), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT11), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n220), .A3(G134), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n225), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT64), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n228), .ZN(new_n232));
  AND4_X1   g046(.A1(KEYINPUT64), .A2(new_n232), .A3(new_n230), .A4(new_n217), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n224), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n235));
  OR2_X1    g049(.A1(new_n229), .A2(new_n230), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n233), .B2(new_n231), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n238));
  XNOR2_X1  g052(.A(G143), .B(G146), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT0), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(new_n213), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AND4_X1   g057(.A1(KEYINPUT0), .A2(new_n203), .A3(new_n205), .A4(G128), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n238), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n241), .ZN(new_n246));
  INV_X1    g060(.A(new_n242), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n206), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n239), .A2(KEYINPUT0), .A3(G128), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT70), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n234), .A2(new_n235), .B1(new_n237), .B2(new_n251), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n224), .B(KEYINPUT71), .C1(new_n231), .C2(new_n233), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n201), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n234), .A2(KEYINPUT67), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n224), .B(new_n256), .C1(new_n231), .C2(new_n233), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n243), .A2(new_n244), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n237), .A2(new_n258), .ZN(new_n259));
  AND4_X1   g073(.A1(new_n201), .A2(new_n255), .A3(new_n257), .A4(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n200), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n252), .A2(new_n199), .A3(new_n253), .ZN(new_n262));
  NOR2_X1   g076(.A1(G237), .A2(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n261), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT31), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n233), .A2(new_n231), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n212), .A2(new_n215), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n223), .A2(G131), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n235), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n237), .A2(new_n251), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(new_n253), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(new_n200), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n234), .A2(KEYINPUT67), .B1(new_n237), .B2(new_n258), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n199), .B1(new_n278), .B2(new_n257), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT28), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n234), .A2(new_n199), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT28), .B1(new_n281), .B2(new_n275), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n267), .B(KEYINPUT72), .Z(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n276), .A2(KEYINPUT30), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n278), .A2(new_n201), .A3(new_n257), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n277), .B1(new_n290), .B2(new_n200), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n267), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n269), .A2(new_n287), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(G472), .A2(G902), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n294), .A2(KEYINPUT32), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT32), .B1(new_n294), .B2(new_n295), .ZN(new_n297));
  INV_X1    g111(.A(G472), .ZN(new_n298));
  INV_X1    g112(.A(new_n267), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n199), .B1(new_n288), .B2(new_n289), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(new_n277), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n301), .B(new_n302), .C1(new_n284), .C2(new_n286), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT28), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n276), .A2(new_n200), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(new_n262), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(new_n282), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n299), .A2(new_n302), .ZN(new_n308));
  AOI21_X1  g122(.A(G902), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n298), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n296), .A2(new_n297), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G217), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(G234), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n194), .B1(new_n207), .B2(new_n208), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n213), .A2(G119), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT73), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT24), .B(G110), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g134(.A1(KEYINPUT24), .A2(G110), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT24), .A2(G110), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(KEYINPUT74), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n208), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT66), .A2(G128), .ZN(new_n326));
  OAI21_X1  g140(.A(G119), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n328));
  INV_X1    g142(.A(new_n316), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n317), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n327), .A2(KEYINPUT23), .A3(new_n329), .ZN(new_n332));
  OR3_X1    g146(.A1(new_n194), .A2(KEYINPUT23), .A3(G128), .ZN(new_n333));
  AOI21_X1  g147(.A(G110), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT76), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n317), .A2(new_n324), .A3(new_n330), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n332), .A2(new_n333), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(G110), .ZN(new_n339));
  INV_X1    g153(.A(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G125), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G140), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT16), .ZN(new_n344));
  OR3_X1    g158(.A1(new_n342), .A2(KEYINPUT16), .A3(G140), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G146), .ZN(new_n346));
  XNOR2_X1  g160(.A(G125), .B(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n202), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n335), .A2(new_n339), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(G146), .B1(new_n344), .B2(new_n345), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI211_X1 g168(.A(new_n351), .B(G146), .C1(new_n344), .C2(new_n345), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n317), .A2(new_n330), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(new_n320), .A3(new_n323), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n338), .A2(G110), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n350), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT77), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n350), .A2(new_n363), .A3(new_n360), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT22), .B(G137), .ZN(new_n365));
  INV_X1    g179(.A(G953), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n366), .A2(G221), .A3(G234), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n365), .B(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n362), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  AOI211_X1 g183(.A(new_n363), .B(new_n368), .C1(new_n350), .C2(new_n360), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT25), .B1(new_n372), .B2(new_n313), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n374));
  AOI211_X1 g188(.A(new_n374), .B(G902), .C1(new_n369), .C2(new_n371), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n314), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n372), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n314), .A2(G902), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT78), .B1(new_n311), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT32), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n292), .B1(new_n291), .B2(new_n267), .ZN(new_n385));
  NOR4_X1   g199(.A1(new_n300), .A2(KEYINPUT31), .A3(new_n277), .A4(new_n299), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n285), .B1(new_n280), .B2(new_n283), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n295), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n384), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n294), .A2(KEYINPUT32), .A3(new_n295), .ZN(new_n391));
  INV_X1    g205(.A(new_n310), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n364), .A2(new_n368), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n363), .B1(new_n350), .B2(new_n360), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n313), .B1(new_n397), .B2(new_n370), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n374), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n372), .A2(KEYINPUT25), .A3(new_n313), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n380), .B1(new_n401), .B2(new_n314), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n393), .A2(new_n394), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G221), .ZN(new_n404));
  XOR2_X1   g218(.A(KEYINPUT9), .B(G234), .Z(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n313), .ZN(new_n406));
  INV_X1    g220(.A(G469), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(new_n313), .ZN(new_n408));
  XOR2_X1   g222(.A(G110), .B(G140), .Z(new_n409));
  INV_X1    g223(.A(G227), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(G953), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n409), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n213), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n215), .B1(new_n417), .B2(new_n239), .ZN(new_n418));
  INV_X1    g232(.A(G101), .ZN(new_n419));
  INV_X1    g233(.A(G104), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G107), .ZN(new_n421));
  INV_X1    g235(.A(G107), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n422), .A2(KEYINPUT3), .A3(G104), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT3), .B1(new_n422), .B2(G104), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n419), .B(new_n421), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(G104), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n419), .B1(new_n421), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AND4_X1   g242(.A1(new_n416), .A2(new_n418), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n422), .A2(G104), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT3), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n420), .B2(G107), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n422), .A2(KEYINPUT3), .A3(G104), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n427), .B1(new_n434), .B2(new_n419), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n416), .B1(new_n435), .B2(new_n418), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n415), .B1(new_n429), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT4), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(KEYINPUT82), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n434), .A2(new_n419), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n434), .A2(new_n419), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n439), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n434), .B2(new_n419), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n251), .ZN(new_n446));
  INV_X1    g260(.A(new_n237), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n415), .B1(new_n212), .B2(new_n215), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n435), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n437), .A2(new_n446), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n445), .A2(new_n251), .B1(new_n435), .B2(new_n448), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n453), .A2(KEYINPUT84), .A3(new_n437), .A4(new_n447), .ZN(new_n454));
  OAI22_X1  g268(.A1(new_n429), .A2(new_n436), .B1(new_n271), .B2(new_n435), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(KEYINPUT12), .A3(new_n237), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n425), .A2(new_n428), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n459), .A2(G128), .B1(new_n203), .B2(new_n205), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n214), .A2(new_n203), .A3(new_n205), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT83), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n435), .A2(new_n416), .A3(new_n418), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n212), .A2(new_n215), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n463), .A2(new_n464), .B1(new_n465), .B2(new_n458), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n457), .B1(new_n466), .B2(new_n447), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n452), .A2(new_n454), .B1(new_n456), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n414), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n452), .A2(new_n454), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n453), .A2(new_n437), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n237), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n414), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n467), .A2(new_n456), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT81), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n470), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n408), .B1(new_n479), .B2(G469), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n466), .A2(new_n457), .A3(new_n447), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT12), .B1(new_n455), .B2(new_n237), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n467), .A2(KEYINPUT85), .A3(new_n456), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n471), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n475), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n471), .A2(new_n414), .A3(new_n473), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n487), .A2(new_n407), .A3(new_n313), .A4(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n406), .B1(new_n480), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G143), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n204), .A2(KEYINPUT92), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n492), .A2(new_n493), .A3(G214), .A4(new_n263), .ZN(new_n494));
  INV_X1    g308(.A(G237), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n366), .A3(G214), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n204), .A2(KEYINPUT92), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n494), .A2(G131), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT17), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n498), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n230), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(new_n499), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n501), .B(new_n505), .C1(new_n354), .C2(new_n355), .ZN(new_n506));
  XNOR2_X1  g320(.A(G113), .B(G122), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(new_n420), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n347), .B(new_n202), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n494), .A2(new_n498), .A3(KEYINPUT18), .A4(G131), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n510), .A2(new_n503), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n506), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT19), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n347), .B(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n346), .B1(new_n516), .B2(G146), .ZN(new_n517));
  AOI21_X1  g331(.A(G131), .B1(new_n494), .B2(new_n498), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n500), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n513), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n508), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  NOR2_X1   g338(.A1(G475), .A2(G902), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n525), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT20), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n523), .A2(KEYINPUT93), .A3(new_n524), .A4(new_n525), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n533));
  INV_X1    g347(.A(new_n514), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n508), .B1(new_n506), .B2(new_n513), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n313), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G475), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n532), .A2(new_n537), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT94), .ZN(new_n540));
  INV_X1    g354(.A(G478), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n196), .B2(G122), .ZN(new_n545));
  INV_X1    g359(.A(G122), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(KEYINPUT95), .A3(G116), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI221_X1 g362(.A(new_n548), .B1(KEYINPUT14), .B2(new_n422), .C1(G116), .C2(new_n546), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n209), .A2(G143), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT96), .B1(new_n213), .B2(G143), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n204), .A3(G128), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n216), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n216), .B1(new_n550), .B2(new_n554), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n549), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n422), .B1(new_n548), .B2(KEYINPUT14), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n545), .A2(new_n547), .B1(new_n196), .B2(G122), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n554), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT97), .B(KEYINPUT13), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT98), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n566), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n554), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n566), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n567), .A2(new_n570), .A3(new_n550), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G134), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n560), .A2(new_n422), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n560), .A2(new_n422), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n555), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n405), .A2(G217), .A3(new_n366), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n564), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n576), .B1(G134), .B2(new_n572), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n558), .A2(new_n563), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n543), .B1(new_n585), .B2(new_n313), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n313), .A3(new_n543), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(KEYINPUT99), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n590));
  AOI211_X1 g404(.A(G902), .B(new_n542), .C1(new_n581), .C2(new_n584), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n590), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(G952), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n594), .A2(KEYINPUT100), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(KEYINPUT100), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n366), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(G234), .A2(G237), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT21), .B(G898), .Z(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(G902), .A3(G953), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND4_X1   g417(.A1(new_n538), .A2(new_n540), .A3(new_n593), .A4(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(G214), .B1(G237), .B2(G902), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(G116), .B(G119), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT5), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n608), .B(G113), .C1(KEYINPUT5), .C2(new_n195), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n192), .A2(new_n607), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n435), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(G101), .A3(new_n443), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n425), .A2(new_n439), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n613), .B1(new_n614), .B2(new_n441), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n611), .B1(new_n615), .B2(new_n199), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT86), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT6), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT86), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n619), .B(new_n611), .C1(new_n615), .C2(new_n199), .ZN(new_n620));
  XNOR2_X1  g434(.A(G110), .B(G122), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n617), .A2(new_n618), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT88), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n621), .B1(new_n616), .B2(KEYINPUT86), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT88), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n625), .A2(new_n626), .A3(new_n618), .A4(new_n620), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n366), .A2(G224), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(G125), .B1(new_n243), .B2(new_n244), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n271), .A2(G125), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n465), .A2(new_n342), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n629), .A3(new_n631), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT89), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n617), .A2(new_n620), .A3(new_n622), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n611), .B(new_n621), .C1(new_n615), .C2(new_n199), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n640), .A2(KEYINPUT6), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT87), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n639), .A2(KEYINPUT87), .A3(new_n641), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n628), .B(new_n638), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT7), .ZN(new_n645));
  OAI22_X1  g459(.A1(new_n632), .A2(new_n633), .B1(new_n645), .B2(new_n630), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n635), .A2(KEYINPUT7), .A3(new_n629), .A4(new_n631), .ZN(new_n647));
  OAI21_X1  g461(.A(G113), .B1(new_n195), .B2(KEYINPUT5), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT90), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n608), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n650), .B1(new_n649), .B2(new_n608), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n458), .B1(new_n651), .B2(new_n610), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n609), .A2(new_n458), .A3(new_n610), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n621), .B(KEYINPUT8), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n646), .B(new_n647), .C1(new_n652), .C2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n640), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n313), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT91), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n644), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(G210), .B1(G237), .B2(G902), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n644), .A2(new_n659), .A3(new_n661), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n606), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n490), .A2(new_n604), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n383), .A2(new_n403), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G101), .ZN(G3));
  INV_X1    g482(.A(new_n406), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n479), .A2(G469), .ZN(new_n670));
  INV_X1    g484(.A(new_n408), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n489), .A3(new_n671), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n402), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n644), .A2(new_n661), .A3(new_n659), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n661), .B1(new_n644), .B2(new_n659), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n605), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n585), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT33), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT33), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n585), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n678), .A2(G478), .A3(new_n313), .A4(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n541), .B1(new_n677), .B2(G902), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n533), .B1(new_n532), .B2(new_n537), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n603), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n676), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n388), .A2(new_n389), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n298), .B1(new_n294), .B2(new_n313), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n673), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT34), .B(G104), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G6));
  XOR2_X1   g507(.A(new_n603), .B(KEYINPUT101), .Z(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n605), .B(new_n695), .C1(new_n674), .C2(new_n675), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n673), .A2(new_n690), .A3(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n589), .A2(new_n592), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n530), .A2(new_n526), .B1(new_n536), .B2(G475), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT35), .B(G107), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G9));
  INV_X1    g518(.A(new_n314), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n399), .B2(new_n400), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n368), .A2(KEYINPUT36), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT102), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n361), .B(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n379), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n706), .A2(KEYINPUT103), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n712));
  INV_X1    g526(.A(new_n710), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n712), .B1(new_n376), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n665), .A2(new_n669), .A3(new_n672), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n715), .A2(new_n716), .A3(new_n604), .A4(new_n690), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G110), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n717), .B(new_n719), .ZN(G12));
  OAI21_X1  g534(.A(new_n600), .B1(G900), .B2(new_n602), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n701), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n715), .A2(new_n716), .A3(new_n393), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G128), .ZN(G30));
  OAI21_X1  g539(.A(KEYINPUT103), .B1(new_n706), .B2(new_n710), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n376), .A2(new_n712), .A3(new_n713), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n593), .B1(new_n540), .B2(new_n538), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n605), .A3(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n721), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n490), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT40), .ZN(new_n734));
  INV_X1    g548(.A(new_n268), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n285), .B1(new_n262), .B2(new_n305), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n313), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G472), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n390), .A2(new_n391), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n674), .A2(new_n675), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT38), .ZN(new_n742));
  OR4_X1    g556(.A1(new_n730), .A2(new_n734), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G143), .ZN(G45));
  OAI211_X1 g558(.A(new_n683), .B(new_n721), .C1(new_n684), .C2(new_n685), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n715), .A2(new_n716), .A3(new_n393), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT106), .B(G146), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G48));
  NAND3_X1  g563(.A1(new_n487), .A2(new_n313), .A3(new_n488), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(G469), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n751), .A2(new_n669), .A3(new_n489), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n687), .A2(new_n393), .A3(new_n402), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  NAND4_X1  g569(.A1(new_n589), .A2(new_n592), .A3(new_n700), .A4(new_n695), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n706), .A2(new_n756), .A3(new_n380), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n393), .A2(new_n757), .A3(new_n665), .A4(new_n752), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n751), .A2(new_n489), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n676), .A2(new_n761), .A3(new_n406), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n762), .A2(new_n393), .A3(KEYINPUT107), .A4(new_n757), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G116), .ZN(G18));
  NAND4_X1  g579(.A1(new_n715), .A2(new_n393), .A3(new_n604), .A4(new_n762), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G119), .ZN(G21));
  NAND2_X1  g581(.A1(new_n294), .A2(new_n313), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n286), .B1(new_n306), .B2(new_n282), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n269), .A2(new_n293), .A3(new_n769), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n768), .A2(G472), .B1(new_n295), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n752), .A3(new_n402), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n665), .A2(new_n729), .A3(new_n695), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT108), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n770), .A2(new_n295), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n382), .A2(new_n775), .A3(new_n689), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n699), .B1(new_n684), .B2(new_n685), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n696), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n776), .A2(new_n778), .A3(new_n779), .A4(new_n752), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G122), .ZN(G24));
  NAND2_X1  g596(.A1(new_n745), .A2(KEYINPUT109), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n540), .A2(new_n538), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n785), .A3(new_n683), .A4(new_n721), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n715), .A2(new_n787), .A3(new_n762), .A4(new_n771), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G125), .ZN(G27));
  INV_X1    g603(.A(KEYINPUT42), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n390), .A2(new_n391), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n310), .B1(new_n791), .B2(KEYINPUT111), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n688), .B2(KEYINPUT32), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n382), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n783), .A2(new_n786), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n663), .A2(new_n605), .A3(new_n664), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT110), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n663), .A2(new_n799), .A3(new_n605), .A4(new_n664), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n490), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n790), .B1(new_n795), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n311), .A2(new_n382), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n798), .A2(new_n490), .A3(new_n800), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n805), .A3(new_n790), .A4(new_n787), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G131), .ZN(G33));
  NAND3_X1  g623(.A1(new_n804), .A2(new_n805), .A3(new_n723), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G134), .ZN(G36));
  NOR2_X1   g625(.A1(new_n684), .A2(new_n685), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n683), .ZN(new_n813));
  NAND2_X1  g627(.A1(KEYINPUT112), .A2(KEYINPUT43), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g629(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n817), .B(new_n715), .C1(new_n688), .C2(new_n689), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT44), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n798), .A2(new_n800), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n818), .B2(new_n819), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n479), .A2(KEYINPUT45), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n407), .B1(new_n479), .B2(KEYINPUT45), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n408), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n826), .A2(KEYINPUT46), .ZN(new_n827));
  INV_X1    g641(.A(new_n489), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n826), .B2(KEYINPUT46), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n406), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n820), .A2(new_n822), .A3(new_n732), .A4(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  XOR2_X1   g646(.A(new_n830), .B(KEYINPUT47), .Z(new_n833));
  NAND3_X1  g647(.A1(new_n311), .A2(new_n382), .A3(new_n746), .ZN(new_n834));
  OR3_X1    g648(.A1(new_n833), .A2(new_n821), .A3(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G140), .ZN(G42));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  INV_X1    g651(.A(new_n600), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n817), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n742), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n839), .A2(new_n840), .A3(new_n605), .A4(new_n772), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n821), .A2(new_n406), .A3(new_n761), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n402), .A2(new_n842), .A3(new_n838), .A4(new_n740), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n784), .A2(new_n683), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n837), .A2(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n771), .A2(new_n726), .A3(new_n727), .ZN(new_n846));
  INV_X1    g660(.A(new_n839), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n842), .ZN(new_n848));
  OAI221_X1 g662(.A(new_n845), .B1(new_n837), .B2(new_n841), .C1(new_n846), .C2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n751), .A2(new_n406), .A3(new_n489), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n833), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n847), .A2(new_n776), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n821), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT116), .Z(new_n854));
  AOI21_X1  g668(.A(new_n849), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT51), .Z(new_n856));
  AND3_X1   g670(.A1(new_n393), .A2(new_n394), .A3(new_n402), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n394), .B1(new_n393), .B2(new_n402), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n859), .A2(new_n666), .B1(new_n760), .B2(new_n763), .ZN(new_n860));
  INV_X1    g674(.A(new_n683), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n812), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n673), .A2(new_n862), .A3(new_n690), .A4(new_n697), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n717), .A2(new_n766), .A3(new_n863), .A4(new_n753), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n587), .A2(new_n588), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n812), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT115), .B1(new_n866), .B2(new_n696), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n673), .A2(new_n867), .A3(new_n690), .ZN(new_n868));
  OR3_X1    g682(.A1(new_n866), .A2(new_n696), .A3(KEYINPUT115), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n868), .A2(new_n869), .B1(new_n774), .B2(new_n780), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n860), .A2(new_n864), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n296), .A2(new_n297), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n392), .B(new_n794), .C1(new_n872), .C2(new_n793), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n402), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n805), .A2(new_n787), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT42), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n796), .A2(new_n846), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n700), .A2(new_n587), .A3(new_n588), .A4(new_n721), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n728), .A2(new_n311), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n805), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n876), .A2(new_n880), .A3(new_n806), .A4(new_n810), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n871), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n777), .A2(new_n676), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n706), .A2(new_n710), .A3(new_n722), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n739), .A3(new_n490), .A4(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n724), .A2(new_n788), .A3(new_n747), .A4(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n665), .A2(new_n726), .A3(new_n490), .A4(new_n727), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n889), .B(new_n393), .C1(new_n723), .C2(new_n746), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(KEYINPUT52), .A3(new_n788), .A4(new_n885), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n882), .A2(KEYINPUT53), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n847), .A2(new_n795), .A3(new_n842), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT48), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n852), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n597), .B1(new_n904), .B2(new_n762), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n843), .A2(new_n862), .ZN(new_n907));
  AND4_X1   g721(.A1(new_n903), .A2(new_n905), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n856), .A2(new_n900), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(G952), .B2(G953), .ZN(new_n910));
  NOR4_X1   g724(.A1(new_n813), .A2(new_n382), .A3(new_n606), .A4(new_n406), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT113), .Z(new_n912));
  XNOR2_X1  g726(.A(new_n761), .B(KEYINPUT49), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n912), .A2(new_n739), .A3(new_n840), .A4(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT114), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n910), .A2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n366), .A2(G952), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n313), .B1(new_n895), .B2(new_n896), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(G210), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n643), .A2(new_n642), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n624), .B2(new_n627), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(new_n638), .Z(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT55), .Z(new_n925));
  AOI21_X1  g739(.A(new_n917), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n918), .B(KEYINPUT117), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n662), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n925), .A2(KEYINPUT56), .ZN(new_n929));
  OAI211_X1 g743(.A(KEYINPUT118), .B(new_n926), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT118), .ZN(new_n931));
  INV_X1    g745(.A(new_n926), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n929), .B1(new_n927), .B2(new_n662), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(G51));
  XOR2_X1   g749(.A(new_n408), .B(KEYINPUT57), .Z(new_n936));
  OAI211_X1 g750(.A(new_n487), .B(new_n488), .C1(new_n900), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n927), .A2(new_n825), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n917), .B1(new_n937), .B2(new_n938), .ZN(G54));
  INV_X1    g753(.A(new_n917), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n927), .A2(KEYINPUT58), .A3(G475), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n523), .ZN(new_n942));
  AND4_X1   g756(.A1(KEYINPUT58), .A2(new_n927), .A3(G475), .A4(new_n523), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(G60));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n945));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT59), .Z(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n898), .B2(new_n899), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n678), .A2(new_n680), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n945), .B1(new_n952), .B2(new_n940), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n945), .B(new_n940), .C1(new_n949), .C2(new_n951), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n949), .A2(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n953), .A2(new_n956), .ZN(G63));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT120), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT60), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT53), .B1(new_n882), .B2(new_n892), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n805), .A2(new_n715), .A3(new_n771), .A4(new_n787), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n311), .A2(new_n878), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n805), .A3(new_n715), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n810), .A3(new_n964), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n965), .A2(new_n803), .A3(new_n807), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n869), .A2(new_n690), .A3(new_n673), .A4(new_n867), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n764), .A2(new_n781), .A3(new_n667), .A4(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n717), .A2(new_n766), .A3(new_n863), .A4(new_n753), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND4_X1   g784(.A1(KEYINPUT53), .A2(new_n966), .A3(new_n892), .A4(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n960), .B1(new_n961), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT121), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT121), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n974), .B(new_n960), .C1(new_n961), .C2(new_n971), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n709), .ZN(new_n977));
  AOI21_X1  g791(.A(KEYINPUT122), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n973), .A2(new_n377), .A3(new_n975), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n940), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT123), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n709), .B1(new_n973), .B2(new_n975), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(KEYINPUT122), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n981), .A2(new_n982), .A3(new_n983), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n982), .A2(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n940), .B(new_n979), .C1(new_n984), .C2(KEYINPUT122), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n984), .A2(KEYINPUT122), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n987), .B(new_n988), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n986), .A2(new_n991), .ZN(G66));
  AOI21_X1  g806(.A(new_n366), .B1(new_n601), .B2(G224), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n871), .B(KEYINPUT124), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(new_n366), .ZN(new_n995));
  INV_X1    g809(.A(G898), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n923), .B1(new_n996), .B2(G953), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT125), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n995), .B(new_n998), .ZN(G69));
  AND2_X1   g813(.A1(new_n890), .A2(new_n788), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n743), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT62), .Z(new_n1002));
  INV_X1    g816(.A(new_n862), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n733), .B(new_n821), .C1(new_n1003), .C2(new_n866), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n859), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT126), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1002), .A2(new_n831), .A3(new_n835), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n366), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n290), .B(new_n516), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(G900), .B2(G953), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n830), .A2(new_n732), .A3(new_n795), .A4(new_n883), .ZN(new_n1012));
  AND4_X1   g826(.A1(new_n808), .A2(new_n1012), .A3(new_n810), .A4(new_n1000), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n835), .A2(new_n831), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1011), .B1(new_n1014), .B2(G953), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n366), .B1(G227), .B2(G900), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n1009), .B2(KEYINPUT127), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1016), .B(new_n1018), .Z(G72));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT63), .Z(new_n1021));
  OAI21_X1  g835(.A(new_n1021), .B1(new_n1007), .B2(new_n994), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n1022), .B(new_n267), .C1(new_n277), .C2(new_n300), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1021), .B1(new_n1014), .B2(new_n994), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1024), .A2(new_n299), .A3(new_n291), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n268), .A2(new_n301), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n897), .A2(new_n1021), .A3(new_n1026), .ZN(new_n1027));
  AND4_X1   g841(.A1(new_n940), .A2(new_n1023), .A3(new_n1025), .A4(new_n1027), .ZN(G57));
endmodule


