//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT11), .B(G169gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  AND2_X1   g008(.A1(KEYINPUT85), .A2(G1gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT16), .B1(KEYINPUT85), .B2(G1gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n208), .B1(new_n212), .B2(KEYINPUT86), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(G1gat), .B2(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI221_X1 g014(.A(new_n212), .B1(KEYINPUT86), .B2(new_n208), .C1(G1gat), .C2(new_n209), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G29gat), .A2(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(G43gat), .A2(G50gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(G43gat), .A2(G50gat), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n227), .A3(KEYINPUT15), .ZN(new_n228));
  INV_X1    g027(.A(G50gat), .ZN(new_n229));
  AND2_X1   g028(.A1(KEYINPUT83), .A2(G43gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(KEYINPUT83), .A2(G43gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G43gat), .ZN(new_n233));
  AND2_X1   g032(.A1(KEYINPUT84), .A2(G50gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(KEYINPUT84), .A2(G50gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT15), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT15), .B1(new_n225), .B2(new_n226), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n238), .A2(new_n222), .A3(new_n220), .A4(new_n223), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n228), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n217), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G229gat), .A2(G233gat), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n242), .B(KEYINPUT13), .Z(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n240), .A2(KEYINPUT17), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT17), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n247), .B(new_n228), .C1(new_n237), .C2(new_n239), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n217), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n215), .A2(new_n216), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT87), .B1(new_n251), .B2(new_n240), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(new_n217), .A3(KEYINPUT87), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n253), .A2(new_n254), .B1(G229gat), .B2(G233gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n245), .B1(new_n255), .B2(KEYINPUT18), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n254), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n257), .A2(KEYINPUT18), .A3(new_n242), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n207), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n255), .A2(KEYINPUT18), .ZN(new_n260));
  INV_X1    g059(.A(new_n207), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(KEYINPUT18), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .A4(new_n245), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G141gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G148gat), .ZN(new_n270));
  INV_X1    g069(.A(G148gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G141gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT2), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n268), .A2(new_n276), .A3(new_n274), .ZN(new_n277));
  INV_X1    g076(.A(new_n266), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n274), .ZN(new_n280));
  INV_X1    g079(.A(new_n274), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT73), .B1(new_n281), .B2(new_n266), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n280), .A2(new_n282), .A3(new_n275), .A4(new_n273), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT1), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  XNOR2_X1  g088(.A(G127gat), .B(G134gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT67), .B(G113gat), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n288), .B(new_n290), .C1(new_n293), .C2(new_n287), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n285), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT4), .ZN(new_n298));
  NAND2_X1  g097(.A1(G225gat), .A2(G233gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n277), .A2(new_n283), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n277), .B2(new_n283), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT3), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n295), .B1(new_n284), .B2(KEYINPUT3), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n303), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(KEYINPUT3), .A3(new_n301), .ZN(new_n310));
  INV_X1    g109(.A(new_n307), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT75), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n298), .B(new_n299), .C1(new_n308), .C2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT5), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n309), .A2(new_n301), .A3(new_n295), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n297), .ZN(new_n316));
  INV_X1    g115(.A(new_n299), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n284), .A2(new_n295), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT4), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT75), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(KEYINPUT5), .A3(new_n299), .ZN(new_n326));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT0), .ZN(new_n328));
  XNOR2_X1  g127(.A(G57gat), .B(G85gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n328), .B(new_n329), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n320), .A2(new_n326), .A3(KEYINPUT6), .A4(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n320), .A2(new_n326), .A3(new_n331), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT6), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n331), .B1(new_n320), .B2(new_n326), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G64gat), .B(G92gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G197gat), .B(G204gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT22), .ZN(new_n343));
  INV_X1    g142(.A(G211gat), .ZN(new_n344));
  INV_X1    g143(.A(G218gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT70), .ZN(new_n348));
  XOR2_X1   g147(.A(G211gat), .B(G218gat), .Z(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n349), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT70), .A3(new_n347), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G226gat), .A2(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n357), .B1(new_n358), .B2(KEYINPUT24), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n359), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  OR2_X1    g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(KEYINPUT24), .A3(new_n358), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT25), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n360), .ZN(new_n368));
  INV_X1    g167(.A(new_n359), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n369), .A3(new_n366), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT27), .B(G183gat), .ZN(new_n373));
  INV_X1    g172(.A(G190gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(KEYINPUT65), .B(KEYINPUT28), .Z(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n373), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n358), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n361), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n357), .B1(new_n381), .B2(KEYINPUT26), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT66), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n383), .A2(KEYINPUT66), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n382), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI22_X1  g185(.A1(new_n367), .A2(new_n372), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n356), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n370), .B(new_n371), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n379), .A2(new_n358), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n385), .A2(new_n384), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n391), .B(new_n377), .C1(new_n392), .C2(new_n382), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n355), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n354), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n387), .A2(new_n356), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n390), .B2(new_n393), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n396), .B(new_n353), .C1(new_n397), .C2(new_n356), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n341), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n399), .A2(KEYINPUT71), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT30), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(KEYINPUT71), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n395), .A2(new_n398), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n404), .A2(new_n340), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n399), .B2(KEYINPUT30), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n337), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G22gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT31), .B(G50gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n285), .A2(new_n304), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n354), .B1(new_n414), .B2(new_n388), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT76), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n416), .B1(new_n353), .B2(KEYINPUT29), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n350), .A2(KEYINPUT76), .A3(new_n388), .A4(new_n352), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n304), .A3(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n302), .A2(new_n303), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n415), .B1(new_n421), .B2(KEYINPUT77), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT77), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n423), .A3(new_n420), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(G228gat), .ZN(new_n426));
  INV_X1    g225(.A(G233gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n415), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n351), .A2(new_n347), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n388), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n351), .A2(new_n347), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n304), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n428), .B1(new_n434), .B2(new_n284), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n413), .B1(new_n429), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n428), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n422), .B2(new_n424), .ZN(new_n439));
  INV_X1    g238(.A(new_n436), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n439), .A2(new_n440), .A3(new_n412), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n411), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n412), .B1(new_n439), .B2(new_n440), .ZN(new_n443));
  INV_X1    g242(.A(new_n424), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n423), .B1(new_n419), .B2(new_n420), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n444), .A2(new_n445), .A3(new_n415), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n436), .B(new_n413), .C1(new_n446), .C2(new_n438), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n447), .A3(new_n410), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n408), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n387), .A2(new_n296), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n390), .A2(new_n393), .A3(new_n295), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G227gat), .A2(G233gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT34), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n454), .B(KEYINPUT64), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(KEYINPUT34), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G15gat), .B(G43gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n451), .A2(new_n452), .A3(new_n457), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(KEYINPUT32), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT68), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n464), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n464), .B(KEYINPUT32), .C1(new_n467), .C2(new_n463), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n460), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n460), .A3(new_n471), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT36), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT69), .B1(new_n470), .B2(new_n471), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n476), .B1(new_n456), .B2(new_n459), .ZN(new_n477));
  AOI211_X1 g276(.A(KEYINPUT69), .B(new_n460), .C1(new_n470), .C2(new_n471), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n475), .B1(new_n479), .B2(KEYINPUT36), .ZN(new_n480));
  INV_X1    g279(.A(new_n448), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n410), .B1(new_n443), .B2(new_n447), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n313), .A2(new_n314), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n318), .B1(new_n325), .B2(new_n299), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n403), .A2(new_n406), .B1(new_n486), .B2(new_n331), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT39), .B1(new_n316), .B2(new_n317), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n298), .B1(new_n308), .B2(new_n312), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(new_n317), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT39), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n491), .A3(new_n317), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n330), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT78), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT78), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n495), .A3(new_n330), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n490), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n487), .B1(new_n497), .B2(KEYINPUT40), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  AOI211_X1 g298(.A(new_n499), .B(new_n490), .C1(new_n494), .C2(new_n496), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n483), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n330), .B1(new_n484), .B2(new_n485), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(new_n334), .A3(new_n333), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT80), .B1(new_n503), .B2(new_n332), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n395), .A2(KEYINPUT37), .A3(new_n398), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n505), .A2(new_n341), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT79), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n404), .B2(new_n508), .ZN(new_n509));
  AOI211_X1 g308(.A(KEYINPUT79), .B(KEYINPUT37), .C1(new_n395), .C2(new_n398), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT38), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT38), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n506), .B(new_n513), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n512), .A2(new_n400), .A3(new_n402), .A4(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n332), .A2(KEYINPUT80), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n504), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n450), .B(new_n480), .C1(new_n501), .C2(new_n517), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n442), .B(new_n448), .C1(new_n477), .C2(new_n478), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT35), .B1(new_n519), .B2(new_n408), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n516), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT81), .ZN(new_n522));
  INV_X1    g321(.A(new_n474), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(new_n472), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n473), .A2(KEYINPUT81), .A3(new_n474), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n403), .A2(new_n406), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n483), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n520), .B1(new_n521), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n265), .B1(new_n518), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT96), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT94), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT92), .ZN(new_n534));
  XOR2_X1   g333(.A(G99gat), .B(G106gat), .Z(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT91), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT8), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(G99gat), .B2(G106gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(G85gat), .A2(G92gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT8), .ZN(new_n543));
  OR2_X1    g342(.A1(G85gat), .A2(G92gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT91), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547));
  INV_X1    g346(.A(G85gat), .ZN(new_n548));
  INV_X1    g347(.A(G92gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n536), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n551), .ZN(new_n554));
  AOI211_X1 g353(.A(new_n535), .B(new_n554), .C1(new_n541), .C2(new_n545), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n534), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n543), .A2(KEYINPUT91), .A3(new_n544), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT91), .B1(new_n543), .B2(new_n544), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n552), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n535), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n552), .B(new_n536), .C1(new_n557), .C2(new_n558), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(KEYINPUT92), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n556), .A2(new_n240), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n560), .A2(KEYINPUT92), .A3(new_n561), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT92), .B1(new_n560), .B2(new_n561), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n249), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT93), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n556), .A2(new_n562), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(KEYINPUT93), .A3(new_n249), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n565), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n533), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT90), .ZN(new_n578));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n578), .B(new_n579), .Z(new_n580));
  AOI21_X1  g379(.A(new_n580), .B1(new_n573), .B2(new_n575), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n563), .A2(new_n564), .ZN(new_n582));
  AOI221_X4 g381(.A(new_n569), .B1(new_n246), .B2(new_n248), .C1(new_n556), .C2(new_n562), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT93), .B1(new_n571), .B2(new_n249), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(KEYINPUT94), .A3(new_n574), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n576), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT95), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n576), .A2(new_n581), .A3(new_n586), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n580), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n585), .A2(new_n574), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n582), .B(new_n575), .C1(new_n583), .C2(new_n584), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n532), .B1(new_n591), .B2(new_n596), .ZN(new_n597));
  AOI211_X1 g396(.A(KEYINPUT96), .B(new_n595), .C1(new_n588), .C2(new_n590), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT9), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(G57gat), .A2(G64gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(G57gat), .A2(G64gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT88), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(G71gat), .B2(G78gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G71gat), .B(G78gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n609), .A3(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G127gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n251), .B1(KEYINPUT21), .B2(new_n613), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT89), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G155gat), .ZN(new_n623));
  XOR2_X1   g422(.A(G183gat), .B(G211gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n620), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n599), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n613), .B1(new_n553), .B2(new_n555), .ZN(new_n631));
  INV_X1    g430(.A(G230gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n427), .ZN(new_n633));
  INV_X1    g432(.A(new_n612), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n609), .B1(new_n605), .B2(new_n607), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n636), .A2(new_n560), .A3(new_n561), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n631), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n639), .A2(KEYINPUT97), .ZN(new_n640));
  INV_X1    g439(.A(new_n633), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n556), .A2(new_n562), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT10), .B1(new_n631), .B2(new_n637), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n639), .A2(KEYINPUT97), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n640), .A2(new_n646), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n649), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n555), .A2(new_n553), .A3(new_n613), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n636), .B1(new_n561), .B2(new_n560), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n642), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n556), .A2(new_n562), .A3(new_n643), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n633), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n652), .B1(new_n657), .B2(new_n639), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n531), .A2(new_n630), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n337), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(G1gat), .Z(G1324gat));
  INV_X1    g462(.A(new_n661), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n208), .B1(new_n664), .B2(new_n527), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT16), .B(G8gat), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n661), .A2(new_n407), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT42), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(KEYINPUT42), .B2(new_n667), .ZN(G1325gat));
  OAI21_X1  g468(.A(G15gat), .B1(new_n661), .B2(new_n480), .ZN(new_n670));
  INV_X1    g469(.A(new_n526), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(G15gat), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n661), .B2(new_n672), .ZN(G1326gat));
  AND2_X1   g472(.A1(new_n531), .A2(new_n449), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n630), .A3(new_n660), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  NOR3_X1   g476(.A1(new_n573), .A2(new_n533), .A3(new_n575), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n594), .A2(new_n592), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n589), .B1(new_n680), .B2(new_n576), .ZN(new_n681));
  INV_X1    g480(.A(new_n590), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n596), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT96), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n591), .A2(new_n532), .A3(new_n596), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n518), .B2(new_n530), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n628), .A2(new_n659), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n264), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n691), .A2(G29gat), .A3(new_n337), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT45), .Z(new_n693));
  OAI21_X1  g492(.A(new_n480), .B1(new_n501), .B2(new_n517), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n450), .A2(KEYINPUT98), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n408), .A2(new_n449), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n530), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n699), .A2(new_n700), .A3(new_n599), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n687), .A2(new_n700), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n690), .ZN(new_n704));
  OAI21_X1  g503(.A(G29gat), .B1(new_n704), .B2(new_n337), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n693), .A2(new_n705), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n704), .B2(new_n407), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n701), .A2(new_n702), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n689), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(KEYINPUT101), .A3(new_n527), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n708), .A2(G36gat), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n527), .A2(new_n219), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n691), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT99), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(KEYINPUT100), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT100), .B(KEYINPUT46), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n712), .B(new_n717), .C1(new_n715), .C2(new_n718), .ZN(G1329gat));
  INV_X1    g518(.A(new_n480), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n710), .B(new_n720), .C1(new_n231), .C2(new_n230), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n230), .A2(new_n231), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n691), .B2(new_n671), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT47), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n721), .A2(new_n726), .A3(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1330gat));
  NOR2_X1   g527(.A1(new_n234), .A2(new_n235), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n710), .B2(new_n449), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n599), .A2(new_n688), .A3(new_n729), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n674), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OR3_X1    g533(.A1(new_n730), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n731), .B1(new_n730), .B2(new_n734), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1331gat));
  AND4_X1   g536(.A1(new_n265), .A2(new_n699), .A3(new_n630), .A4(new_n659), .ZN(new_n738));
  INV_X1    g537(.A(new_n337), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(KEYINPUT102), .B(G57gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1332gat));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n527), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT49), .B(G64gat), .Z(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n743), .B2(new_n745), .ZN(G1333gat));
  NAND2_X1  g545(.A1(new_n738), .A2(new_n720), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n671), .A2(G71gat), .ZN(new_n748));
  AOI22_X1  g547(.A1(new_n747), .A2(G71gat), .B1(new_n738), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g549(.A1(new_n738), .A2(new_n449), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g551(.A1(new_n628), .A2(new_n264), .A3(new_n660), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n703), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n739), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G85gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n628), .A2(new_n264), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n699), .A2(new_n599), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n699), .A2(KEYINPUT51), .A3(new_n599), .A4(new_n757), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT103), .Z(new_n763));
  NAND3_X1  g562(.A1(new_n739), .A2(new_n548), .A3(new_n659), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n756), .B1(new_n763), .B2(new_n764), .ZN(G1336gat));
  NAND3_X1  g564(.A1(new_n760), .A2(KEYINPUT104), .A3(new_n761), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n758), .A2(new_n767), .A3(new_n759), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n407), .A2(G92gat), .A3(new_n660), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT105), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT105), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n766), .A2(new_n772), .A3(new_n768), .A4(new_n769), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n527), .B(new_n753), .C1(new_n701), .C2(new_n702), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n771), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT52), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  INV_X1    g577(.A(new_n769), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n775), .B(new_n778), .C1(new_n762), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(G1337gat));
  NAND2_X1  g580(.A1(new_n754), .A2(new_n720), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT106), .B(G99gat), .Z(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n671), .A2(new_n660), .A3(new_n783), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT107), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n763), .B2(new_n786), .ZN(G1338gat));
  NOR3_X1   g586(.A1(new_n483), .A2(G106gat), .A3(new_n660), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n766), .A2(new_n768), .A3(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n449), .B(new_n753), .C1(new_n701), .C2(new_n702), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(G106gat), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT53), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  INV_X1    g592(.A(new_n788), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n762), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n792), .B1(new_n791), .B2(new_n795), .ZN(G1339gat));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n655), .A2(new_n633), .A3(new_n656), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n646), .A2(new_n798), .A3(KEYINPUT54), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n652), .B1(new_n646), .B2(KEYINPUT54), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n649), .B1(new_n657), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n646), .A2(new_n798), .A3(KEYINPUT54), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT55), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n801), .A2(new_n651), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n801), .A2(KEYINPUT108), .A3(new_n651), .A4(new_n805), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n264), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n241), .A2(new_n244), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n257), .B2(new_n242), .ZN(new_n812));
  INV_X1    g611(.A(new_n205), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n263), .A2(new_n659), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n598), .B2(new_n597), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n263), .A2(new_n814), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n808), .A2(new_n818), .A3(new_n809), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n684), .A2(new_n820), .A3(new_n685), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n628), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  NOR4_X1   g621(.A1(new_n599), .A2(new_n629), .A3(new_n264), .A4(new_n659), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(new_n449), .A3(new_n671), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n337), .A2(new_n527), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n265), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n684), .A2(new_n685), .B1(new_n815), .B2(new_n810), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n597), .A2(new_n598), .A3(new_n819), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n629), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n686), .A2(new_n265), .A3(new_n628), .A4(new_n660), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n337), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n519), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n527), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n264), .A2(new_n293), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT109), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n828), .A2(new_n839), .ZN(G1340gat));
  OAI21_X1  g639(.A(G120gat), .B1(new_n827), .B2(new_n660), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n287), .A3(new_n659), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT110), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n827), .B2(new_n629), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n836), .A2(new_n617), .A3(new_n628), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1342gat));
  NOR2_X1   g646(.A1(new_n686), .A2(new_n527), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OR3_X1    g648(.A1(new_n835), .A2(G134gat), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT111), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n825), .A2(new_n599), .A3(new_n826), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n850), .A2(KEYINPUT56), .B1(new_n853), .B2(G134gat), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1343gat));
  XNOR2_X1  g654(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n739), .B1(new_n822), .B2(new_n823), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n480), .A2(new_n449), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT115), .B(new_n739), .C1(new_n822), .C2(new_n823), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n861), .A2(new_n407), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n265), .A2(G141gat), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n858), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n803), .A2(new_n804), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n640), .A2(new_n649), .A3(new_n650), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n869), .A2(new_n797), .B1(new_n870), .B2(new_n646), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n264), .A2(new_n805), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n815), .A2(KEYINPUT112), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT112), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n263), .A2(new_n874), .A3(new_n659), .A4(new_n814), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n597), .B2(new_n598), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT113), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT113), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n876), .B(new_n879), .C1(new_n597), .C2(new_n598), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n821), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n823), .B1(new_n881), .B2(new_n629), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n483), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT114), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n877), .A2(KEYINPUT113), .B1(new_n599), .B2(new_n820), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n628), .B1(new_n888), .B2(new_n880), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n887), .B(new_n884), .C1(new_n889), .C2(new_n823), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n883), .B1(new_n824), .B2(new_n483), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n480), .A2(new_n826), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n264), .A3(new_n893), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n857), .B(new_n868), .C1(G141gat), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(G141gat), .ZN(new_n896));
  INV_X1    g695(.A(new_n868), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n856), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n895), .A2(new_n898), .ZN(G1344gat));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n892), .A2(new_n893), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n900), .B(G148gat), .C1(new_n901), .C2(new_n660), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n818), .A2(new_n805), .A3(new_n871), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n599), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n877), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n628), .B1(new_n905), .B2(KEYINPUT119), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n907), .A3(new_n877), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n823), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n883), .B1(new_n909), .B2(new_n483), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n831), .A2(new_n832), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n884), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n893), .A2(new_n659), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n271), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n902), .B1(new_n900), .B2(new_n915), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n865), .A2(G148gat), .A3(new_n660), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n917), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(G1345gat));
  NAND4_X1  g719(.A1(new_n892), .A2(G155gat), .A3(new_n628), .A4(new_n893), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n862), .B1(new_n833), .B2(KEYINPUT115), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n922), .A2(new_n407), .A3(new_n628), .A4(new_n861), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(KEYINPUT120), .ZN(new_n924));
  INV_X1    g723(.A(G155gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n923), .B2(KEYINPUT120), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n921), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(KEYINPUT121), .B(new_n921), .C1(new_n924), .C2(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1346gat));
  OAI21_X1  g730(.A(G162gat), .B1(new_n901), .B2(new_n686), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n849), .A2(G162gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n922), .A2(new_n861), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT122), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n739), .A2(new_n407), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT123), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n825), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(G169gat), .B1(new_n939), .B2(new_n265), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT124), .Z(new_n941));
  AND2_X1   g740(.A1(new_n911), .A2(new_n937), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n834), .ZN(new_n943));
  OR3_X1    g742(.A1(new_n943), .A2(G169gat), .A3(new_n265), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n941), .A2(new_n944), .ZN(G1348gat));
  INV_X1    g744(.A(G176gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n946), .B1(new_n943), .B2(new_n660), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT125), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n939), .A2(new_n946), .A3(new_n660), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(G1349gat));
  OAI21_X1  g749(.A(G183gat), .B1(new_n939), .B2(new_n629), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n628), .A2(new_n373), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n943), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g753(.A(G190gat), .B1(new_n939), .B2(new_n686), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n599), .A2(new_n374), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n943), .B2(new_n957), .ZN(G1351gat));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n863), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n264), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n938), .A2(new_n480), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n962), .B1(new_n910), .B2(new_n912), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n264), .A2(G197gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  AOI21_X1  g764(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n960), .A2(new_n659), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n967), .B(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(G204gat), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n963), .A2(new_n659), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n960), .A2(new_n344), .A3(new_n628), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n974));
  AOI211_X1 g773(.A(new_n974), .B(new_n344), .C1(new_n963), .C2(new_n628), .ZN(new_n975));
  INV_X1    g774(.A(new_n962), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n913), .A2(new_n628), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n977), .B2(G211gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n973), .B1(new_n975), .B2(new_n978), .ZN(G1354gat));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n599), .B1(new_n963), .B2(new_n980), .ZN(new_n981));
  AOI211_X1 g780(.A(KEYINPUT127), .B(new_n962), .C1(new_n910), .C2(new_n912), .ZN(new_n982));
  OAI21_X1  g781(.A(G218gat), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n960), .A2(new_n345), .A3(new_n599), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1355gat));
endmodule


