//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT68), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT70), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT69), .B(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G137), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n465), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OAI221_X1 g051(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n465), .C2(G112), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n474), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  OR3_X1    g056(.A1(new_n480), .A2(KEYINPUT71), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT71), .B1(new_n480), .B2(new_n481), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n478), .B1(new_n482), .B2(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(new_n460), .A2(KEYINPUT69), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n485), .B(new_n487), .C1(new_n472), .C2(new_n473), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT4), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n464), .A2(new_n465), .A3(new_n491), .A4(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n472), .B2(new_n473), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n464), .A2(KEYINPUT72), .A3(new_n497), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(G50), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT73), .B(G88), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT74), .ZN(new_n515));
  XOR2_X1   g090(.A(KEYINPUT6), .B(G651), .Z(new_n516));
  XOR2_X1   g091(.A(KEYINPUT73), .B(G88), .Z(new_n517));
  NAND2_X1  g092(.A1(new_n508), .A2(new_n509), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n516), .B1(new_n519), .B2(new_n505), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n515), .A2(new_n522), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT76), .B(G89), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n513), .A2(new_n530), .B1(G63), .B2(G651), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n531), .B2(new_n510), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n516), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n513), .A2(KEYINPUT75), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n534), .A2(G543), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n532), .B1(G51), .B2(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(new_n536), .A2(G52), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n524), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n510), .A2(new_n516), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT77), .B(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n538), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(new_n536), .A2(G43), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n524), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n541), .A2(G81), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT78), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n510), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n541), .A2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n534), .A2(G53), .A3(G543), .A4(new_n535), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G299));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n544), .B(new_n569), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  NAND4_X1  g146(.A1(new_n534), .A2(G49), .A3(G543), .A4(new_n535), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n541), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n508), .B2(new_n509), .ZN(new_n577));
  AND2_X1   g152(.A1(G73), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n508), .B2(new_n509), .ZN(new_n583));
  AND2_X1   g158(.A1(G48), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n513), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n579), .A2(new_n580), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n541), .A2(G85), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n534), .A2(G543), .A3(new_n535), .ZN(new_n592));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n590), .B1(new_n524), .B2(new_n591), .C1(new_n592), .C2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(new_n541), .A2(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n536), .A2(G54), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n518), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n524), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n544), .B(KEYINPUT79), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G284));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n567), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n567), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(new_n601), .ZN(new_n609));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G860), .ZN(G148));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n550), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n601), .A2(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g191(.A1(new_n460), .A2(G2104), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n464), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(G123), .A2(new_n475), .B1(new_n479), .B2(G135), .ZN(new_n623));
  OAI221_X1 g198(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n465), .C2(G111), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT81), .B(G2096), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n622), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(KEYINPUT83), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(KEYINPUT83), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n639), .B(new_n640), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n637), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n637), .B2(new_n638), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n630), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n637), .A2(new_n638), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(new_n641), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n637), .A2(new_n638), .A3(new_n642), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n629), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n645), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g228(.A1(new_n645), .A2(new_n649), .A3(KEYINPUT84), .A4(new_n650), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT85), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n650), .B1(new_n645), .B2(new_n649), .ZN(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n656), .B1(new_n655), .B2(new_n659), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(G401));
  INV_X1    g237(.A(KEYINPUT18), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n621), .ZN(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(G2096), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n677), .A2(new_n682), .A3(new_n680), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n682), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n685));
  AOI211_X1 g260(.A(new_n681), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n684), .B2(new_n685), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G1971), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G6), .B(G305), .S(G16), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT32), .B(G1981), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  AND2_X1   g276(.A1(new_n694), .A2(G23), .ZN(new_n702));
  NAND2_X1  g277(.A1(G288), .A2(KEYINPUT89), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT89), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n572), .A2(new_n573), .A3(new_n704), .A4(new_n574), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n702), .B1(new_n706), .B2(G16), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT33), .B(G1976), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n708), .ZN(new_n711));
  AND3_X1   g286(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n710), .B1(new_n709), .B2(new_n711), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n698), .B(new_n701), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  OAI221_X1 g295(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n465), .C2(G107), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT87), .ZN(new_n722));
  AOI22_X1  g297(.A1(G119), .A2(new_n475), .B1(new_n479), .B2(G131), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n720), .B1(new_n725), .B2(new_n719), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G24), .B(G290), .S(G16), .Z(new_n730));
  XOR2_X1   g305(.A(KEYINPUT88), .B(G1986), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(KEYINPUT91), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n718), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT91), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(KEYINPUT36), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n736), .A2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n694), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT103), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT23), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n567), .B2(new_n694), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT104), .ZN(new_n745));
  INV_X1    g320(.A(G1956), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(G2090), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n719), .A2(G35), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n719), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT29), .Z(new_n752));
  OAI211_X1 g327(.A(new_n747), .B(new_n748), .C1(new_n749), .C2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT105), .ZN(new_n754));
  NOR2_X1   g329(.A1(G168), .A2(new_n694), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n694), .B2(G21), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT98), .ZN(new_n759));
  NOR2_X1   g334(.A1(G5), .A2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT99), .Z(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n544), .B2(new_n694), .ZN(new_n762));
  INV_X1    g337(.A(G1961), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT100), .Z(new_n765));
  NAND3_X1  g340(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT95), .B(KEYINPUT25), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(new_n465), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n479), .A2(G139), .ZN(new_n771));
  AND3_X1   g346(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G29), .B2(G33), .ZN(new_n774));
  INV_X1    g349(.A(G2072), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n763), .B2(new_n762), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n757), .A2(new_n756), .B1(new_n774), .B2(new_n775), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n759), .A2(new_n765), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT26), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n475), .B2(G129), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n479), .A2(G141), .B1(G105), .B2(new_n617), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT96), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  MUX2_X1   g364(.A(G32), .B(new_n789), .S(G29), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT27), .B(G1996), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT97), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n790), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n719), .A2(G27), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G164), .B2(new_n719), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT101), .B(G2078), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G34), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n798), .A2(KEYINPUT24), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(KEYINPUT24), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n719), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G160), .B2(new_n719), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2084), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT30), .B(G28), .ZN(new_n804));
  OR2_X1    g379(.A1(KEYINPUT31), .A2(G11), .ZN(new_n805));
  NAND2_X1  g380(.A1(KEYINPUT31), .A2(G11), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n804), .A2(new_n719), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n625), .B2(new_n719), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n793), .A2(new_n797), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n779), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT102), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n475), .A2(G128), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT92), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n479), .A2(G140), .ZN(new_n816));
  NOR2_X1   g391(.A1(G104), .A2(G2105), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT93), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n719), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT94), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n719), .A2(G26), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT28), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G2067), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n694), .A2(G19), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n551), .B2(new_n694), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1341), .ZN(new_n831));
  INV_X1    g406(.A(G1348), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n609), .A2(G16), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G4), .B2(G16), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n831), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n752), .A2(new_n749), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n834), .A2(new_n832), .ZN(new_n837));
  AND4_X1   g412(.A1(new_n828), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n811), .A2(KEYINPUT102), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n754), .A2(new_n812), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n739), .A2(new_n740), .A3(new_n840), .ZN(G311));
  NOR2_X1   g416(.A1(new_n740), .A2(new_n840), .ZN(new_n842));
  INV_X1    g417(.A(new_n739), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(G150));
  AOI22_X1  g419(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(new_n524), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT106), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n541), .A2(G93), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G55), .ZN(new_n851));
  OAI22_X1  g426(.A1(new_n846), .A2(new_n847), .B1(new_n592), .B2(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n853), .A2(KEYINPUT107), .A3(new_n550), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n550), .A2(KEYINPUT107), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT107), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n546), .A2(new_n856), .A3(new_n548), .A4(new_n549), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n850), .A2(new_n852), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n601), .A2(new_n610), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  INV_X1    g439(.A(G860), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n858), .A2(new_n865), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  XOR2_X1   g445(.A(new_n625), .B(G160), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G162), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n821), .A2(new_n503), .ZN(new_n873));
  OAI21_X1  g448(.A(G164), .B1(new_n815), .B2(new_n820), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n475), .A2(G130), .ZN(new_n876));
  OAI221_X1 g451(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n465), .C2(G118), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n479), .A2(G142), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n873), .A2(new_n879), .A3(new_n874), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n722), .A2(KEYINPUT109), .A3(new_n723), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT109), .B1(new_n722), .B2(new_n723), .ZN(new_n885));
  OR3_X1    g460(.A1(new_n884), .A2(new_n885), .A3(new_n619), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n619), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n881), .A2(new_n887), .A3(new_n886), .A4(new_n882), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n786), .A2(KEYINPUT108), .A3(new_n788), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT108), .B1(new_n786), .B2(new_n788), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n772), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n785), .B2(new_n772), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n889), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n889), .B2(new_n890), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n872), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT110), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g474(.A(KEYINPUT110), .B(new_n872), .C1(new_n895), .C2(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n895), .A2(new_n896), .A3(new_n872), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n902), .A2(G37), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(KEYINPUT111), .B(KEYINPUT40), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(G395));
  XNOR2_X1  g481(.A(G299), .B(new_n601), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT41), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n860), .B(new_n614), .Z(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT42), .ZN(new_n913));
  INV_X1    g488(.A(new_n706), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n914), .A2(G290), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(G290), .ZN(new_n916));
  XNOR2_X1  g491(.A(G305), .B(G303), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n915), .B2(new_n916), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n910), .A2(new_n921), .A3(new_n911), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n913), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n920), .B1(new_n913), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n853), .A2(new_n612), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(G295));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n926), .ZN(G331));
  INV_X1    g503(.A(G37), .ZN(new_n929));
  NAND2_X1  g504(.A1(G286), .A2(new_n544), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(G301), .B2(G286), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n860), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n603), .A2(G168), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(new_n854), .A3(new_n859), .A4(new_n930), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n601), .B(new_n567), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n931), .A2(KEYINPUT112), .A3(new_n860), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT112), .B1(new_n931), .B2(new_n860), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n937), .B1(new_n940), .B2(new_n908), .ZN(new_n941));
  INV_X1    g516(.A(new_n920), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n929), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI211_X1 g518(.A(new_n920), .B(new_n937), .C1(new_n940), .C2(new_n908), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT43), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n942), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n935), .B(KEYINPUT41), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n934), .B2(new_n932), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n934), .A2(new_n935), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n932), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n931), .A2(KEYINPUT112), .A3(new_n860), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n920), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n946), .A2(new_n954), .A3(new_n955), .A4(new_n929), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n945), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AND4_X1   g534(.A1(KEYINPUT43), .A2(new_n946), .A3(new_n929), .A4(new_n954), .ZN(new_n960));
  INV_X1    g535(.A(new_n934), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n951), .B2(new_n952), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n936), .B1(new_n962), .B2(new_n947), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n963), .B2(new_n920), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT43), .B1(new_n964), .B2(new_n946), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n959), .A2(new_n966), .ZN(G397));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(G1384), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n503), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n465), .ZN(new_n971));
  INV_X1    g546(.A(G125), .ZN(new_n972));
  INV_X1    g547(.A(new_n472), .ZN(new_n973));
  INV_X1    g548(.A(new_n473), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n469), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n977), .A2(new_n463), .A3(G40), .A4(new_n466), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n970), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n493), .B2(new_n502), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n981), .A2(KEYINPUT45), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n757), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT119), .ZN(new_n984));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n503), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n987));
  INV_X1    g562(.A(G2084), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n981), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n987), .A2(new_n988), .A3(new_n979), .A4(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT119), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n992), .B(new_n757), .C1(new_n980), .C2(new_n982), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n984), .A2(G168), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n995), .B1(KEYINPUT124), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(KEYINPUT124), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n994), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n984), .A2(new_n991), .A3(new_n993), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(G8), .A3(G286), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n999), .B1(new_n994), .B2(new_n997), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT125), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n994), .A2(new_n997), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n998), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT125), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n1002), .A4(new_n1000), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT62), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1005), .A2(new_n1012), .A3(new_n1009), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G303), .A2(G8), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1016), .A2(KEYINPUT116), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT116), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n980), .B2(new_n982), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n986), .A2(new_n968), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n978), .B1(new_n503), .B2(new_n969), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(KEYINPUT114), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n697), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n990), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n979), .B1(new_n981), .B2(new_n989), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(KEYINPUT115), .A3(new_n749), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n987), .A2(new_n749), .A3(new_n979), .A4(new_n990), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1026), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1020), .A2(new_n1034), .A3(G8), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  INV_X1    g611(.A(G1981), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n586), .B2(new_n588), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n581), .A2(new_n585), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1039), .A2(G1981), .A3(new_n587), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1036), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n995), .B1(new_n979), .B2(new_n981), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n586), .A2(new_n1037), .A3(new_n588), .ZN(new_n1043));
  OAI21_X1  g618(.A(G1981), .B1(new_n1039), .B2(new_n587), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n703), .A2(G1976), .A3(new_n705), .ZN(new_n1047));
  INV_X1    g622(.A(G1976), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT52), .B1(G288), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1042), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1042), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT52), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT117), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(new_n1055), .A3(KEYINPUT52), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1051), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1035), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1017), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1062), .B2(new_n995), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n987), .A2(new_n979), .A3(new_n990), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n980), .A2(new_n982), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(G2078), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1064), .A2(new_n763), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(G2078), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(new_n1069), .B2(KEYINPUT53), .ZN(new_n1070));
  AND4_X1   g645(.A1(new_n603), .A2(new_n1058), .A3(new_n1063), .A4(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1011), .A2(new_n1013), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1064), .A2(new_n832), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n979), .A2(new_n981), .A3(new_n827), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(KEYINPUT60), .A3(new_n1074), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n609), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n563), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n567), .B(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1064), .A2(new_n746), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1065), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1083), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1079), .B1(new_n1090), .B2(KEYINPUT61), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT58), .B(G1341), .Z(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n986), .B2(new_n978), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(G1996), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n551), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT59), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1083), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(KEYINPUT61), .A3(new_n1087), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1078), .A2(new_n609), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1097), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n601), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1100), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT123), .B1(new_n1106), .B2(new_n1087), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT123), .B(new_n1087), .C1(new_n1089), .C2(new_n1104), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n1091), .A2(new_n1103), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1070), .A2(new_n603), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1068), .B(G301), .C1(new_n1069), .C2(KEYINPUT53), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT54), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1070), .A2(G171), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1112), .A2(KEYINPUT54), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1110), .A2(new_n1116), .A3(new_n1010), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n993), .A2(new_n991), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n992), .B1(new_n1094), .B2(new_n757), .ZN(new_n1121));
  OAI211_X1 g696(.A(G8), .B(G168), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1063), .A2(new_n1035), .A3(new_n1057), .A4(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1061), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n1034), .B2(G8), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1001), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1124), .A2(new_n1125), .B1(new_n1058), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1035), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1057), .ZN(new_n1132));
  INV_X1    g707(.A(G288), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1046), .A2(new_n1048), .A3(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1040), .B(KEYINPUT118), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1042), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1132), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1119), .B1(new_n1130), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1058), .A2(new_n1129), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1138), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(KEYINPUT121), .A3(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1072), .A2(new_n1118), .A3(new_n1139), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n982), .A2(new_n979), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1147), .A2(G1996), .A3(new_n784), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT113), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n821), .B(G2067), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(G1996), .B2(new_n789), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1149), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n725), .A2(new_n727), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n725), .A2(new_n727), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1147), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G290), .B(G1986), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n1147), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1145), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1146), .B1(new_n1150), .B2(new_n785), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT46), .B1(new_n1146), .B2(G1996), .ZN(new_n1161));
  OR3_X1    g736(.A1(new_n1146), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1164));
  XNOR2_X1  g739(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n821), .A2(new_n827), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1146), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1156), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1146), .A2(G1986), .A3(G290), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT48), .Z(new_n1171));
  AOI211_X1 g746(.A(new_n1165), .B(new_n1168), .C1(new_n1169), .C2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1159), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g748(.A1(G227), .A2(new_n458), .ZN(new_n1175));
  OAI21_X1  g749(.A(new_n1175), .B1(new_n660), .B2(new_n661), .ZN(new_n1176));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1177));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g752(.A(KEYINPUT127), .B(new_n1175), .C1(new_n660), .C2(new_n661), .ZN(new_n1179));
  AOI21_X1  g753(.A(G229), .B1(new_n901), .B2(new_n903), .ZN(new_n1180));
  AND4_X1   g754(.A1(new_n957), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(G308));
  NAND4_X1  g755(.A1(new_n957), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(G225));
endmodule


