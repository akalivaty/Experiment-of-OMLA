//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT65), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G137), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n469), .B(KEYINPUT67), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n459), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n472), .A3(G125), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n468), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n467), .A2(new_n474), .ZN(G160));
  AND2_X1   g050(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(new_n468), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n471), .A2(new_n472), .A3(G138), .A4(new_n468), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n464), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g068(.A1(KEYINPUT70), .A2(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT70), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2105), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n489), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n502), .B1(new_n510), .B2(G651), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  AOI211_X1 g087(.A(KEYINPUT72), .B(new_n512), .C1(new_n508), .C2(new_n509), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n514), .B1(new_n512), .B2(KEYINPUT71), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT6), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(G50), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n507), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR3_X1   g097(.A1(new_n511), .A2(new_n513), .A3(new_n522), .ZN(G166));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n516), .A2(KEYINPUT6), .A3(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(KEYINPUT6), .B1(new_n516), .B2(G651), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n515), .A2(KEYINPUT73), .A3(new_n517), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n530), .A2(G543), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n525), .B(new_n526), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n515), .A2(new_n517), .B1(new_n505), .B2(new_n506), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n535), .A2(G89), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n504), .B1(new_n518), .B2(new_n527), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n541), .A2(G51), .A3(new_n531), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n525), .B1(new_n542), .B2(new_n526), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n524), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n526), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n546), .A2(KEYINPUT75), .A3(new_n534), .A4(new_n539), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(G168));
  XNOR2_X1  g123(.A(KEYINPUT76), .B(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n535), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  OAI221_X1 g127(.A(new_n550), .B1(new_n512), .B2(new_n551), .C1(new_n532), .C2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND3_X1  g129(.A1(new_n541), .A2(G43), .A3(new_n531), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT5), .B(G543), .Z(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n535), .A2(G81), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n555), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(KEYINPUT77), .B2(KEYINPUT9), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n530), .A2(G543), .A3(new_n531), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n557), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G91), .B2(new_n535), .ZN(new_n577));
  INV_X1    g152(.A(new_n572), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n541), .A2(new_n531), .A3(new_n578), .A4(new_n570), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n573), .A2(new_n577), .A3(new_n579), .ZN(G299));
  AND2_X1   g155(.A1(new_n544), .A2(new_n547), .ZN(G286));
  OR3_X1    g156(.A1(new_n511), .A2(new_n513), .A3(new_n522), .ZN(G303));
  NAND2_X1  g157(.A1(new_n535), .A2(G87), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n532), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n541), .A2(KEYINPUT78), .A3(G49), .A4(new_n531), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G288));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n505), .B2(new_n506), .ZN(new_n593));
  AND2_X1   g168(.A1(G73), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n518), .A2(G48), .A3(G543), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n518), .A2(G86), .A3(new_n507), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n595), .A2(KEYINPUT79), .A3(new_n596), .A4(new_n597), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(G305));
  NAND2_X1  g178(.A1(new_n535), .A2(G85), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G47), .ZN(new_n606));
  OAI221_X1 g181(.A(new_n604), .B1(new_n512), .B2(new_n605), .C1(new_n532), .C2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n532), .A2(KEYINPUT81), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n541), .A2(new_n610), .A3(new_n531), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n609), .A2(G54), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n614));
  AND4_X1   g189(.A1(new_n614), .A2(new_n518), .A3(G92), .A4(new_n507), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n535), .B2(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(new_n512), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n518), .A2(G92), .A3(new_n507), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT80), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n535), .A2(new_n614), .A3(G92), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n621), .A2(KEYINPUT10), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g198(.A1(new_n612), .A2(new_n617), .A3(new_n619), .A4(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n608), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n608), .B1(new_n625), .B2(G868), .ZN(G321));
  NOR2_X1   g202(.A1(G299), .A2(G868), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g204(.A(new_n628), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n625), .B1(new_n631), .B2(G860), .ZN(G148));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n562), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n624), .A2(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n633), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n479), .A2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n481), .A2(G123), .ZN(new_n639));
  OR2_X1    g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n640), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n642), .A2(G2096), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(G2096), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT12), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2100), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n643), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT82), .Z(G156));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT84), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2430), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(G14), .B1(new_n661), .B2(new_n664), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(G401));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT17), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT86), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n671), .B1(new_n672), .B2(new_n668), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(KEYINPUT85), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(KEYINPUT85), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n669), .A2(new_n672), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n670), .A2(new_n672), .A3(new_n668), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT18), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n674), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2096), .B(G2100), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(KEYINPUT87), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(KEYINPUT87), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  OR3_X1    g264(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n687), .B2(new_n688), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(KEYINPUT89), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(KEYINPUT89), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n690), .A2(new_n695), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n691), .A2(new_n695), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT88), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n697), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G1991), .B(G1996), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n706), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n705), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n708), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n709), .A2(new_n713), .ZN(G229));
  XOR2_X1   g289(.A(KEYINPUT100), .B(G28), .Z(new_n715));
  AOI21_X1  g290(.A(G29), .B1(new_n715), .B2(KEYINPUT30), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(KEYINPUT30), .B2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT31), .B(G11), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(G164), .A2(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G27), .B2(G29), .ZN(new_n721));
  INV_X1    g296(.A(G2078), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n724), .A2(G5), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G301), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1961), .ZN(new_n727));
  OAI221_X1 g302(.A(new_n723), .B1(new_n722), .B2(new_n721), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n724), .A2(G19), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n563), .B2(new_n724), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(G1341), .Z(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  AND2_X1   g307(.A1(KEYINPUT24), .A2(G34), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(KEYINPUT24), .B2(G34), .ZN(new_n734));
  OAI22_X1  g309(.A1(G160), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(G2084), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(G2084), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n642), .A2(new_n732), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n731), .A2(new_n736), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n728), .B(new_n739), .C1(new_n727), .C2(new_n726), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n732), .A2(G26), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT28), .Z(new_n742));
  INV_X1    g317(.A(KEYINPUT96), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n476), .A2(new_n477), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(new_n468), .ZN(new_n745));
  INV_X1    g320(.A(G140), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n479), .A2(KEYINPUT96), .A3(G140), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G116), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n481), .B2(G128), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n742), .B1(new_n754), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G2067), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n740), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n479), .A2(G141), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n481), .A2(G129), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT26), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  AND2_X1   g338(.A1(G105), .A2(G2104), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n762), .A2(new_n763), .B1(new_n468), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n758), .A2(new_n759), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT99), .ZN(new_n767));
  MUX2_X1   g342(.A(G32), .B(new_n767), .S(G29), .Z(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT27), .B(G1996), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G2090), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n732), .A2(G35), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n485), .B2(G29), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT29), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n768), .A2(new_n770), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n724), .A2(G21), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G168), .B2(new_n724), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(G1966), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(G1966), .ZN(new_n779));
  NOR2_X1   g354(.A1(G4), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n625), .B2(G16), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT95), .B(G1348), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n775), .A2(new_n778), .A3(new_n779), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n732), .A2(G33), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  AND2_X1   g362(.A1(new_n471), .A2(new_n472), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n788), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n787), .B1(new_n789), .B2(new_n468), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n479), .B2(G139), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT97), .Z(new_n792));
  OAI21_X1  g367(.A(new_n785), .B1(new_n792), .B2(new_n732), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT98), .B(G2072), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n793), .B(new_n794), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n724), .A2(G20), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT23), .ZN(new_n797));
  INV_X1    g372(.A(G299), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n724), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT101), .B(G1956), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n799), .B(new_n800), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n768), .A2(new_n770), .B1(new_n771), .B2(new_n774), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n757), .A2(new_n784), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n732), .A2(G25), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT90), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n481), .A2(G119), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(KEYINPUT91), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT91), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n481), .A2(new_n809), .A3(G119), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n812));
  INV_X1    g387(.A(G107), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(G2105), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n479), .B2(G131), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n806), .B1(new_n816), .B2(G29), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT92), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G1991), .Z(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT94), .ZN(new_n822));
  OR2_X1    g397(.A1(G290), .A2(KEYINPUT93), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n724), .B1(G290), .B2(KEYINPUT93), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n823), .A2(new_n824), .B1(new_n724), .B2(G24), .ZN(new_n825));
  INV_X1    g400(.A(G1986), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n820), .A2(new_n821), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT36), .ZN(new_n830));
  MUX2_X1   g405(.A(G6), .B(G305), .S(G16), .Z(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT32), .B(G1981), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n724), .A2(G22), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G166), .B2(new_n724), .ZN(new_n836));
  INV_X1    g411(.A(G1971), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n724), .A2(G23), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n590), .B2(new_n724), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT33), .B(G1976), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n833), .A2(new_n834), .A3(new_n838), .A4(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT34), .ZN(new_n844));
  OR3_X1    g419(.A1(new_n829), .A2(new_n830), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n830), .B1(new_n829), .B2(new_n844), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n804), .A2(new_n845), .A3(new_n846), .ZN(G150));
  INV_X1    g422(.A(G150), .ZN(G311));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n541), .A2(G55), .A3(new_n531), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  INV_X1    g426(.A(G93), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n851), .A2(new_n512), .B1(new_n520), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n849), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(G80), .A2(G543), .ZN(new_n855));
  INV_X1    g430(.A(G67), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n557), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n857), .A2(G651), .B1(G93), .B2(new_n535), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n541), .A2(G55), .A3(new_n531), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(KEYINPUT103), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G860), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT37), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n625), .A2(G559), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT38), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n854), .A2(new_n860), .A3(new_n562), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n850), .A2(new_n853), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(new_n562), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n858), .A2(new_n859), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n563), .A2(KEYINPUT102), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n866), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n865), .B(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n874));
  INV_X1    g449(.A(G860), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n873), .B2(KEYINPUT39), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n863), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT104), .ZN(G145));
  XNOR2_X1  g453(.A(new_n642), .B(KEYINPUT105), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(G160), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n467), .B2(new_n474), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n881), .A2(new_n882), .A3(G162), .ZN(new_n883));
  AOI21_X1  g458(.A(G162), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n792), .A2(new_n766), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(new_n792), .B2(new_n767), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n816), .A2(new_n646), .ZN(new_n888));
  INV_X1    g463(.A(new_n646), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n811), .B2(new_n815), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n479), .A2(G142), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n481), .A2(G130), .ZN(new_n893));
  OR2_X1    g468(.A1(G106), .A2(G2105), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n894), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n749), .A2(new_n500), .A3(new_n753), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n500), .B1(new_n749), .B2(new_n753), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n896), .A3(new_n898), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n891), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n891), .B1(new_n901), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n887), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n901), .A2(new_n903), .ZN(new_n908));
  INV_X1    g483(.A(new_n891), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n887), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n904), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n885), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n907), .A2(new_n912), .A3(new_n885), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n914), .A2(KEYINPUT40), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n915), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n919), .B2(new_n913), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n917), .A2(new_n920), .ZN(G395));
  INV_X1    g496(.A(KEYINPUT111), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n866), .A2(new_n869), .A3(new_n871), .ZN(new_n923));
  INV_X1    g498(.A(new_n635), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n872), .A2(new_n635), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT106), .B1(new_n624), .B2(new_n798), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n617), .A2(new_n619), .A3(new_n623), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n930), .A2(new_n931), .A3(G299), .A4(new_n612), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n617), .A2(new_n619), .A3(new_n623), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n609), .A2(G54), .A3(new_n611), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n798), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT107), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n624), .A2(new_n938), .A3(new_n798), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n928), .B1(new_n933), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n928), .B1(new_n929), .B2(new_n932), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n936), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n927), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n929), .A2(new_n932), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n925), .A2(new_n926), .B1(new_n945), .B2(new_n936), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n944), .A2(KEYINPUT110), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n590), .A2(G290), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT108), .B1(new_n600), .B2(new_n602), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n598), .A2(new_n599), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n601), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(G303), .A3(new_n953), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n951), .A2(new_n952), .A3(new_n601), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n952), .B1(new_n951), .B2(new_n601), .ZN(new_n956));
  OAI21_X1  g531(.A(G166), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n590), .A2(G290), .ZN(new_n958));
  AND4_X1   g533(.A1(new_n949), .A2(new_n954), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n954), .A2(new_n957), .B1(new_n949), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n948), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n954), .A2(new_n957), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n949), .A2(new_n958), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n954), .A2(new_n957), .A3(new_n949), .A4(new_n958), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(KEYINPUT109), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(KEYINPUT42), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT42), .B1(new_n964), .B2(new_n965), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT110), .B1(new_n944), .B2(new_n946), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n947), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n969), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n925), .A2(new_n926), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n624), .A2(new_n938), .A3(new_n798), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n938), .B1(new_n624), .B2(new_n798), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT41), .B1(new_n977), .B2(new_n945), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n945), .A2(KEYINPUT41), .A3(new_n936), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n946), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n973), .A2(new_n982), .A3(KEYINPUT110), .ZN(new_n983));
  OAI21_X1  g558(.A(G868), .B1(new_n972), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n861), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(G868), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n922), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n980), .A2(new_n989), .A3(new_n981), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n980), .B2(new_n981), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n991), .B2(new_n973), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n944), .A2(new_n946), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(new_n989), .A3(new_n969), .A4(new_n967), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n633), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n995), .A2(KEYINPUT111), .A3(new_n986), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n988), .A2(new_n996), .ZN(G295));
  NAND2_X1  g572(.A1(new_n984), .A2(new_n987), .ZN(G331));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n945), .A2(new_n936), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n544), .A2(new_n547), .A3(G301), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G301), .B1(new_n544), .B2(new_n547), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n872), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G168), .A2(G171), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n923), .B1(new_n1005), .B2(new_n1001), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1000), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n872), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n923), .A3(new_n1001), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n977), .A4(new_n942), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1000), .A2(new_n928), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n959), .A2(new_n948), .A3(new_n960), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT109), .B1(new_n964), .B2(new_n965), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G37), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1007), .A2(KEYINPUT112), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n961), .A2(new_n966), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1009), .B(new_n1008), .C1(new_n978), .C2(new_n979), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1020), .B(new_n1000), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT43), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1020), .B1(new_n1026), .B2(new_n1000), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1015), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT43), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n915), .A4(new_n1022), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n999), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n915), .A3(new_n1022), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1022), .A2(new_n1029), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1032), .A2(KEYINPUT43), .B1(new_n1033), .B2(new_n1016), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1031), .B1(new_n999), .B2(new_n1034), .ZN(G397));
  INV_X1    g610(.A(G40), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n467), .A2(new_n474), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT45), .B1(new_n500), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(G1996), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT127), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(KEYINPUT46), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(KEYINPUT46), .ZN(new_n1044));
  MUX2_X1   g619(.A(new_n1041), .B(new_n1043), .S(new_n1044), .Z(new_n1045));
  INV_X1    g620(.A(G2067), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n754), .B(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n766), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1040), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1045), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g626(.A(new_n1051), .B(KEYINPUT47), .Z(new_n1052));
  NAND2_X1  g627(.A1(new_n766), .A2(G1996), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1047), .B(new_n1053), .C1(G1996), .C2(new_n767), .ZN(new_n1054));
  XOR2_X1   g629(.A(new_n816), .B(new_n819), .Z(new_n1055));
  OAI21_X1  g630(.A(new_n1050), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1040), .A2(G290), .A3(G1986), .ZN(new_n1057));
  XOR2_X1   g632(.A(new_n1057), .B(KEYINPUT48), .Z(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n811), .A2(new_n819), .A3(new_n815), .ZN(new_n1060));
  OAI22_X1  g635(.A1(new_n1054), .A2(new_n1060), .B1(G2067), .B2(new_n754), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1050), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1052), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G303), .A2(G8), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1065), .B(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n500), .A2(new_n1038), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT45), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n1038), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(KEYINPUT114), .A3(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n500), .A2(new_n1038), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(KEYINPUT45), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1037), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n837), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1069), .A2(KEYINPUT50), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1081), .A2(new_n771), .A3(new_n1037), .A4(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT120), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G137), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1085), .B1(new_n461), .B2(new_n463), .ZN(new_n1086));
  INV_X1    g661(.A(new_n466), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n468), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n470), .A2(new_n473), .ZN(new_n1089));
  OAI211_X1 g664(.A(G40), .B(new_n1088), .C1(new_n1089), .C2(new_n468), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT120), .B(new_n1083), .C1(new_n1091), .C2(G1971), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G8), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1068), .B1(new_n1084), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n590), .B2(G1976), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT115), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1098), .B(new_n1095), .C1(new_n590), .C2(G1976), .ZN(new_n1099));
  OAI21_X1  g674(.A(G8), .B1(new_n1090), .B2(new_n1069), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(G1976), .B2(new_n590), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n598), .A2(KEYINPUT49), .ZN(new_n1103));
  INV_X1    g678(.A(G1981), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n595), .B2(KEYINPUT116), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT49), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n595), .A2(new_n1106), .A3(new_n596), .A4(new_n597), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1105), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n1100), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n588), .A2(new_n589), .ZN(new_n1111));
  INV_X1    g686(.A(new_n585), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(G1976), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G8), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1037), .B2(new_n1074), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1095), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1102), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1114), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1119), .B2(new_n1067), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1094), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1090), .A2(new_n1069), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT124), .B(KEYINPUT58), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(G1341), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G1996), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n1091), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT59), .B1(new_n1127), .B2(new_n562), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n1129));
  AOI211_X1 g704(.A(G1996), .B(new_n1090), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1129), .B(new_n563), .C1(new_n1130), .C2(new_n1125), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT56), .B(G2072), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n1038), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1135), .A2(new_n1039), .A3(new_n1075), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1069), .A2(KEYINPUT114), .A3(new_n1070), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1037), .B(new_n1134), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1081), .A2(new_n1037), .A3(new_n1082), .ZN(new_n1142));
  INV_X1    g717(.A(G1956), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1138), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1141), .B1(new_n1138), .B2(new_n1144), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1133), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n625), .A2(KEYINPUT60), .ZN(new_n1148));
  INV_X1    g723(.A(G1348), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1142), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1122), .A2(new_n1046), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n625), .A2(KEYINPUT60), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1148), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1150), .A2(KEYINPUT60), .A3(new_n625), .A4(new_n1151), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1138), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1091), .A2(new_n1134), .B1(new_n1143), .B2(new_n1142), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT123), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1159));
  OR2_X1    g734(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n1161));
  NAND2_X1  g736(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(KEYINPUT61), .B(new_n1157), .C1(new_n1158), .C2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1132), .A2(new_n1147), .A3(new_n1156), .A4(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n624), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1167), .B1(new_n1157), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT125), .B(KEYINPUT54), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n1091), .A2(new_n722), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT53), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1172), .A2(new_n1173), .B1(new_n727), .B2(new_n1142), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1071), .A2(new_n1037), .A3(new_n1072), .ZN(new_n1175));
  OR3_X1    g750(.A1(new_n1175), .A2(new_n1173), .A3(G2078), .ZN(new_n1176));
  AOI21_X1  g751(.A(G301), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1088), .A2(KEYINPUT126), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1088), .A2(KEYINPUT126), .ZN(new_n1179));
  NOR4_X1   g754(.A1(new_n474), .A2(new_n1173), .A3(new_n1036), .A4(G2078), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1077), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1142), .A2(new_n727), .ZN(new_n1182));
  AOI211_X1 g757(.A(G2078), .B(new_n1090), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1181), .B(new_n1182), .C1(new_n1183), .C2(KEYINPUT53), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1184), .A2(G171), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1171), .B1(new_n1177), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(G1966), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1175), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(G2084), .B2(new_n1142), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1190), .A2(G168), .ZN(new_n1191));
  OAI21_X1  g766(.A(G8), .B1(new_n1189), .B2(G286), .ZN(new_n1192));
  OAI21_X1  g767(.A(KEYINPUT51), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1192), .A2(KEYINPUT51), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT54), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1195), .B1(new_n1184), .B2(G171), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1174), .A2(G301), .A3(new_n1176), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1193), .A2(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1170), .A2(new_n1186), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT62), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1193), .A2(new_n1194), .A3(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1201), .A2(new_n1203), .A3(new_n1177), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1121), .B1(new_n1199), .B2(new_n1204), .ZN(new_n1205));
  NOR3_X1   g780(.A1(new_n1190), .A2(G286), .A3(new_n1114), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1083), .B1(new_n1091), .B2(G1971), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1067), .A2(G8), .A3(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1206), .A2(new_n1208), .A3(KEYINPUT63), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT122), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1067), .B1(G8), .B2(new_n1207), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1210), .B1(new_n1211), .B2(new_n1118), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1118), .ZN(new_n1213));
  OAI211_X1 g788(.A(new_n1213), .B(KEYINPUT122), .C1(new_n1119), .C2(new_n1067), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1209), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1094), .A2(new_n1120), .A3(new_n1206), .ZN(new_n1216));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n1216), .B2(KEYINPUT121), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT121), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1094), .A2(new_n1120), .A3(new_n1218), .A4(new_n1206), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1215), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n1208), .A2(new_n1118), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1110), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT118), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1223), .B1(G288), .B2(G1976), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  NOR3_X1   g800(.A1(G288), .A2(new_n1223), .A3(G1976), .ZN(new_n1226));
  OAI22_X1  g801(.A1(new_n1225), .A2(new_n1226), .B1(G1981), .B2(new_n598), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n1115), .B(KEYINPUT117), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1221), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n1229), .B(KEYINPUT119), .ZN(new_n1230));
  NOR3_X1   g805(.A1(new_n1205), .A2(new_n1220), .A3(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g806(.A(G290), .B(new_n826), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1056), .B1(new_n1040), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT113), .ZN(new_n1234));
  XNOR2_X1  g809(.A(new_n1233), .B(new_n1234), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1064), .B1(new_n1231), .B2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g811(.A(new_n684), .B(G319), .C1(new_n665), .C2(new_n666), .ZN(new_n1238));
  AOI21_X1  g812(.A(new_n1238), .B1(new_n709), .B2(new_n713), .ZN(new_n1239));
  OAI21_X1  g813(.A(new_n1239), .B1(new_n919), .B2(new_n913), .ZN(new_n1240));
  NOR2_X1   g814(.A1(new_n1240), .A2(new_n1034), .ZN(G308));
  OR2_X1    g815(.A1(new_n1240), .A2(new_n1034), .ZN(G225));
endmodule


