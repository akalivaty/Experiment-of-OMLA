//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  AND2_X1   g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n210), .A2(G20), .A3(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n205), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n208), .B(new_n212), .C1(KEYINPUT1), .C2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(KEYINPUT1), .B2(new_n219), .ZN(G361));
  XNOR2_X1  g0021(.A(G238), .B(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT2), .B(G226), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(G264), .B(G270), .Z(new_n227));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n226), .B(new_n229), .ZN(G358));
  XNOR2_X1  g0030(.A(G50), .B(G68), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G58), .B(G77), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XNOR2_X1  g0034(.A(G107), .B(G116), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G351));
  NAND3_X1  g0037(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n238));
  NAND2_X1  g0038(.A1(G1), .A2(G13), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT73), .B(G116), .ZN(new_n241));
  INV_X1    g0041(.A(G33), .ZN(new_n242));
  NOR3_X1   g0042(.A1(new_n241), .A2(G20), .A3(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT23), .ZN(new_n244));
  INV_X1    g0044(.A(G20), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n244), .B1(new_n245), .B2(G107), .ZN(new_n246));
  INV_X1    g0046(.A(G107), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(KEYINPUT23), .A3(G20), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n243), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n245), .B(G87), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT22), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT24), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n249), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n254), .B1(new_n249), .B2(new_n253), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n240), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(KEYINPUT25), .A3(new_n247), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(KEYINPUT25), .B1(new_n261), .B2(new_n247), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n259), .A2(G33), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n260), .A2(new_n265), .A3(new_n239), .A4(new_n238), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n263), .A2(new_n264), .B1(new_n247), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n258), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(G257), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  OAI211_X1 g0071(.A(G250), .B(new_n271), .C1(new_n250), .C2(new_n251), .ZN(new_n272));
  INV_X1    g0072(.A(G294), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n270), .B(new_n272), .C1(new_n242), .C2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n239), .B1(G33), .B2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n259), .A2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT5), .B(G41), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G264), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n279), .A2(new_n278), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n211), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n276), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT78), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n274), .A2(new_n275), .B1(new_n280), .B2(G264), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT78), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n290), .A3(new_n286), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(G169), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n289), .A2(G179), .A3(new_n286), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n269), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT79), .ZN(new_n296));
  AOI21_X1  g0096(.A(G190), .B1(new_n288), .B2(new_n291), .ZN(new_n297));
  AOI21_X1  g0097(.A(G200), .B1(new_n289), .B2(new_n286), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n296), .B1(new_n299), .B2(new_n269), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n249), .A2(new_n253), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT24), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n255), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n267), .B1(new_n303), .B2(new_n240), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(KEYINPUT79), .C1(new_n297), .C2(new_n298), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n295), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G41), .ZN(new_n307));
  INV_X1    g0107(.A(G45), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n259), .A2(new_n309), .B1(new_n211), .B2(new_n284), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n310), .A2(KEYINPUT68), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(KEYINPUT68), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(G238), .ZN(new_n313));
  NOR2_X1   g0113(.A1(G41), .A2(G45), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT64), .B1(new_n314), .B2(G1), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT64), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n316), .B(new_n259), .C1(G41), .C2(G45), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n285), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n223), .A2(G1698), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(G226), .B2(G1698), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n250), .A2(new_n251), .ZN(new_n322));
  INV_X1    g0122(.A(G97), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n321), .A2(new_n322), .B1(new_n242), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n275), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n313), .A2(new_n319), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT13), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n313), .A2(new_n328), .A3(new_n319), .A4(new_n325), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT14), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(G169), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT70), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n327), .B2(new_n329), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT70), .A3(new_n331), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G179), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n336), .A2(new_n331), .B1(new_n330), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G68), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n261), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT12), .ZN(new_n345));
  INV_X1    g0145(.A(new_n240), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n260), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT65), .B1(new_n245), .B2(G1), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT65), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(new_n259), .A3(G20), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n348), .A2(G68), .A3(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(G20), .A2(G33), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(G50), .B1(G20), .B2(new_n343), .ZN(new_n355));
  INV_X1    g0155(.A(G77), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n245), .A2(G33), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT11), .A3(new_n240), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n345), .A2(new_n353), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT11), .B1(new_n358), .B2(new_n240), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n342), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n327), .A2(G190), .A3(new_n329), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n362), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n327), .B2(new_n329), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT69), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n368), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT69), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n365), .A4(new_n362), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n364), .A2(new_n373), .ZN(new_n374));
  XOR2_X1   g0174(.A(KEYINPUT8), .B(G58), .Z(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n352), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n376), .A2(new_n347), .B1(new_n260), .B2(new_n375), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT7), .B1(new_n322), .B2(new_n245), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n242), .ZN(new_n381));
  NAND2_X1  g0181(.A1(KEYINPUT3), .A2(G33), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n381), .A2(KEYINPUT7), .A3(new_n245), .A4(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G58), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n343), .ZN(new_n387));
  NOR2_X1   g0187(.A1(G58), .A2(G68), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n354), .A2(G159), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT16), .B1(new_n385), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n381), .A2(new_n245), .A3(new_n382), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n343), .B1(new_n396), .B2(new_n383), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n389), .A2(KEYINPUT16), .A3(new_n390), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n240), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n378), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n318), .A2(new_n285), .B1(new_n310), .B2(G232), .ZN(new_n401));
  INV_X1    g0201(.A(G223), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n271), .ZN(new_n403));
  INV_X1    g0203(.A(G226), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G1698), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n403), .B(new_n405), .C1(new_n250), .C2(new_n251), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G87), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n275), .ZN(new_n409));
  INV_X1    g0209(.A(G190), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n401), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(G200), .B1(new_n401), .B2(new_n409), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT71), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n400), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n398), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n346), .B1(new_n385), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT16), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n397), .B2(new_n391), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n377), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n310), .A2(G232), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n319), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n211), .A2(new_n284), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n406), .B2(new_n407), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n367), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n401), .A2(new_n409), .A3(new_n410), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT71), .B1(new_n420), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT17), .B1(new_n415), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  OAI21_X1  g0230(.A(G169), .B1(new_n422), .B2(new_n424), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n401), .A2(new_n409), .A3(G179), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n400), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n430), .B1(new_n400), .B2(new_n433), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n420), .A2(new_n427), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n429), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G50), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n349), .B2(new_n351), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n348), .A2(new_n443), .B1(new_n442), .B2(new_n261), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT8), .B(G58), .ZN(new_n445));
  INV_X1    g0245(.A(G150), .ZN(new_n446));
  INV_X1    g0246(.A(new_n354), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n445), .A2(new_n357), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n245), .B1(new_n388), .B2(new_n442), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n240), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT9), .ZN(new_n452));
  INV_X1    g0252(.A(new_n319), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(G226), .B2(new_n310), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n322), .A2(new_n271), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n455), .A2(G223), .B1(G77), .B2(new_n322), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n381), .A2(new_n382), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(G222), .A3(new_n271), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n454), .B1(new_n459), .B2(new_n423), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G200), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n452), .B(new_n461), .C1(new_n410), .C2(new_n460), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT10), .ZN(new_n463));
  INV_X1    g0263(.A(new_n451), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n460), .B2(new_n335), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(G179), .B2(new_n460), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n447), .A2(KEYINPUT66), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n447), .A2(KEYINPUT66), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n469), .A2(new_n445), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT15), .B(G87), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n472), .A2(new_n357), .B1(new_n245), .B2(new_n356), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n346), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n352), .A2(G77), .ZN(new_n476));
  OAI22_X1  g0276(.A1(new_n476), .A2(new_n347), .B1(G77), .B2(new_n260), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n455), .A2(G238), .B1(G107), .B2(new_n322), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n457), .A2(G232), .A3(new_n271), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n275), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n453), .B1(G244), .B2(new_n310), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n478), .B1(new_n485), .B2(new_n367), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n486), .A2(KEYINPUT67), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(G190), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(KEYINPUT67), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n478), .B1(new_n484), .B2(new_n335), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(G179), .B2(new_n484), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NOR4_X1   g0293(.A1(new_n374), .A2(new_n441), .A3(new_n467), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n457), .A2(new_n245), .A3(G68), .ZN(new_n495));
  NAND3_X1  g0295(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n245), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n203), .B2(G87), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n357), .A2(new_n323), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n495), .B(new_n498), .C1(KEYINPUT19), .C2(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(new_n240), .B1(new_n261), .B2(new_n472), .ZN(new_n501));
  INV_X1    g0301(.A(new_n266), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G87), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(G238), .B(new_n271), .C1(new_n250), .C2(new_n251), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n505), .B(new_n506), .C1(new_n242), .C2(new_n241), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n275), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n285), .A2(new_n278), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n423), .A2(G250), .A3(new_n277), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G200), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n275), .B2(new_n507), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT74), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n515), .A3(G190), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n514), .B2(G190), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n504), .B(new_n512), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n472), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n502), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n501), .A2(new_n521), .B1(new_n514), .B2(new_n339), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n511), .A2(new_n335), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n519), .A2(KEYINPUT75), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT75), .B1(new_n519), .B2(new_n524), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n280), .A2(G257), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n286), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n457), .A2(G250), .A3(G1698), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G283), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(G244), .B(new_n271), .C1(new_n250), .C2(new_n251), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(KEYINPUT72), .A3(new_n535), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT72), .B1(new_n534), .B2(new_n535), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n533), .B(new_n536), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n530), .B1(new_n540), .B2(new_n275), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n339), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n247), .A2(KEYINPUT6), .A3(G97), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n323), .A2(new_n247), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(new_n202), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n543), .B1(new_n545), .B2(KEYINPUT6), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(G20), .B1(G77), .B2(new_n354), .ZN(new_n547));
  OAI21_X1  g0347(.A(G107), .B1(new_n379), .B2(new_n384), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n346), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n502), .A2(G97), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(G97), .B2(new_n260), .ZN(new_n551));
  OR2_X1    g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n542), .B(new_n552), .C1(G169), .C2(new_n541), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n532), .B(new_n245), .C1(G33), .C2(new_n323), .ZN(new_n554));
  INV_X1    g0354(.A(G116), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT73), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT73), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G116), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n240), .B(new_n554), .C1(new_n559), .C2(new_n245), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT20), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n241), .A2(G20), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(KEYINPUT20), .A3(new_n240), .A4(new_n554), .ZN(new_n564));
  INV_X1    g0364(.A(G13), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(G1), .ZN(new_n566));
  INV_X1    g0366(.A(new_n563), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n562), .A2(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OR3_X1    g0368(.A1(new_n266), .A2(KEYINPUT76), .A3(new_n555), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT76), .B1(new_n266), .B2(new_n555), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n280), .A2(G270), .B1(new_n282), .B2(new_n285), .ZN(new_n573));
  OAI211_X1 g0373(.A(G264), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n574));
  OAI211_X1 g0374(.A(G257), .B(new_n271), .C1(new_n250), .C2(new_n251), .ZN(new_n575));
  INV_X1    g0375(.A(G303), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n457), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n275), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n335), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n572), .A2(new_n579), .A3(KEYINPUT21), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n573), .A2(G179), .A3(new_n578), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n572), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT21), .B1(new_n572), .B2(new_n579), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n572), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n367), .B1(new_n573), .B2(new_n578), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT77), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n573), .A2(G190), .A3(new_n578), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n586), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n571), .A3(new_n568), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT77), .B1(new_n592), .B2(new_n587), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n540), .A2(new_n275), .ZN(new_n595));
  INV_X1    g0395(.A(new_n530), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(G190), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n549), .A2(new_n551), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(new_n598), .C1(new_n367), .C2(new_n541), .ZN(new_n599));
  AND4_X1   g0399(.A1(new_n553), .A2(new_n585), .A3(new_n594), .A4(new_n599), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n306), .A2(new_n494), .A3(new_n528), .A4(new_n600), .ZN(G372));
  OAI21_X1  g0401(.A(new_n414), .B1(new_n400), .B2(new_n413), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n420), .A2(KEYINPUT71), .A3(new_n427), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n439), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n440), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n369), .A2(new_n372), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n606), .A2(new_n492), .ZN(new_n607));
  AOI211_X1 g0407(.A(new_n604), .B(new_n605), .C1(new_n607), .C2(new_n364), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n400), .A2(new_n433), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT18), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n434), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n463), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n612), .A2(new_n466), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n513), .A2(KEYINPUT80), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT80), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n509), .B2(new_n510), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n508), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n522), .B1(new_n618), .B2(G169), .ZN(new_n619));
  XOR2_X1   g0419(.A(new_n619), .B(KEYINPUT82), .Z(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(G200), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n504), .B(new_n621), .C1(new_n517), .C2(new_n518), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n553), .A2(new_n599), .A3(new_n619), .A4(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n300), .B2(new_n305), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n269), .A2(new_n294), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(KEYINPUT81), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT81), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n269), .B2(new_n294), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n585), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n620), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n519), .A2(new_n524), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT75), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n553), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n525), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g0435(.A(KEYINPUT83), .B(KEYINPUT26), .Z(new_n636));
  NAND2_X1  g0436(.A1(new_n622), .A2(new_n619), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(new_n553), .ZN(new_n638));
  OAI22_X1  g0438(.A1(new_n635), .A2(new_n636), .B1(new_n638), .B2(KEYINPUT26), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n630), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n494), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n613), .A2(new_n641), .ZN(G369));
  NAND2_X1  g0442(.A1(new_n566), .A2(new_n245), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n572), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n585), .A2(new_n594), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n585), .B2(new_n649), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G330), .ZN(new_n652));
  XOR2_X1   g0452(.A(new_n652), .B(KEYINPUT84), .Z(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n648), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n306), .B1(new_n304), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n625), .B2(new_n655), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT85), .Z(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n585), .A2(new_n648), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n306), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n626), .A2(new_n628), .A3(new_n648), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n660), .A2(new_n665), .ZN(G399));
  NOR3_X1   g0466(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n206), .A2(new_n307), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(G1), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n209), .B2(new_n668), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n635), .A2(new_n636), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n638), .A2(KEYINPUT26), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n620), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n623), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n300), .A2(new_n305), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n625), .A2(new_n585), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT89), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n624), .A2(KEYINPUT89), .A3(new_n677), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n674), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT90), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT29), .A4(new_n655), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n682), .A2(KEYINPUT29), .A3(new_n655), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n648), .B1(new_n630), .B2(new_n639), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT90), .B1(new_n686), .B2(KEYINPUT29), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n306), .A2(new_n600), .A3(new_n528), .A4(new_n655), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT31), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n655), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT86), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n514), .A2(new_n289), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n514), .B2(new_n289), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n541), .B(new_n581), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT30), .ZN(new_n698));
  AOI21_X1  g0498(.A(G179), .B1(new_n573), .B2(new_n578), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n699), .A2(new_n617), .A3(new_n287), .ZN(new_n700));
  INV_X1    g0500(.A(new_n541), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n697), .A2(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT87), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n514), .A2(new_n289), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT86), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n694), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(KEYINPUT30), .A3(new_n541), .A4(new_n581), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n702), .B2(new_n703), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n692), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n697), .A2(new_n698), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n700), .A2(new_n701), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT88), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT88), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n702), .A2(new_n715), .A3(new_n708), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n655), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n690), .B(new_n710), .C1(new_n717), .C2(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n689), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n671), .B1(new_n721), .B2(G1), .ZN(G364));
  NOR2_X1   g0522(.A1(new_n565), .A2(G20), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n259), .B1(new_n723), .B2(G45), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n668), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n653), .B(new_n728), .C1(G330), .C2(new_n651), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT91), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n206), .B(new_n457), .C1(G355), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT91), .B1(new_n203), .B2(G87), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n731), .A2(new_n732), .B1(G116), .B2(new_n206), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n233), .A2(new_n308), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n322), .A2(new_n206), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n308), .B2(new_n210), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n733), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n239), .B1(G20), .B2(new_n335), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n727), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n245), .A2(new_n410), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n367), .A2(G179), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n322), .B1(new_n747), .B2(new_n576), .ZN(new_n748));
  NAND3_X1  g0548(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n410), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n748), .B1(G326), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(G179), .A3(new_n367), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n245), .A2(G190), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n746), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n753), .A2(G322), .B1(new_n756), .B2(G283), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n754), .A2(G179), .A3(new_n367), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G179), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n754), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n759), .A2(G311), .B1(new_n762), .B2(G329), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n245), .B1(new_n760), .B2(G190), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n749), .A2(G190), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT33), .B(G317), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n765), .A2(G294), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n751), .A2(new_n757), .A3(new_n763), .A4(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n750), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n442), .A2(new_n770), .B1(new_n752), .B2(new_n386), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n759), .A2(KEYINPUT92), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n759), .A2(KEYINPUT92), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n771), .B1(new_n776), .B2(G77), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT93), .Z(new_n778));
  XNOR2_X1  g0578(.A(new_n764), .B(KEYINPUT94), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G97), .ZN(new_n780));
  INV_X1    g0580(.A(G87), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n457), .B1(new_n747), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(G107), .B2(new_n756), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n761), .A2(KEYINPUT32), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(G68), .B2(new_n766), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT32), .B1(new_n761), .B2(new_n784), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n780), .A2(new_n783), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n769), .B1(new_n778), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n744), .B1(new_n789), .B2(new_n741), .ZN(new_n790));
  INV_X1    g0590(.A(new_n740), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n651), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n729), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G396));
  NOR2_X1   g0594(.A1(new_n492), .A2(new_n648), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n648), .B1(new_n475), .B2(new_n477), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n490), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n795), .B1(new_n797), .B2(new_n492), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n686), .B(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n727), .B1(new_n799), .B2(new_n719), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n719), .B2(new_n799), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n753), .A2(G143), .B1(G137), .B2(new_n750), .ZN(new_n802));
  INV_X1    g0602(.A(new_n766), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n802), .B1(new_n446), .B2(new_n803), .C1(new_n775), .C2(new_n784), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT34), .Z(new_n805));
  NOR2_X1   g0605(.A1(new_n764), .A2(new_n386), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n457), .B1(new_n747), .B2(new_n442), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n756), .A2(G68), .ZN(new_n808));
  INV_X1    g0608(.A(G132), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n809), .B2(new_n761), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n805), .A2(new_n806), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n776), .A2(new_n559), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n322), .B1(new_n747), .B2(new_n247), .C1(new_n576), .C2(new_n770), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G283), .B2(new_n766), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n752), .A2(new_n273), .B1(new_n761), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G87), .B2(new_n756), .ZN(new_n817));
  AND4_X1   g0617(.A1(new_n780), .A2(new_n812), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n741), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n741), .A2(new_n738), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT95), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n728), .B1(new_n822), .B2(new_n356), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n819), .B(new_n823), .C1(new_n798), .C2(new_n739), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n801), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G384));
  NAND2_X1  g0626(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n239), .A2(new_n245), .A3(new_n555), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n546), .B2(KEYINPUT35), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT96), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT36), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n210), .B(G77), .C1(new_n386), .C2(new_n343), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n442), .A2(G68), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n259), .B(G13), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n795), .B1(new_n686), .B2(new_n798), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  INV_X1    g0640(.A(new_n646), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT97), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n417), .A2(new_n419), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(new_n378), .ZN(new_n844));
  AOI211_X1 g0644(.A(KEYINPUT97), .B(new_n377), .C1(new_n417), .C2(new_n419), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n840), .B1(new_n441), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n433), .B1(new_n844), .B2(new_n845), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n846), .A2(new_n849), .A3(new_n602), .A4(new_n603), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT37), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT37), .B1(new_n400), .B2(new_n433), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n400), .A2(new_n841), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n602), .A2(new_n852), .A3(new_n603), .A4(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT98), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT98), .ZN(new_n856));
  AND4_X1   g0656(.A1(new_n602), .A2(new_n852), .A3(new_n603), .A4(new_n853), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(new_n850), .C2(KEYINPUT37), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n848), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n604), .A2(new_n611), .A3(new_n605), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(new_n846), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n602), .A2(new_n603), .ZN(new_n863));
  INV_X1    g0663(.A(new_n433), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n400), .A2(KEYINPUT97), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n843), .A2(new_n842), .A3(new_n378), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n862), .B1(new_n868), .B2(new_n846), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n856), .B1(new_n869), .B2(new_n857), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n851), .A2(KEYINPUT98), .A3(new_n854), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n861), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n859), .B1(new_n872), .B2(KEYINPUT38), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n363), .B(new_n648), .C1(new_n606), .C2(new_n342), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n362), .A2(new_n655), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n340), .B1(new_n334), .B2(new_n337), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n373), .B(new_n876), .C1(new_n877), .C2(new_n362), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n839), .A2(new_n873), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n437), .B2(new_n841), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT38), .B1(new_n860), .B2(new_n846), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n870), .B2(new_n871), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  INV_X1    g0684(.A(new_n853), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n609), .A2(new_n853), .A3(new_n438), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n441), .A2(new_n885), .B1(new_n887), .B2(new_n854), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n884), .B1(new_n888), .B2(KEYINPUT38), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n883), .A2(KEYINPUT99), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT99), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n854), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n860), .B2(new_n853), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT39), .B1(new_n893), .B2(new_n840), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n891), .B1(new_n859), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n855), .A2(new_n858), .B1(new_n860), .B2(new_n846), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n840), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n884), .B1(new_n898), .B2(new_n859), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT100), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT99), .B1(new_n883), .B2(new_n889), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n859), .A2(new_n891), .A3(new_n894), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT100), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n364), .A2(new_n648), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n881), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n688), .A2(new_n494), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n613), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n909), .B(new_n911), .Z(new_n912));
  NAND2_X1  g0712(.A1(new_n879), .A2(new_n798), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n713), .A2(KEYINPUT88), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n715), .B1(new_n702), .B2(new_n708), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n692), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n690), .B(new_n916), .C1(new_n717), .C2(KEYINPUT31), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT101), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n648), .B1(new_n914), .B2(new_n915), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n691), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT101), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n920), .A2(new_n921), .A3(new_n690), .A4(new_n916), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n913), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n873), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n893), .A2(new_n840), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n859), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n925), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n923), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n918), .A2(new_n922), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n494), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n931), .A2(new_n933), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(G330), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n912), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n259), .B2(new_n723), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n912), .A2(new_n936), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n837), .B1(new_n938), .B2(new_n939), .ZN(G367));
  OAI211_X1 g0740(.A(new_n553), .B(new_n599), .C1(new_n598), .C2(new_n655), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n553), .B2(new_n655), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT102), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT44), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n942), .B(new_n665), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n665), .A2(new_n942), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT45), .Z(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(new_n659), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n659), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n662), .B1(new_n657), .B2(new_n661), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n653), .B(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n720), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n668), .B(KEYINPUT41), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n724), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n659), .A2(new_n942), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n663), .A2(new_n942), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n553), .B1(new_n941), .B2(new_n625), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n961), .A2(KEYINPUT42), .B1(new_n655), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(KEYINPUT42), .B2(new_n961), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT43), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n504), .A2(new_n655), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n637), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n620), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n964), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n965), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n960), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n959), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(G283), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n775), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n747), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(KEYINPUT46), .A3(G116), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n977), .B1(new_n323), .B2(new_n755), .C1(new_n978), .C2(new_n761), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT46), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n747), .B2(new_n241), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n247), .B2(new_n764), .C1(new_n803), .C2(new_n273), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n322), .B1(new_n752), .B2(new_n576), .C1(new_n815), .C2(new_n770), .ZN(new_n983));
  NOR4_X1   g0783(.A1(new_n975), .A2(new_n979), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT104), .Z(new_n985));
  AOI22_X1  g0785(.A1(G58), .A2(new_n976), .B1(new_n762), .B2(G137), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n446), .B2(new_n752), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n322), .B1(new_n756), .B2(G77), .ZN(new_n988));
  INV_X1    g0788(.A(G143), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n988), .B1(new_n770), .B2(new_n989), .C1(new_n784), .C2(new_n803), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n987), .B(new_n990), .C1(G50), .C2(new_n776), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n779), .A2(G68), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n985), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT47), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n741), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n968), .A2(new_n740), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n742), .B1(new_n206), .B2(new_n472), .C1(new_n229), .C2(new_n735), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n998), .A2(KEYINPUT103), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(KEYINPUT103), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n999), .A2(new_n1000), .A3(new_n728), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n996), .A2(new_n997), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n973), .A2(new_n1002), .ZN(G387));
  NAND2_X1  g0803(.A1(new_n721), .A2(new_n956), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n720), .A2(new_n955), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n726), .A3(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n752), .A2(new_n442), .B1(new_n758), .B2(new_n343), .ZN(new_n1007));
  XOR2_X1   g0807(.A(KEYINPUT106), .B(G150), .Z(new_n1008));
  OAI22_X1  g0808(.A1(new_n1008), .A2(new_n761), .B1(new_n747), .B2(new_n356), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n779), .A2(new_n520), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n457), .B1(new_n755), .B2(new_n323), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n375), .B2(new_n766), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n750), .A2(G159), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n750), .A2(G322), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n753), .A2(G317), .B1(G311), .B2(new_n766), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n775), .C2(new_n576), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT48), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n976), .A2(G294), .B1(new_n765), .B2(G283), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT49), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(KEYINPUT107), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n457), .B1(new_n762), .B2(G326), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n241), .C2(new_n755), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1024), .A2(KEYINPUT107), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1015), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n741), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n667), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(new_n206), .A3(new_n457), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(G107), .B2(new_n206), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n226), .A2(new_n308), .ZN(new_n1034));
  AOI211_X1 g0834(.A(G45), .B(new_n1031), .C1(G68), .C2(G77), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n445), .A2(G50), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n735), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1033), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n727), .B1(new_n1039), .B2(new_n743), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT105), .Z(new_n1041));
  OAI211_X1 g0841(.A(new_n1030), .B(new_n1041), .C1(new_n657), .C2(new_n791), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1006), .B(new_n1042), .C1(new_n724), .C2(new_n955), .ZN(G393));
  NAND3_X1  g0843(.A1(new_n953), .A2(new_n721), .A3(new_n956), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT108), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n951), .A2(new_n1045), .A3(new_n952), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n950), .A2(new_n659), .A3(KEYINPUT108), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n1004), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1044), .A2(new_n726), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n725), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n742), .B1(new_n323), .B2(new_n206), .C1(new_n236), .C2(new_n735), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n727), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n978), .A2(new_n770), .B1(new_n752), .B2(new_n815), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT52), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n322), .B1(new_n755), .B2(new_n247), .C1(new_n803), .C2(new_n576), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n559), .B2(new_n765), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n758), .A2(new_n273), .B1(new_n747), .B2(new_n974), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G322), .B2(new_n762), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n457), .B1(new_n755), .B2(new_n781), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n747), .A2(new_n343), .B1(new_n761), .B2(new_n989), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(G50), .C2(new_n766), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n779), .A2(G77), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n445), .C2(new_n775), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n753), .A2(G159), .B1(G150), .B2(new_n750), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1060), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1053), .B1(new_n1068), .B2(new_n741), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n942), .B2(new_n791), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1049), .A2(new_n1051), .A3(new_n1070), .ZN(G390));
  INV_X1    g0871(.A(new_n908), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n879), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1072), .B1(new_n838), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n900), .A2(new_n906), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n928), .A2(new_n908), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n797), .A2(new_n492), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n682), .A2(new_n655), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n795), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1076), .B1(new_n1081), .B2(new_n1073), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n718), .A2(new_n879), .A3(G330), .A4(new_n798), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1075), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n908), .B(new_n928), .C1(new_n1080), .C2(new_n879), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n905), .B1(new_n901), .B2(new_n904), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1088), .B2(new_n1074), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n879), .A2(new_n798), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n932), .A2(G330), .A3(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(KEYINPUT109), .B(new_n1084), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1091), .B1(new_n1075), .B2(new_n1082), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT109), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1088), .A2(new_n738), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n821), .A2(new_n375), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n808), .B1(new_n555), .B2(new_n752), .C1(new_n273), .C2(new_n761), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n457), .B1(new_n976), .B2(G87), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n770), .B2(new_n974), .C1(new_n247), .C2(new_n803), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1099), .B(new_n1101), .C1(G97), .C2(new_n776), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n779), .A2(G159), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT54), .B(G143), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n775), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1008), .A2(new_n747), .ZN(new_n1106));
  XOR2_X1   g0906(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n1107));
  XNOR2_X1  g0907(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n766), .A2(G137), .B1(new_n750), .B2(G128), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n322), .B1(new_n762), .B2(G125), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n442), .B2(new_n755), .C1(new_n809), .C2(new_n752), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1105), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1102), .A2(new_n1064), .B1(new_n1103), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n728), .B(new_n1098), .C1(new_n1115), .C2(new_n741), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1096), .A2(new_n725), .B1(new_n1097), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT111), .ZN(new_n1118));
  AOI211_X1 g0918(.A(KEYINPUT109), .B(new_n1091), .C1(new_n1075), .C2(new_n1082), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1075), .A2(new_n1082), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1091), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1094), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1119), .B1(new_n1122), .B2(new_n1084), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n718), .A2(G330), .A3(new_n798), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n1073), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT110), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1124), .A2(KEYINPUT110), .A3(new_n1073), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1091), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n839), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n932), .A2(G330), .A3(new_n798), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n1073), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1078), .A2(new_n1083), .A3(new_n1079), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1130), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n932), .A2(G330), .A3(new_n494), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n910), .A2(new_n613), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1118), .B(new_n726), .C1(new_n1123), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(KEYINPUT112), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1129), .A2(new_n839), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n910), .A2(new_n613), .A3(new_n1136), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT112), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1123), .A2(new_n1140), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1139), .A2(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1075), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1148), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1143), .B1(new_n1149), .B2(new_n1119), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1118), .B1(new_n1150), .B2(new_n726), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1117), .B1(new_n1147), .B2(new_n1151), .ZN(G378));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1142), .B1(new_n1096), .B2(new_n1143), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT115), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n464), .A2(new_n646), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n467), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1158), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n463), .B2(new_n466), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1157), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1159), .A2(new_n1161), .A3(new_n1157), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1155), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(KEYINPUT115), .A3(new_n1162), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n926), .A2(G330), .A3(new_n930), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n930), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT40), .B1(new_n923), .B2(new_n873), .ZN(new_n1171));
  INV_X1    g0971(.A(G330), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1169), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n909), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n926), .A2(G330), .A3(new_n930), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1174), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1088), .A2(new_n1072), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1169), .C1(new_n1180), .C2(new_n881), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1153), .B1(new_n1154), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1137), .B1(new_n1123), .B2(new_n1138), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1182), .A2(new_n1153), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n668), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1182), .A2(new_n724), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n820), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n727), .B1(G50), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1168), .A2(new_n739), .ZN(new_n1191));
  INV_X1    g0991(.A(G128), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n752), .A2(new_n1192), .B1(new_n747), .B2(new_n1104), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G137), .B2(new_n759), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n766), .A2(G132), .B1(new_n750), .B2(G125), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n779), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1194), .B(new_n1195), .C1(new_n446), .C2(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n242), .B(new_n307), .C1(new_n755), .C2(new_n784), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G124), .B2(new_n762), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n457), .A2(G41), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n356), .B2(new_n747), .C1(new_n803), .C2(new_n323), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G116), .B2(new_n750), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n520), .A2(new_n759), .B1(new_n756), .B2(G58), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n753), .A2(G107), .B1(new_n762), .B2(G283), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1205), .A2(new_n992), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT58), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G50), .B(new_n1203), .C1(new_n242), .C2(new_n307), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT114), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1202), .A2(new_n1210), .A3(new_n1211), .A4(new_n1213), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1190), .B(new_n1191), .C1(new_n741), .C2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1188), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1187), .A2(new_n1216), .ZN(G375));
  NAND2_X1  g1017(.A1(new_n1073), .A2(new_n738), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n727), .B1(new_n821), .B2(G68), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n753), .A2(G137), .B1(new_n762), .B2(G128), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n446), .B2(new_n758), .C1(new_n784), .C2(new_n747), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n809), .A2(new_n770), .B1(new_n803), .B2(new_n1104), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n457), .B1(new_n755), .B2(new_n386), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT116), .Z(new_n1225));
  OAI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(new_n442), .C2(new_n1196), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n776), .A2(G107), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n322), .B1(new_n755), .B2(new_n356), .C1(new_n803), .C2(new_n241), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G294), .B2(new_n750), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n752), .A2(new_n974), .B1(new_n761), .B2(new_n576), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G97), .B2(new_n976), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1227), .A2(new_n1011), .A3(new_n1229), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1226), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1219), .B1(new_n1233), .B2(new_n741), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1135), .A2(new_n725), .B1(new_n1218), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n958), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1235), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT117), .Z(G381));
  NOR4_X1   g1041(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1242));
  INV_X1    g1042(.A(G387), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NOR4_X1   g1044(.A1(new_n1244), .A2(G375), .A3(G378), .A4(G381), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT118), .ZN(G407));
  NAND2_X1  g1046(.A1(new_n647), .A2(G213), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(G375), .A2(G378), .A3(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT119), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(G213), .A3(new_n1249), .ZN(G409));
  AND3_X1   g1050(.A1(new_n1177), .A2(new_n1181), .A3(new_n1238), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1138), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1142), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT120), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT121), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n724), .B1(new_n1182), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1177), .A2(new_n1181), .A3(KEYINPUT121), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1215), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1184), .A2(KEYINPUT120), .A3(new_n1251), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1255), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT111), .B1(new_n1252), .B2(new_n668), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n1146), .A3(new_n1139), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1263), .A3(new_n1117), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G378), .A2(new_n1187), .A3(new_n1216), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT122), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT122), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1271), .B(new_n1237), .C1(new_n1143), .C2(new_n1267), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n668), .B1(new_n1269), .B2(KEYINPUT60), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1274), .A2(G384), .A3(new_n1235), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G384), .B1(new_n1274), .B2(new_n1235), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1266), .A2(new_n1247), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(KEYINPUT124), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1266), .A2(new_n1247), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1247), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(G2897), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(KEYINPUT123), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1277), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1284), .B1(new_n1277), .B2(new_n1285), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1282), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1266), .A2(new_n1247), .A3(new_n1277), .A4(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1281), .A2(new_n1289), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1288), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1296), .A2(new_n1281), .A3(KEYINPUT125), .A4(new_n1292), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(G393), .B(new_n793), .ZN(new_n1298));
  OR2_X1    g1098(.A1(G390), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G390), .A2(new_n1298), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1243), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1243), .A2(new_n1300), .A3(new_n1299), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(KEYINPUT126), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT126), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1303), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(new_n1301), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1295), .A2(new_n1297), .A3(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1278), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1311), .A2(KEYINPUT63), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1306), .A2(new_n1301), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(KEYINPUT63), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .A4(new_n1296), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1310), .A2(new_n1315), .ZN(G405));
  XNOR2_X1  g1116(.A(G375), .B(G378), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1277), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1318), .A2(KEYINPUT127), .ZN(new_n1319));
  AND2_X1   g1119(.A1(new_n1318), .A2(KEYINPUT127), .ZN(new_n1320));
  OR3_X1    g1120(.A1(new_n1317), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1319), .B1(new_n1317), .B2(new_n1320), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1323), .B(new_n1308), .ZN(G402));
endmodule


