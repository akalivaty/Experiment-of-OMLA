//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  INV_X1    g006(.A(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(KEYINPUT26), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT27), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(G190gat), .B1(new_n216), .B2(KEYINPUT67), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT28), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT28), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n219), .A2(new_n224), .A3(G190gat), .ZN(new_n225));
  OAI221_X1 g024(.A(new_n206), .B1(new_n210), .B2(new_n214), .C1(new_n223), .C2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n212), .A2(KEYINPUT23), .B1(new_n211), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n206), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n209), .B2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n230), .A2(KEYINPUT66), .A3(new_n235), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n234), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n232), .A2(KEYINPUT64), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n206), .A2(new_n242), .A3(new_n231), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n240), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n209), .A2(new_n237), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n211), .A3(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n236), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n235), .A2(new_n238), .A3(new_n229), .A4(new_n228), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n239), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G226gat), .ZN(new_n253));
  INV_X1    g052(.A(G233gat), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n226), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT22), .ZN(new_n258));
  INV_X1    g057(.A(G211gat), .ZN(new_n259));
  INV_X1    g058(.A(G218gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n257), .A3(new_n261), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(KEYINPUT70), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n262), .A2(new_n268), .A3(new_n264), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n253), .A2(new_n254), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(KEYINPUT29), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n272), .B1(new_n226), .B2(new_n252), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n256), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n270), .ZN(new_n275));
  INV_X1    g074(.A(new_n273), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(new_n255), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n205), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n270), .B1(new_n256), .B2(new_n273), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n275), .A3(new_n255), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(new_n280), .A3(new_n204), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(KEYINPUT30), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n279), .A2(new_n280), .A3(new_n283), .A4(new_n204), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n286));
  OR2_X1    g085(.A1(KEYINPUT71), .A2(G148gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(KEYINPUT71), .A2(G148gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(G141gat), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G141gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G148gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n293), .B1(new_n296), .B2(KEYINPUT2), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G148gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G141gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n291), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n296), .A2(new_n293), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G127gat), .B(G134gat), .Z(new_n307));
  XNOR2_X1  g106(.A(G113gat), .B(G120gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(KEYINPUT1), .B2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(G113gat), .B(G120gat), .Z(new_n310));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311));
  XNOR2_X1  g110(.A(G127gat), .B(G134gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n286), .B1(new_n306), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n309), .A2(new_n313), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n292), .A2(new_n297), .B1(new_n303), .B2(new_n304), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT4), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n316), .B1(KEYINPUT3), .B2(new_n306), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT72), .B(KEYINPUT3), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  AND4_X1   g123(.A1(new_n322), .A2(new_n298), .A3(new_n305), .A4(new_n323), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n320), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT5), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n306), .B(new_n314), .ZN(new_n330));
  INV_X1    g129(.A(new_n327), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G1gat), .B(G29gat), .Z(new_n334));
  XNOR2_X1  g133(.A(G57gat), .B(G85gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n320), .A2(new_n326), .A3(new_n329), .A4(new_n327), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n333), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n333), .B2(new_n339), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT6), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n341), .A2(KEYINPUT6), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n285), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n265), .A2(KEYINPUT75), .A3(new_n266), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n266), .A2(KEYINPUT75), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n323), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n306), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n298), .A2(new_n305), .A3(new_n323), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT73), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n317), .A2(new_n322), .A3(new_n323), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT29), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n350), .B1(new_n354), .B2(new_n275), .ZN(new_n355));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n347), .B1(new_n324), .B2(new_n325), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n270), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n267), .A2(new_n347), .A3(new_n269), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n356), .B1(new_n361), .B2(new_n306), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n355), .A2(new_n356), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G22gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n306), .ZN(new_n367));
  INV_X1    g166(.A(new_n356), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n367), .B(new_n368), .C1(new_n354), .C2(new_n275), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n357), .A2(new_n270), .B1(new_n306), .B2(new_n349), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n369), .B(new_n364), .C1(new_n370), .C2(new_n368), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G78gat), .B(G106gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT31), .B(G50gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n374), .B(new_n375), .Z(new_n376));
  AOI21_X1  g175(.A(new_n366), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n376), .ZN(new_n378));
  AOI211_X1 g177(.A(KEYINPUT77), .B(new_n378), .C1(new_n371), .C2(new_n372), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n365), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT76), .B1(new_n363), .B2(new_n364), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT77), .B1(new_n381), .B2(new_n378), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n363), .B(G22gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n373), .A2(new_n366), .A3(new_n376), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n344), .A2(new_n380), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G227gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(new_n254), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n226), .A2(new_n252), .A3(new_n316), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n316), .B1(new_n226), .B2(new_n252), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT68), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT68), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n393), .B(new_n388), .C1(new_n389), .C2(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT32), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n226), .A2(new_n252), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n314), .ZN(new_n398));
  INV_X1    g197(.A(new_n388), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n226), .A2(new_n252), .A3(new_n316), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT34), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT33), .B1(new_n392), .B2(new_n394), .ZN(new_n404));
  XNOR2_X1  g203(.A(G15gat), .B(G43gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT69), .ZN(new_n406));
  INV_X1    g205(.A(G71gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(G99gat), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n403), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n401), .B(KEYINPUT34), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n409), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n396), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(new_n411), .A3(new_n414), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n403), .B1(new_n404), .B2(new_n409), .ZN(new_n418));
  INV_X1    g217(.A(new_n396), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(KEYINPUT36), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT36), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n419), .B1(new_n417), .B2(new_n418), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n285), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT39), .B1(new_n330), .B2(new_n331), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n320), .A2(new_n326), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n331), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n314), .B1(new_n317), .B2(new_n360), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(new_n352), .B2(new_n353), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n331), .B1(new_n432), .B2(new_n319), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n433), .A2(KEYINPUT39), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n430), .A2(KEYINPUT40), .A3(new_n434), .A4(new_n338), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT40), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n338), .B1(new_n433), .B2(KEYINPUT39), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(new_n429), .ZN(new_n438));
  INV_X1    g237(.A(new_n341), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n380), .A2(new_n385), .B1(new_n426), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT80), .B1(new_n342), .B2(new_n343), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n343), .A2(KEYINPUT80), .ZN(new_n443));
  INV_X1    g242(.A(new_n281), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n279), .A2(new_n280), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT37), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n204), .B1(new_n279), .B2(new_n280), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT37), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n204), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(KEYINPUT79), .B(KEYINPUT38), .Z(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n444), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n448), .B1(new_n274), .B2(KEYINPUT78), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(KEYINPUT78), .B2(new_n445), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n455), .B(new_n451), .C1(new_n447), .C2(new_n449), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n442), .A2(new_n443), .A3(new_n453), .A4(new_n456), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n421), .A2(new_n425), .B1(new_n441), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n380), .A2(new_n385), .ZN(new_n459));
  OR3_X1    g258(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT6), .ZN(new_n460));
  INV_X1    g259(.A(new_n343), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n460), .A2(new_n461), .B1(new_n284), .B2(new_n282), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n459), .A2(new_n462), .A3(new_n420), .A4(new_n416), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n423), .A2(new_n424), .ZN(new_n465));
  XOR2_X1   g264(.A(KEYINPUT81), .B(KEYINPUT35), .Z(new_n466));
  NAND2_X1  g265(.A1(new_n285), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n467), .B1(new_n442), .B2(new_n443), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n468), .A3(new_n459), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n386), .A2(new_n458), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G15gat), .B(G22gat), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n471), .A2(G1gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT16), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n473), .B2(G1gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(KEYINPUT86), .A2(G8gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n477));
  INV_X1    g276(.A(G8gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n472), .A2(new_n474), .A3(new_n480), .A4(new_n475), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(G43gat), .A2(G50gat), .ZN(new_n483));
  NOR2_X1   g282(.A1(G43gat), .A2(G50gat), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT15), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G29gat), .A2(G36gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT82), .ZN(new_n489));
  NOR4_X1   g288(.A1(new_n489), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n491));
  INV_X1    g290(.A(G36gat), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT82), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n488), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n487), .B1(new_n494), .B2(KEYINPUT83), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT83), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(new_n488), .C1(new_n490), .C2(new_n493), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n485), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT14), .ZN(new_n499));
  INV_X1    g298(.A(G29gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n492), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n488), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(new_n485), .A3(new_n486), .ZN(new_n503));
  INV_X1    g302(.A(G43gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT84), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G43gat), .ZN(new_n507));
  INV_X1    g306(.A(G50gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n483), .A2(KEYINPUT15), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT85), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT85), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n513), .A3(new_n510), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n503), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n498), .A2(KEYINPUT17), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n517));
  INV_X1    g316(.A(new_n485), .ZN(new_n518));
  INV_X1    g317(.A(new_n488), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n489), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n491), .A2(KEYINPUT82), .A3(new_n492), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n486), .B1(new_n522), .B2(new_n496), .ZN(new_n523));
  INV_X1    g322(.A(new_n497), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n515), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n517), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n482), .B1(new_n516), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n494), .A2(KEYINPUT83), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(new_n497), .A3(new_n486), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n515), .B1(new_n531), .B2(new_n518), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n529), .B1(new_n532), .B2(new_n482), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n528), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n479), .A2(new_n481), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT17), .B1(new_n498), .B2(new_n515), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n525), .A2(new_n517), .A3(new_n526), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n535), .B1(new_n541), .B2(new_n533), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n529), .B(KEYINPUT13), .Z(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n525), .A2(new_n526), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n538), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n532), .A2(new_n482), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n537), .A2(new_n542), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G197gat), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT11), .B(G169gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT12), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n540), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n533), .B1(new_n558), .B2(new_n482), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n548), .B1(new_n559), .B2(new_n536), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(new_n555), .A3(new_n542), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT88), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT41), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(KEYINPUT95), .A2(G99gat), .A3(G106gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(KEYINPUT8), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G99gat), .ZN(new_n573));
  INV_X1    g372(.A(G106gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n568), .ZN(new_n576));
  OAI21_X1  g375(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n577));
  AND2_X1   g376(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT7), .ZN(new_n580));
  INV_X1    g379(.A(G85gat), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n580), .A2(new_n581), .A3(G92gat), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n572), .B(new_n576), .C1(new_n579), .C2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n580), .A2(new_n581), .ZN(new_n585));
  NAND2_X1  g384(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(G92gat), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n577), .A2(new_n578), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n576), .B1(new_n589), .B2(new_n572), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n567), .B1(new_n545), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n558), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n593), .B2(new_n591), .ZN(new_n594));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n565), .A2(new_n566), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT93), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT94), .ZN(new_n601));
  XOR2_X1   g400(.A(G134gat), .B(G162gat), .Z(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n597), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n594), .A2(new_n595), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n603), .B1(new_n606), .B2(new_n596), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G71gat), .B(G78gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT89), .ZN(new_n610));
  OR2_X1    g409(.A1(G71gat), .A2(G78gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT89), .ZN(new_n612));
  NAND2_X1  g411(.A1(G71gat), .A2(G78gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n615));
  INV_X1    g414(.A(G57gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(G64gat), .ZN(new_n617));
  INV_X1    g416(.A(G64gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(G57gat), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n615), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n610), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G57gat), .B(G64gat), .ZN(new_n622));
  OAI211_X1 g421(.A(KEYINPUT89), .B(new_n609), .C1(new_n622), .C2(new_n615), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n482), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n294), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n635));
  NAND3_X1  g434(.A1(new_n621), .A2(new_n635), .A3(new_n623), .ZN(new_n636));
  AND2_X1   g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(G127gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(G183gat), .B(G211gat), .Z(new_n643));
  NOR2_X1   g442(.A1(new_n640), .A2(G127gat), .ZN(new_n644));
  OR3_X1    g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n642), .B2(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n634), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n632), .A2(new_n646), .A3(new_n645), .A4(new_n633), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT97), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G230gat), .A2(G233gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT98), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n623), .B(new_n621), .C1(new_n584), .C2(new_n590), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT10), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n572), .B1(new_n579), .B2(new_n582), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(new_n568), .A3(new_n575), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n624), .A2(new_n660), .A3(new_n583), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n591), .A2(KEYINPUT10), .A3(new_n624), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n656), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n655), .B1(new_n657), .B2(new_n661), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n654), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT99), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n668), .B(new_n654), .C1(new_n664), .C2(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n655), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n662), .B2(new_n663), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n654), .B1(new_n665), .B2(KEYINPUT96), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n673), .B(new_n674), .C1(KEYINPUT96), .C2(new_n665), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n608), .A2(new_n650), .A3(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n470), .A2(new_n564), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n342), .A2(new_n343), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n426), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n473), .A2(new_n478), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n478), .B2(new_n684), .ZN(new_n688));
  MUX2_X1   g487(.A(new_n687), .B(new_n688), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g488(.A(new_n679), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n425), .A2(new_n421), .ZN(new_n691));
  OAI21_X1  g490(.A(G15gat), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n465), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(G15gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n690), .B2(new_n694), .ZN(G1326gat));
  NOR2_X1   g494(.A1(new_n470), .A2(new_n564), .ZN(new_n696));
  INV_X1    g495(.A(new_n459), .ZN(new_n697));
  INV_X1    g496(.A(new_n678), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  NOR3_X1   g500(.A1(new_n608), .A2(new_n650), .A3(new_n676), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n696), .A2(new_n500), .A3(new_n680), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT44), .B1(new_n470), .B2(new_n608), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n464), .A2(new_n469), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n441), .A2(new_n457), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n386), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n344), .A2(new_n380), .A3(new_n385), .A4(KEYINPUT101), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n691), .A2(new_n707), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n604), .B1(new_n597), .B2(new_n598), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n606), .A2(new_n603), .A3(new_n596), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n716));
  NAND3_X1  g515(.A1(new_n712), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n705), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n650), .B(KEYINPUT100), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n555), .B1(new_n560), .B2(new_n542), .ZN(new_n720));
  AND4_X1   g519(.A1(new_n555), .A2(new_n537), .A3(new_n542), .A4(new_n549), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n719), .A2(new_n722), .A3(new_n676), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n680), .ZN(new_n725));
  OAI21_X1  g524(.A(G29gat), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n704), .A2(new_n726), .ZN(G1328gat));
  AND2_X1   g526(.A1(new_n696), .A2(new_n702), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n729));
  AOI21_X1  g528(.A(G36gat), .B1(new_n729), .B2(KEYINPUT46), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n426), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n729), .A2(KEYINPUT46), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G36gat), .B1(new_n724), .B2(new_n285), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1329gat));
  NAND2_X1  g534(.A1(new_n505), .A2(new_n507), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n728), .A2(new_n465), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n724), .A2(new_n691), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(new_n737), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g541(.A(KEYINPUT47), .B(new_n738), .C1(new_n739), .C2(new_n737), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1330gat));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n508), .A3(new_n697), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(KEYINPUT48), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT104), .B1(new_n724), .B2(new_n459), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G50gat), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n724), .A2(KEYINPUT104), .A3(new_n459), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n724), .A2(new_n459), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n745), .B1(new_n751), .B2(new_n508), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT48), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(new_n754), .ZN(G1331gat));
  NAND4_X1  g554(.A1(new_n608), .A2(new_n722), .A3(new_n650), .A4(new_n676), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n706), .B2(new_n711), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n680), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g558(.A1(new_n757), .A2(new_n426), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  AND2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n760), .B2(new_n761), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT105), .ZN(G1333gat));
  INV_X1    g564(.A(new_n691), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n407), .B1(new_n757), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n693), .A2(G71gat), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n757), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g569(.A1(new_n757), .A2(new_n697), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g571(.A(new_n608), .B1(new_n706), .B2(new_n711), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n650), .A2(new_n562), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(KEYINPUT51), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT51), .B1(new_n773), .B2(new_n774), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n676), .A2(new_n581), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n778), .A2(new_n725), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n774), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n677), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n705), .B2(new_n717), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n581), .B1(new_n784), .B2(new_n680), .ZN(new_n785));
  OR3_X1    g584(.A1(new_n780), .A2(new_n785), .A3(KEYINPUT106), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT106), .B1(new_n780), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1336gat));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  INV_X1    g588(.A(G92gat), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n784), .B2(new_n426), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n677), .A2(new_n285), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n790), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n712), .A2(new_n715), .A3(new_n774), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n795), .B1(new_n798), .B2(new_n775), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n791), .A2(KEYINPUT108), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT108), .ZN(new_n801));
  INV_X1    g600(.A(new_n716), .ZN(new_n802));
  AOI211_X1 g601(.A(new_n608), .B(new_n802), .C1(new_n706), .C2(new_n711), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n691), .A2(new_n707), .A3(new_n386), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n706), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n806), .B2(new_n715), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n426), .B(new_n782), .C1(new_n803), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G92gat), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n790), .B(new_n794), .C1(new_n776), .C2(new_n777), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n801), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n793), .B1(new_n800), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT108), .B1(new_n791), .B2(new_n799), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(new_n809), .B2(KEYINPUT107), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n809), .A2(new_n810), .A3(new_n801), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n816), .ZN(G1337gat));
  INV_X1    g616(.A(new_n784), .ZN(new_n818));
  OAI21_X1  g617(.A(G99gat), .B1(new_n818), .B2(new_n691), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n465), .A2(new_n573), .A3(new_n676), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n778), .B2(new_n820), .ZN(G1338gat));
  NAND2_X1  g620(.A1(new_n676), .A2(new_n574), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n778), .A2(new_n459), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n574), .B1(new_n784), .B2(new_n697), .ZN(new_n824));
  OR3_X1    g623(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT53), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT53), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1339gat));
  INV_X1    g626(.A(G113gat), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n725), .A2(new_n426), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n465), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n831));
  OR3_X1    g630(.A1(new_n678), .A2(KEYINPUT109), .A3(new_n562), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT109), .B1(new_n678), .B2(new_n562), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n529), .B1(new_n528), .B2(new_n546), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n546), .A2(new_n547), .A3(new_n544), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n554), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n676), .A2(new_n561), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n672), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n662), .A2(new_n663), .A3(new_n656), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g642(.A(KEYINPUT54), .B(new_n656), .C1(new_n662), .C2(new_n663), .ZN(new_n844));
  INV_X1    g643(.A(new_n654), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n844), .A2(KEYINPUT110), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n662), .A2(new_n663), .ZN(new_n848));
  INV_X1    g647(.A(new_n656), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n840), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n847), .B1(new_n850), .B2(new_n654), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n843), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n842), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n672), .A3(new_n840), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT110), .B1(new_n844), .B2(new_n845), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n850), .A2(new_n847), .A3(new_n654), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n852), .B(new_n675), .C1(new_n857), .C2(KEYINPUT55), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n838), .B1(new_n858), .B2(new_n722), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT111), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n861), .B(new_n838), .C1(new_n858), .C2(new_n722), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n608), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n561), .A2(new_n837), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n608), .A2(new_n858), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n719), .B1(new_n867), .B2(KEYINPUT112), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n715), .B1(new_n859), .B2(KEYINPUT111), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n865), .B1(new_n869), .B2(new_n862), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT112), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n834), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n831), .B1(new_n873), .B2(new_n697), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n832), .A2(new_n833), .ZN(new_n875));
  INV_X1    g674(.A(new_n719), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n870), .B2(new_n871), .ZN(new_n877));
  AOI211_X1 g676(.A(KEYINPUT112), .B(new_n865), .C1(new_n869), .C2(new_n862), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(KEYINPUT113), .A3(new_n459), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n830), .B1(new_n874), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n828), .B1(new_n881), .B2(new_n563), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n722), .A2(G113gat), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n693), .A2(new_n697), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n879), .A2(new_n680), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT114), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n879), .A2(new_n888), .A3(new_n680), .A4(new_n885), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n426), .B(new_n884), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT115), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n830), .ZN(new_n892));
  INV_X1    g691(.A(new_n880), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT113), .B1(new_n879), .B2(new_n459), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n563), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G113gat), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n887), .A2(new_n889), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n285), .A3(new_n883), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n891), .A2(new_n900), .ZN(G1340gat));
  NOR2_X1   g700(.A1(new_n677), .A2(G120gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n897), .A2(new_n285), .A3(new_n902), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n676), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n904), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT116), .B1(new_n904), .B2(G120gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(G1341gat));
  INV_X1    g706(.A(G127gat), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n897), .A2(new_n908), .A3(new_n285), .A4(new_n650), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n881), .A2(new_n719), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n908), .ZN(G1342gat));
  OAI211_X1 g710(.A(new_n715), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n608), .A2(G134gat), .A3(new_n426), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n887), .B2(new_n889), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n916));
  AOI22_X1  g715(.A1(G134gat), .A2(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n897), .A2(new_n913), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT117), .B1(new_n918), .B2(KEYINPUT56), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n915), .A2(new_n920), .A3(new_n916), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n919), .B2(new_n921), .ZN(G1343gat));
  NAND2_X1  g721(.A1(new_n691), .A2(new_n829), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT118), .ZN(new_n924));
  XOR2_X1   g723(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n925));
  AOI21_X1  g724(.A(new_n925), .B1(new_n879), .B2(new_n697), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n648), .A2(new_n649), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n677), .A2(new_n864), .ZN(new_n928));
  INV_X1    g727(.A(new_n858), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n563), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n866), .B1(new_n930), .B2(new_n715), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n834), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n932), .A2(new_n933), .A3(new_n459), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n924), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G141gat), .B1(new_n935), .B2(new_n564), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n766), .A2(new_n459), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n285), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n873), .A2(new_n725), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n563), .A2(new_n290), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT120), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT58), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n936), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT58), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n562), .B(new_n924), .C1(new_n926), .C2(new_n934), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n945), .A2(G141gat), .B1(new_n939), .B2(new_n941), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(G1344gat));
  NAND4_X1  g746(.A1(new_n939), .A2(new_n287), .A3(new_n288), .A4(new_n676), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n948), .B(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT59), .B1(new_n287), .B2(new_n288), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n951), .B1(new_n935), .B2(new_n677), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT59), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n678), .A2(new_n563), .A3(KEYINPUT122), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n698), .B2(new_n564), .ZN(new_n956));
  AOI211_X1 g755(.A(new_n954), .B(new_n956), .C1(new_n931), .C2(new_n927), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n933), .B1(new_n957), .B2(new_n459), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n879), .A2(new_n697), .A3(new_n925), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n924), .A2(new_n676), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n299), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n952), .B1(new_n953), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n950), .A2(new_n963), .ZN(G1345gat));
  OAI21_X1  g763(.A(G155gat), .B1(new_n935), .B2(new_n876), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n939), .A2(new_n294), .A3(new_n650), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1346gat));
  OAI21_X1  g766(.A(G162gat), .B1(new_n935), .B2(new_n608), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n939), .A2(new_n295), .A3(new_n715), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1347gat));
  NOR2_X1   g769(.A1(new_n873), .A2(new_n680), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(new_n885), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n972), .A2(new_n426), .A3(new_n562), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n680), .A2(new_n285), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT123), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(new_n465), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n977), .B1(new_n874), .B2(new_n880), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n564), .A2(new_n207), .ZN(new_n979));
  AOI22_X1  g778(.A1(new_n973), .A2(new_n207), .B1(new_n978), .B2(new_n979), .ZN(G1348gat));
  NAND3_X1  g779(.A1(new_n972), .A2(new_n208), .A3(new_n794), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n978), .A2(new_n676), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(new_n208), .ZN(G1349gat));
  AOI21_X1  g782(.A(new_n215), .B1(new_n978), .B2(new_n719), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n971), .A2(new_n426), .A3(new_n885), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n985), .A2(new_n219), .A3(new_n927), .ZN(new_n986));
  OAI21_X1  g785(.A(KEYINPUT60), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  OR3_X1    g786(.A1(new_n985), .A2(new_n219), .A3(new_n927), .ZN(new_n988));
  INV_X1    g787(.A(new_n977), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n719), .B(new_n989), .C1(new_n893), .C2(new_n894), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(G183gat), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT60), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n987), .A2(new_n993), .ZN(G1350gat));
  NOR2_X1   g793(.A1(new_n608), .A2(G190gat), .ZN(new_n995));
  INV_X1    g794(.A(new_n995), .ZN(new_n996));
  OR3_X1    g795(.A1(new_n985), .A2(KEYINPUT124), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g796(.A(KEYINPUT124), .B1(new_n985), .B2(new_n996), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g798(.A(new_n715), .B(new_n989), .C1(new_n893), .C2(new_n894), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(G190gat), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT61), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1000), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n999), .A2(new_n1003), .A3(new_n1004), .ZN(G1351gat));
  AND3_X1   g804(.A1(new_n879), .A2(new_n725), .A3(new_n937), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n1006), .A2(new_n426), .ZN(new_n1007));
  AOI21_X1  g806(.A(G197gat), .B1(new_n1007), .B2(new_n562), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n976), .A2(new_n691), .ZN(new_n1009));
  XNOR2_X1  g808(.A(new_n1009), .B(KEYINPUT125), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1010), .B1(new_n958), .B2(new_n959), .ZN(new_n1011));
  AND3_X1   g810(.A1(new_n1011), .A2(G197gat), .A3(new_n563), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n1008), .A2(new_n1012), .ZN(G1352gat));
  INV_X1    g812(.A(G204gat), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1006), .A2(new_n1014), .A3(new_n794), .ZN(new_n1015));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1016));
  XNOR2_X1  g815(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  AOI211_X1 g816(.A(new_n677), .B(new_n1010), .C1(new_n958), .C2(new_n959), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT126), .ZN(new_n1019));
  AND2_X1   g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g819(.A(G204gat), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1021));
  OAI21_X1  g820(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(G1353gat));
  NAND3_X1  g821(.A1(new_n1007), .A2(new_n259), .A3(new_n650), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1011), .A2(new_n650), .ZN(new_n1024));
  AOI21_X1  g823(.A(KEYINPUT63), .B1(new_n1024), .B2(G211gat), .ZN(new_n1025));
  INV_X1    g824(.A(KEYINPUT63), .ZN(new_n1026));
  AOI211_X1 g825(.A(new_n1026), .B(new_n259), .C1(new_n1011), .C2(new_n650), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1023), .B1(new_n1025), .B2(new_n1027), .ZN(G1354gat));
  INV_X1    g827(.A(new_n1010), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n960), .A2(KEYINPUT127), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1030), .A2(new_n715), .ZN(new_n1031));
  NOR2_X1   g830(.A1(new_n1011), .A2(KEYINPUT127), .ZN(new_n1032));
  OAI21_X1  g831(.A(G218gat), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n1007), .A2(new_n260), .A3(new_n715), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n1033), .A2(new_n1034), .ZN(G1355gat));
endmodule


