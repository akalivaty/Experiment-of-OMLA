

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U558 ( .A(n881), .Z(n524) );
  NOR2_X1 U559 ( .A1(n774), .A2(n765), .ZN(n525) );
  INV_X1 U560 ( .A(KEYINPUT30), .ZN(n738) );
  INV_X1 U561 ( .A(n974), .ZN(n765) );
  NOR2_X1 U562 ( .A1(n703), .A2(n702), .ZN(n730) );
  AND2_X1 U563 ( .A1(n766), .A2(n525), .ZN(n767) );
  NOR2_X1 U564 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U565 ( .A1(G164), .A2(G1384), .ZN(n701) );
  XOR2_X1 U566 ( .A(KEYINPUT77), .B(n611), .Z(n970) );
  NOR2_X1 U567 ( .A1(G651), .A2(n657), .ZN(n667) );
  NOR2_X1 U568 ( .A1(n537), .A2(n536), .ZN(G160) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n880) );
  NAND2_X1 U570 ( .A1(n880), .A2(G113), .ZN(n528) );
  INV_X1 U571 ( .A(G2104), .ZN(n529) );
  NOR2_X2 U572 ( .A1(G2105), .A2(n529), .ZN(n876) );
  NAND2_X1 U573 ( .A1(G101), .A2(n876), .ZN(n526) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n526), .Z(n527) );
  NAND2_X1 U575 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U576 ( .A1(n529), .A2(G2105), .ZN(n530) );
  XNOR2_X1 U577 ( .A(n530), .B(KEYINPUT65), .ZN(n881) );
  NAND2_X1 U578 ( .A1(n524), .A2(G125), .ZN(n535) );
  XNOR2_X1 U579 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n532) );
  NOR2_X1 U580 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X2 U582 ( .A(KEYINPUT66), .B(n533), .ZN(n877) );
  NAND2_X1 U583 ( .A1(G137), .A2(n877), .ZN(n534) );
  NAND2_X1 U584 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U585 ( .A1(G651), .A2(G543), .ZN(n538) );
  XNOR2_X1 U586 ( .A(n538), .B(KEYINPUT64), .ZN(n664) );
  NAND2_X1 U587 ( .A1(n664), .A2(G89), .ZN(n539) );
  XNOR2_X1 U588 ( .A(n539), .B(KEYINPUT78), .ZN(n540) );
  XNOR2_X1 U589 ( .A(n540), .B(KEYINPUT4), .ZN(n542) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n657) );
  INV_X1 U591 ( .A(G651), .ZN(n544) );
  NOR2_X1 U592 ( .A1(n657), .A2(n544), .ZN(n663) );
  NAND2_X1 U593 ( .A1(G76), .A2(n663), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U595 ( .A(n543), .B(KEYINPUT5), .ZN(n552) );
  NAND2_X1 U596 ( .A1(G51), .A2(n667), .ZN(n549) );
  INV_X1 U597 ( .A(KEYINPUT68), .ZN(n547) );
  NOR2_X1 U598 ( .A1(G543), .A2(n544), .ZN(n545) );
  XNOR2_X1 U599 ( .A(KEYINPUT1), .B(n545), .ZN(n546) );
  XNOR2_X2 U600 ( .A(n547), .B(n546), .ZN(n668) );
  NAND2_X1 U601 ( .A1(G63), .A2(n668), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U603 ( .A(KEYINPUT6), .B(n550), .Z(n551) );
  NAND2_X1 U604 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U605 ( .A(n553), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U606 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U607 ( .A1(G102), .A2(n876), .ZN(n555) );
  NAND2_X1 U608 ( .A1(G138), .A2(n877), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U610 ( .A1(G114), .A2(n880), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G126), .A2(n524), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U613 ( .A1(n559), .A2(n558), .ZN(G164) );
  XOR2_X1 U614 ( .A(G2451), .B(G2454), .Z(n561) );
  XNOR2_X1 U615 ( .A(G2430), .B(KEYINPUT104), .ZN(n560) );
  XNOR2_X1 U616 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U617 ( .A(n562), .B(G2446), .Z(n564) );
  XNOR2_X1 U618 ( .A(G1348), .B(G1341), .ZN(n563) );
  XNOR2_X1 U619 ( .A(n564), .B(n563), .ZN(n568) );
  XOR2_X1 U620 ( .A(G2438), .B(G2427), .Z(n566) );
  XNOR2_X1 U621 ( .A(G2443), .B(G2435), .ZN(n565) );
  XNOR2_X1 U622 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U623 ( .A(n568), .B(n567), .Z(n569) );
  AND2_X1 U624 ( .A1(G14), .A2(n569), .ZN(G401) );
  AND2_X1 U625 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U626 ( .A1(G99), .A2(n876), .ZN(n571) );
  NAND2_X1 U627 ( .A1(G111), .A2(n880), .ZN(n570) );
  NAND2_X1 U628 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U629 ( .A(KEYINPUT82), .B(n572), .ZN(n575) );
  NAND2_X1 U630 ( .A1(n524), .A2(G123), .ZN(n573) );
  XOR2_X1 U631 ( .A(KEYINPUT18), .B(n573), .Z(n574) );
  NOR2_X1 U632 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U633 ( .A1(G135), .A2(n877), .ZN(n576) );
  NAND2_X1 U634 ( .A1(n577), .A2(n576), .ZN(n941) );
  XOR2_X1 U635 ( .A(G2096), .B(KEYINPUT83), .Z(n578) );
  XNOR2_X1 U636 ( .A(n941), .B(n578), .ZN(n579) );
  OR2_X1 U637 ( .A1(G2100), .A2(n579), .ZN(G156) );
  INV_X1 U638 ( .A(G132), .ZN(G219) );
  INV_X1 U639 ( .A(G82), .ZN(G220) );
  INV_X1 U640 ( .A(G120), .ZN(G236) );
  INV_X1 U641 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U642 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n584) );
  NAND2_X1 U643 ( .A1(n663), .A2(G77), .ZN(n581) );
  NAND2_X1 U644 ( .A1(G90), .A2(n664), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT9), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n584), .B(n583), .ZN(n589) );
  NAND2_X1 U648 ( .A1(n667), .A2(G52), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT70), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G64), .A2(n668), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U652 ( .A1(n589), .A2(n588), .ZN(G171) );
  NAND2_X1 U653 ( .A1(G7), .A2(G661), .ZN(n590) );
  XOR2_X1 U654 ( .A(n590), .B(KEYINPUT10), .Z(n831) );
  NAND2_X1 U655 ( .A1(n831), .A2(G567), .ZN(n591) );
  XOR2_X1 U656 ( .A(KEYINPUT11), .B(n591), .Z(G234) );
  NAND2_X1 U657 ( .A1(n664), .A2(G81), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n592), .B(KEYINPUT12), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n593), .B(KEYINPUT74), .ZN(n595) );
  NAND2_X1 U660 ( .A1(G68), .A2(n663), .ZN(n594) );
  NAND2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U662 ( .A(n596), .B(KEYINPUT13), .ZN(n598) );
  NAND2_X1 U663 ( .A1(G43), .A2(n667), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U665 ( .A1(n668), .A2(G56), .ZN(n599) );
  XOR2_X1 U666 ( .A(KEYINPUT14), .B(n599), .Z(n600) );
  NOR2_X1 U667 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U668 ( .A(KEYINPUT75), .B(n602), .Z(n982) );
  NAND2_X1 U669 ( .A1(n982), .A2(G860), .ZN(G153) );
  INV_X1 U670 ( .A(G171), .ZN(G301) );
  NAND2_X1 U671 ( .A1(G868), .A2(G301), .ZN(n613) );
  NAND2_X1 U672 ( .A1(G92), .A2(n664), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G66), .A2(n668), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U675 ( .A(KEYINPUT76), .B(n605), .ZN(n609) );
  NAND2_X1 U676 ( .A1(G79), .A2(n663), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G54), .A2(n667), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U679 ( .A(KEYINPUT15), .B(n610), .Z(n611) );
  INV_X1 U680 ( .A(n970), .ZN(n713) );
  INV_X1 U681 ( .A(G868), .ZN(n683) );
  NAND2_X1 U682 ( .A1(n713), .A2(n683), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n613), .A2(n612), .ZN(G284) );
  NAND2_X1 U684 ( .A1(n663), .A2(G78), .ZN(n615) );
  NAND2_X1 U685 ( .A1(G91), .A2(n664), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U687 ( .A1(G53), .A2(n667), .ZN(n616) );
  XNOR2_X1 U688 ( .A(KEYINPUT73), .B(n616), .ZN(n617) );
  NOR2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G65), .A2(n668), .ZN(n619) );
  NAND2_X1 U691 ( .A1(n620), .A2(n619), .ZN(G299) );
  NOR2_X1 U692 ( .A1(G286), .A2(n683), .ZN(n621) );
  XOR2_X1 U693 ( .A(KEYINPUT79), .B(n621), .Z(n623) );
  NOR2_X1 U694 ( .A1(G868), .A2(G299), .ZN(n622) );
  NOR2_X1 U695 ( .A1(n623), .A2(n622), .ZN(G297) );
  INV_X1 U696 ( .A(G860), .ZN(n632) );
  NAND2_X1 U697 ( .A1(n632), .A2(G559), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n624), .A2(n970), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n625), .B(KEYINPUT81), .ZN(n627) );
  XOR2_X1 U700 ( .A(KEYINPUT16), .B(KEYINPUT80), .Z(n626) );
  XNOR2_X1 U701 ( .A(n627), .B(n626), .ZN(G148) );
  NOR2_X1 U702 ( .A1(G559), .A2(n713), .ZN(n628) );
  NOR2_X1 U703 ( .A1(n683), .A2(n628), .ZN(n630) );
  NOR2_X1 U704 ( .A1(n982), .A2(G868), .ZN(n629) );
  OR2_X1 U705 ( .A1(n630), .A2(n629), .ZN(G282) );
  NAND2_X1 U706 ( .A1(G559), .A2(n970), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n631), .B(n982), .ZN(n679) );
  NAND2_X1 U708 ( .A1(n632), .A2(n679), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n663), .A2(G80), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G93), .A2(n664), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G55), .A2(n667), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G67), .A2(n668), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n682) );
  XOR2_X1 U716 ( .A(n639), .B(n682), .Z(G145) );
  NAND2_X1 U717 ( .A1(G47), .A2(n667), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G60), .A2(n668), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U720 ( .A1(n663), .A2(G72), .ZN(n643) );
  NAND2_X1 U721 ( .A1(G85), .A2(n664), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n646), .B(KEYINPUT69), .ZN(G290) );
  NAND2_X1 U725 ( .A1(n663), .A2(G73), .ZN(n648) );
  XNOR2_X1 U726 ( .A(KEYINPUT2), .B(KEYINPUT86), .ZN(n647) );
  XNOR2_X1 U727 ( .A(n648), .B(n647), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n667), .A2(G48), .ZN(n650) );
  NAND2_X1 U729 ( .A1(G86), .A2(n664), .ZN(n649) );
  NAND2_X1 U730 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U731 ( .A1(G61), .A2(n668), .ZN(n651) );
  XNOR2_X1 U732 ( .A(KEYINPUT85), .B(n651), .ZN(n652) );
  NOR2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n655), .A2(n654), .ZN(G305) );
  NAND2_X1 U735 ( .A1(G49), .A2(n667), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(KEYINPUT84), .ZN(n662) );
  NAND2_X1 U737 ( .A1(G87), .A2(n657), .ZN(n659) );
  NAND2_X1 U738 ( .A1(G74), .A2(G651), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U740 ( .A1(n668), .A2(n660), .ZN(n661) );
  NAND2_X1 U741 ( .A1(n662), .A2(n661), .ZN(G288) );
  NAND2_X1 U742 ( .A1(n663), .A2(G75), .ZN(n666) );
  NAND2_X1 U743 ( .A1(G88), .A2(n664), .ZN(n665) );
  NAND2_X1 U744 ( .A1(n666), .A2(n665), .ZN(n672) );
  NAND2_X1 U745 ( .A1(G50), .A2(n667), .ZN(n670) );
  NAND2_X1 U746 ( .A1(G62), .A2(n668), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U748 ( .A1(n672), .A2(n671), .ZN(G166) );
  INV_X1 U749 ( .A(G166), .ZN(G303) );
  XOR2_X1 U750 ( .A(G299), .B(G290), .Z(n673) );
  XNOR2_X1 U751 ( .A(n673), .B(G305), .ZN(n676) );
  XOR2_X1 U752 ( .A(KEYINPUT19), .B(KEYINPUT87), .Z(n674) );
  XNOR2_X1 U753 ( .A(G288), .B(n674), .ZN(n675) );
  XOR2_X1 U754 ( .A(n676), .B(n675), .Z(n678) );
  XOR2_X1 U755 ( .A(G303), .B(n682), .Z(n677) );
  XNOR2_X1 U756 ( .A(n678), .B(n677), .ZN(n900) );
  XNOR2_X1 U757 ( .A(n679), .B(n900), .ZN(n680) );
  XNOR2_X1 U758 ( .A(KEYINPUT88), .B(n680), .ZN(n681) );
  NOR2_X1 U759 ( .A1(n683), .A2(n681), .ZN(n685) );
  AND2_X1 U760 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U761 ( .A1(n685), .A2(n684), .ZN(G295) );
  NAND2_X1 U762 ( .A1(G2078), .A2(G2084), .ZN(n686) );
  XOR2_X1 U763 ( .A(KEYINPUT20), .B(n686), .Z(n687) );
  NAND2_X1 U764 ( .A1(G2090), .A2(n687), .ZN(n688) );
  XNOR2_X1 U765 ( .A(KEYINPUT21), .B(n688), .ZN(n689) );
  NAND2_X1 U766 ( .A1(n689), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U767 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U768 ( .A1(G237), .A2(G236), .ZN(n690) );
  NAND2_X1 U769 ( .A1(G69), .A2(n690), .ZN(n691) );
  XNOR2_X1 U770 ( .A(KEYINPUT89), .B(n691), .ZN(n692) );
  NAND2_X1 U771 ( .A1(n692), .A2(G108), .ZN(n836) );
  NAND2_X1 U772 ( .A1(G567), .A2(n836), .ZN(n697) );
  NOR2_X1 U773 ( .A1(G220), .A2(G219), .ZN(n693) );
  XOR2_X1 U774 ( .A(KEYINPUT22), .B(n693), .Z(n694) );
  NOR2_X1 U775 ( .A1(G218), .A2(n694), .ZN(n695) );
  NAND2_X1 U776 ( .A1(G96), .A2(n695), .ZN(n837) );
  NAND2_X1 U777 ( .A1(G2106), .A2(n837), .ZN(n696) );
  NAND2_X1 U778 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U779 ( .A(KEYINPUT90), .B(n698), .ZN(n835) );
  NAND2_X1 U780 ( .A1(G661), .A2(G483), .ZN(n699) );
  XOR2_X1 U781 ( .A(KEYINPUT91), .B(n699), .Z(n700) );
  NOR2_X1 U782 ( .A1(n835), .A2(n700), .ZN(n834) );
  NAND2_X1 U783 ( .A1(n834), .A2(G36), .ZN(G176) );
  XNOR2_X1 U784 ( .A(G1986), .B(G290), .ZN(n978) );
  NAND2_X1 U785 ( .A1(G160), .A2(G40), .ZN(n702) );
  NOR2_X1 U786 ( .A1(n701), .A2(n702), .ZN(n826) );
  NAND2_X1 U787 ( .A1(n978), .A2(n826), .ZN(n816) );
  INV_X1 U788 ( .A(n701), .ZN(n703) );
  INV_X1 U789 ( .A(n730), .ZN(n736) );
  INV_X1 U790 ( .A(G1996), .ZN(n852) );
  NOR2_X1 U791 ( .A1(n736), .A2(n852), .ZN(n705) );
  XOR2_X1 U792 ( .A(KEYINPUT26), .B(KEYINPUT102), .Z(n704) );
  XNOR2_X1 U793 ( .A(n705), .B(n704), .ZN(n707) );
  NAND2_X1 U794 ( .A1(n736), .A2(G1341), .ZN(n706) );
  NAND2_X1 U795 ( .A1(n707), .A2(n706), .ZN(n712) );
  NAND2_X1 U796 ( .A1(G1348), .A2(n736), .ZN(n709) );
  NAND2_X1 U797 ( .A1(G2067), .A2(n730), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n714) );
  NAND2_X1 U799 ( .A1(n713), .A2(n714), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n982), .A2(n710), .ZN(n711) );
  NOR2_X1 U801 ( .A1(n712), .A2(n711), .ZN(n716) );
  NOR2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U803 ( .A1(n716), .A2(n715), .ZN(n722) );
  NAND2_X1 U804 ( .A1(G2072), .A2(n730), .ZN(n717) );
  XOR2_X1 U805 ( .A(KEYINPUT99), .B(n717), .Z(n718) );
  XNOR2_X1 U806 ( .A(KEYINPUT27), .B(n718), .ZN(n720) );
  XOR2_X1 U807 ( .A(G1956), .B(KEYINPUT100), .Z(n999) );
  NOR2_X1 U808 ( .A1(n730), .A2(n999), .ZN(n719) );
  NOR2_X1 U809 ( .A1(n720), .A2(n719), .ZN(n723) );
  INV_X1 U810 ( .A(G299), .ZN(n965) );
  NAND2_X1 U811 ( .A1(n723), .A2(n965), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n727) );
  NOR2_X1 U813 ( .A1(n723), .A2(n965), .ZN(n725) );
  XNOR2_X1 U814 ( .A(KEYINPUT28), .B(KEYINPUT101), .ZN(n724) );
  XNOR2_X1 U815 ( .A(n725), .B(n724), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U817 ( .A(KEYINPUT29), .B(n728), .Z(n735) );
  XNOR2_X1 U818 ( .A(G2078), .B(KEYINPUT97), .ZN(n729) );
  XNOR2_X1 U819 ( .A(n729), .B(KEYINPUT25), .ZN(n922) );
  NOR2_X1 U820 ( .A1(n922), .A2(n736), .ZN(n732) );
  XNOR2_X1 U821 ( .A(G1961), .B(KEYINPUT96), .ZN(n1004) );
  NOR2_X1 U822 ( .A1(n730), .A2(n1004), .ZN(n731) );
  NOR2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n742) );
  NOR2_X1 U824 ( .A1(n742), .A2(G301), .ZN(n733) );
  XOR2_X1 U825 ( .A(KEYINPUT98), .B(n733), .Z(n734) );
  NAND2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n747) );
  NAND2_X1 U827 ( .A1(G8), .A2(n736), .ZN(n774) );
  NOR2_X1 U828 ( .A1(G1966), .A2(n774), .ZN(n758) );
  NOR2_X1 U829 ( .A1(G2084), .A2(n736), .ZN(n755) );
  NOR2_X1 U830 ( .A1(n758), .A2(n755), .ZN(n737) );
  AND2_X1 U831 ( .A1(n737), .A2(G8), .ZN(n739) );
  XNOR2_X1 U832 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U833 ( .A1(G168), .A2(n740), .ZN(n741) );
  XNOR2_X1 U834 ( .A(n741), .B(KEYINPUT103), .ZN(n744) );
  NAND2_X1 U835 ( .A1(n742), .A2(G301), .ZN(n743) );
  NAND2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U837 ( .A(n745), .B(KEYINPUT31), .ZN(n746) );
  NAND2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n756) );
  NAND2_X1 U839 ( .A1(n756), .A2(G286), .ZN(n752) );
  NOR2_X1 U840 ( .A1(G1971), .A2(n774), .ZN(n749) );
  NOR2_X1 U841 ( .A1(G2090), .A2(n736), .ZN(n748) );
  NOR2_X1 U842 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n750), .A2(G303), .ZN(n751) );
  NAND2_X1 U844 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U845 ( .A1(G8), .A2(n753), .ZN(n754) );
  XNOR2_X1 U846 ( .A(n754), .B(KEYINPUT32), .ZN(n762) );
  NAND2_X1 U847 ( .A1(G8), .A2(n755), .ZN(n760) );
  INV_X1 U848 ( .A(n756), .ZN(n757) );
  NOR2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n775) );
  NOR2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n973) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n763) );
  NOR2_X1 U854 ( .A1(n973), .A2(n763), .ZN(n764) );
  NAND2_X1 U855 ( .A1(n775), .A2(n764), .ZN(n766) );
  NAND2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NOR2_X1 U857 ( .A1(KEYINPUT33), .A2(n767), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n973), .A2(KEYINPUT33), .ZN(n768) );
  NOR2_X1 U859 ( .A1(n768), .A2(n774), .ZN(n769) );
  NOR2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U861 ( .A(G1981), .B(G305), .Z(n987) );
  NAND2_X1 U862 ( .A1(n771), .A2(n987), .ZN(n784) );
  NOR2_X1 U863 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XOR2_X1 U864 ( .A(n772), .B(KEYINPUT24), .Z(n773) );
  NOR2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n782) );
  INV_X1 U866 ( .A(n774), .ZN(n780) );
  INV_X1 U867 ( .A(n775), .ZN(n778) );
  NAND2_X1 U868 ( .A1(G166), .A2(G8), .ZN(n776) );
  NOR2_X1 U869 ( .A1(G2090), .A2(n776), .ZN(n777) );
  NOR2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n795) );
  XNOR2_X1 U874 ( .A(KEYINPUT37), .B(G2067), .ZN(n824) );
  NAND2_X1 U875 ( .A1(G104), .A2(n876), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G140), .A2(n877), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(n787), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G116), .A2(n880), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G128), .A2(n524), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U882 ( .A(KEYINPUT92), .B(n790), .Z(n791) );
  XNOR2_X1 U883 ( .A(KEYINPUT35), .B(n791), .ZN(n792) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U885 ( .A(KEYINPUT36), .B(n794), .ZN(n896) );
  NOR2_X1 U886 ( .A1(n824), .A2(n896), .ZN(n939) );
  NAND2_X1 U887 ( .A1(n826), .A2(n939), .ZN(n822) );
  NAND2_X1 U888 ( .A1(n795), .A2(n822), .ZN(n814) );
  NAND2_X1 U889 ( .A1(G107), .A2(n880), .ZN(n797) );
  NAND2_X1 U890 ( .A1(G119), .A2(n524), .ZN(n796) );
  NAND2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U892 ( .A(KEYINPUT93), .B(n798), .ZN(n803) );
  NAND2_X1 U893 ( .A1(G95), .A2(n876), .ZN(n800) );
  NAND2_X1 U894 ( .A1(G131), .A2(n877), .ZN(n799) );
  NAND2_X1 U895 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U896 ( .A(KEYINPUT94), .B(n801), .Z(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n888) );
  AND2_X1 U898 ( .A1(n888), .A2(G1991), .ZN(n812) );
  NAND2_X1 U899 ( .A1(G117), .A2(n880), .ZN(n805) );
  NAND2_X1 U900 ( .A1(G129), .A2(n524), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n876), .A2(G105), .ZN(n806) );
  XOR2_X1 U903 ( .A(KEYINPUT38), .B(n806), .Z(n807) );
  NOR2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n810) );
  NAND2_X1 U905 ( .A1(G141), .A2(n877), .ZN(n809) );
  NAND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n895) );
  AND2_X1 U907 ( .A1(n895), .A2(G1996), .ZN(n811) );
  OR2_X1 U908 ( .A1(n812), .A2(n811), .ZN(n940) );
  AND2_X1 U909 ( .A1(n940), .A2(n826), .ZN(n819) );
  XOR2_X1 U910 ( .A(KEYINPUT95), .B(n819), .Z(n813) );
  NOR2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n829) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n895), .ZN(n952) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U915 ( .A1(G1991), .A2(n888), .ZN(n944) );
  NOR2_X1 U916 ( .A1(n817), .A2(n944), .ZN(n818) );
  NOR2_X1 U917 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U918 ( .A1(n952), .A2(n820), .ZN(n821) );
  XNOR2_X1 U919 ( .A(KEYINPUT39), .B(n821), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n824), .A2(n896), .ZN(n948) );
  NAND2_X1 U922 ( .A1(n825), .A2(n948), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U925 ( .A(KEYINPUT40), .B(n830), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n831), .ZN(G217) );
  INV_X1 U927 ( .A(n831), .ZN(G223) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U929 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U931 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U932 ( .A(n835), .ZN(G319) );
  XNOR2_X1 U933 ( .A(G69), .B(KEYINPUT105), .ZN(G235) );
  INV_X1 U935 ( .A(G108), .ZN(G238) );
  INV_X1 U936 ( .A(G96), .ZN(G221) );
  NOR2_X1 U937 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XOR2_X1 U939 ( .A(G2096), .B(KEYINPUT43), .Z(n839) );
  XNOR2_X1 U940 ( .A(G2090), .B(KEYINPUT42), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U942 ( .A(n840), .B(G2678), .Z(n842) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U945 ( .A(KEYINPUT106), .B(G2100), .Z(n844) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U947 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1971), .B(G1956), .Z(n848) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1966), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U952 ( .A(n849), .B(KEYINPUT41), .Z(n851) );
  XNOR2_X1 U953 ( .A(G1961), .B(G1976), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n856) );
  XOR2_X1 U955 ( .A(G2474), .B(G1981), .Z(n854) );
  XOR2_X1 U956 ( .A(n852), .B(G1991), .Z(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G100), .A2(n876), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G112), .A2(n880), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G124), .A2(n524), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n859), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n877), .A2(G136), .ZN(n860) );
  XOR2_X1 U965 ( .A(KEYINPUT107), .B(n860), .Z(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U967 ( .A1(n864), .A2(n863), .ZN(G162) );
  XOR2_X1 U968 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n866) );
  XNOR2_X1 U969 ( .A(G164), .B(G160), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n894) );
  XNOR2_X1 U971 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G106), .A2(n876), .ZN(n868) );
  NAND2_X1 U973 ( .A1(G142), .A2(n877), .ZN(n867) );
  NAND2_X1 U974 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U975 ( .A(n869), .B(KEYINPUT45), .ZN(n870) );
  XNOR2_X1 U976 ( .A(n871), .B(n870), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G118), .A2(n880), .ZN(n873) );
  NAND2_X1 U978 ( .A1(G130), .A2(n524), .ZN(n872) );
  NAND2_X1 U979 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U980 ( .A1(n875), .A2(n874), .ZN(n892) );
  NAND2_X1 U981 ( .A1(G103), .A2(n876), .ZN(n879) );
  NAND2_X1 U982 ( .A1(G139), .A2(n877), .ZN(n878) );
  NAND2_X1 U983 ( .A1(n879), .A2(n878), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G115), .A2(n880), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G127), .A2(n524), .ZN(n882) );
  NAND2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(KEYINPUT47), .B(n884), .Z(n885) );
  NOR2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U989 ( .A(KEYINPUT110), .B(n887), .Z(n935) );
  XNOR2_X1 U990 ( .A(G162), .B(n888), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n889), .B(n941), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n935), .B(n890), .ZN(n891) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n898) );
  XOR2_X1 U995 ( .A(n896), .B(n895), .Z(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U997 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U998 ( .A(G286), .B(n900), .ZN(n902) );
  XOR2_X1 U999 ( .A(n970), .B(G171), .Z(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n903), .B(n982), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n904), .ZN(G397) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n905), .B(KEYINPUT49), .ZN(n906) );
  NOR2_X1 U1005 ( .A1(G401), .A2(n906), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(n907), .A2(G319), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(KEYINPUT111), .B(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(KEYINPUT112), .B(n911), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(KEYINPUT55), .ZN(n960) );
  XNOR2_X1 U1013 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n912) );
  XNOR2_X1 U1014 ( .A(n912), .B(G34), .ZN(n913) );
  XNOR2_X1 U1015 ( .A(G2084), .B(n913), .ZN(n929) );
  XNOR2_X1 U1016 ( .A(G2090), .B(G35), .ZN(n927) );
  XNOR2_X1 U1017 ( .A(G1991), .B(G25), .ZN(n915) );
  XNOR2_X1 U1018 ( .A(G33), .B(G2072), .ZN(n914) );
  NOR2_X1 U1019 ( .A1(n915), .A2(n914), .ZN(n921) );
  XOR2_X1 U1020 ( .A(G2067), .B(G26), .Z(n916) );
  NAND2_X1 U1021 ( .A1(n916), .A2(G28), .ZN(n919) );
  XNOR2_X1 U1022 ( .A(KEYINPUT116), .B(G1996), .ZN(n917) );
  XNOR2_X1 U1023 ( .A(G32), .B(n917), .ZN(n918) );
  NOR2_X1 U1024 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1025 ( .A1(n921), .A2(n920), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(G27), .B(n922), .ZN(n923) );
  NOR2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1028 ( .A(KEYINPUT53), .B(n925), .ZN(n926) );
  NOR2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(n930), .B(KEYINPUT118), .ZN(n931) );
  XOR2_X1 U1032 ( .A(n960), .B(n931), .Z(n932) );
  OR2_X1 U1033 ( .A1(G29), .A2(n932), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n933), .A2(G11), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(n934), .B(KEYINPUT119), .ZN(n964) );
  XOR2_X1 U1036 ( .A(G164), .B(G2078), .Z(n937) );
  XNOR2_X1 U1037 ( .A(G2072), .B(n935), .ZN(n936) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1039 ( .A(KEYINPUT50), .B(n938), .Z(n958) );
  OR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(G160), .B(G2084), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT113), .B(n945), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n955) );
  XOR2_X1 U1047 ( .A(G2090), .B(G162), .Z(n950) );
  XNOR2_X1 U1048 ( .A(KEYINPUT114), .B(n950), .ZN(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(KEYINPUT51), .B(n953), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT115), .B(n956), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(KEYINPUT52), .B(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n962), .A2(G29), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n1023) );
  INV_X1 U1058 ( .A(G16), .ZN(n1018) );
  XOR2_X1 U1059 ( .A(n1018), .B(KEYINPUT56), .Z(n993) );
  XOR2_X1 U1060 ( .A(G303), .B(G1971), .Z(n969) );
  XOR2_X1 U1061 ( .A(n965), .B(G1956), .Z(n967) );
  XOR2_X1 U1062 ( .A(G171), .B(G1961), .Z(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1065 ( .A(G1348), .B(n970), .Z(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n980) );
  INV_X1 U1067 ( .A(n973), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(KEYINPUT120), .B(n976), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(KEYINPUT121), .B(n981), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(n982), .B(G1341), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(n983), .B(KEYINPUT122), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(KEYINPUT123), .B(n986), .ZN(n991) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(KEYINPUT57), .B(n989), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n1020) );
  XNOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT59), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(n994), .B(G4), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(G6), .B(G1981), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1002) );
  XOR2_X1 U1088 ( .A(G20), .B(n999), .Z(n1000) );
  XNOR2_X1 U1089 ( .A(KEYINPUT124), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n1003), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(n1004), .B(G5), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(G21), .B(G1966), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1015) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G23), .B(G1976), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XOR2_X1 U1099 ( .A(G1986), .B(G24), .Z(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1106 ( .A(n1021), .B(KEYINPUT125), .Z(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(KEYINPUT126), .B(n1024), .Z(n1025) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

