//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0002(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0003(.A(G1), .ZN(new_n204));
  INV_X1    g0004(.A(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n205), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G244), .ZN(new_n216));
  AND2_X1   g0016(.A1(new_n216), .A2(G77), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n207), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n210), .B(new_n215), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT66), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G68), .B(G77), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(new_n236));
  XOR2_X1   g0036(.A(G50), .B(G58), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G200), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT3), .ZN(new_n244));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n250), .B1(new_n251), .B2(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n204), .A2(G274), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT68), .A2(G45), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT68), .A2(G45), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT70), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G41), .A2(G45), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(G1), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n204), .B(KEYINPUT70), .C1(G41), .C2(G45), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n255), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  XOR2_X1   g0067(.A(KEYINPUT69), .B(G226), .Z(new_n268));
  AOI21_X1  g0068(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n243), .B1(new_n256), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT75), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT9), .ZN(new_n273));
  INV_X1    g0073(.A(G50), .ZN(new_n274));
  INV_X1    g0074(.A(G58), .ZN(new_n275));
  INV_X1    g0075(.A(G68), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n277), .A2(G20), .B1(G150), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT71), .ZN(new_n281));
  OR3_X1    g0081(.A1(new_n275), .A2(KEYINPUT71), .A3(KEYINPUT8), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n205), .A2(G33), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n279), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n213), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n204), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n287), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n204), .A2(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G50), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n291), .A2(new_n294), .B1(new_n274), .B2(new_n290), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n273), .B1(new_n288), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n288), .A2(new_n273), .A3(new_n295), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n271), .A2(new_n272), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n256), .A2(new_n269), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n301), .A2(G190), .B1(new_n270), .B2(KEYINPUT75), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n271), .A2(new_n272), .B1(new_n305), .B2(new_n300), .ZN(new_n306));
  INV_X1    g0106(.A(new_n298), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n307), .A2(new_n296), .B1(new_n270), .B2(KEYINPUT75), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT10), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT72), .B(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n301), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n288), .A2(new_n295), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(G169), .C2(new_n301), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT68), .B(G45), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n204), .B(G274), .C1(new_n316), .C2(G41), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G97), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(G226), .A2(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(G232), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(G1698), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n319), .B1(new_n322), .B2(new_n248), .ZN(new_n323));
  INV_X1    g0123(.A(new_n213), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G41), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n317), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G238), .ZN(new_n328));
  AOI211_X1 g0128(.A(new_n328), .B(new_n255), .C1(new_n265), .C2(new_n266), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT13), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT76), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n321), .A2(G1698), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(G226), .B2(G1698), .ZN(new_n333));
  AND2_X1   g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NOR2_X1   g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n318), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n262), .B1(new_n337), .B2(new_n255), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT13), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n267), .A2(G238), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n330), .A2(new_n331), .A3(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n338), .A2(KEYINPUT76), .A3(new_n339), .A4(new_n340), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(G169), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT14), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n342), .A2(new_n346), .A3(G169), .A4(new_n343), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n330), .A2(G179), .A3(new_n341), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n278), .A2(G50), .B1(G20), .B2(new_n276), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n251), .B2(new_n284), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(KEYINPUT77), .A3(new_n287), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT77), .B1(new_n351), .B2(new_n287), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT11), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(new_n287), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT77), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT11), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(new_n352), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT12), .B1(new_n289), .B2(G68), .ZN(new_n361));
  OR3_X1    g0161(.A1(new_n289), .A2(KEYINPUT12), .A3(G68), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n276), .B1(new_n204), .B2(G20), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n361), .A2(new_n362), .B1(new_n291), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n355), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n349), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n330), .A2(G190), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n367), .B2(new_n341), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n342), .A2(G200), .A3(new_n343), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n246), .A2(new_n205), .A3(new_n247), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n246), .A2(KEYINPUT7), .A3(new_n205), .A4(new_n247), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n276), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n275), .A2(new_n276), .ZN(new_n379));
  NOR2_X1   g0179(.A1(G58), .A2(G68), .ZN(new_n380));
  OAI21_X1  g0180(.A(G20), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n278), .A2(G159), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n373), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT78), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n378), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n336), .B2(new_n205), .ZN(new_n388));
  INV_X1    g0188(.A(new_n377), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(KEYINPUT78), .A3(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n384), .A2(new_n387), .A3(new_n392), .A4(new_n287), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n281), .A2(new_n282), .A3(new_n292), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(KEYINPUT79), .ZN(new_n395));
  INV_X1    g0195(.A(new_n291), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n394), .B2(KEYINPUT79), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n395), .A2(new_n397), .B1(new_n290), .B2(new_n283), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT80), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n393), .A2(KEYINPUT80), .A3(new_n398), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n253), .A2(new_n249), .ZN(new_n403));
  INV_X1    g0203(.A(G226), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G1698), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n403), .B(new_n405), .C1(new_n334), .C2(new_n335), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G87), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n326), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(new_n262), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n267), .A2(G232), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G169), .ZN(new_n412));
  INV_X1    g0212(.A(new_n311), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n409), .A2(new_n413), .A3(new_n410), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n401), .A2(new_n402), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT18), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n321), .B(new_n255), .C1(new_n265), .C2(new_n266), .ZN(new_n418));
  NOR4_X1   g0218(.A1(new_n418), .A2(new_n408), .A3(new_n305), .A4(new_n262), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n243), .B1(new_n409), .B2(new_n410), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(new_n393), .A3(new_n398), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n421), .A2(new_n393), .A3(KEYINPUT17), .A4(new_n398), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n401), .A2(new_n427), .A3(new_n402), .A4(new_n415), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n417), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n336), .A2(G107), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n430), .B(new_n431), .C1(new_n252), .C2(new_n328), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n255), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n262), .B1(new_n267), .B2(new_n216), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n311), .ZN(new_n437));
  INV_X1    g0237(.A(new_n278), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n280), .A2(new_n438), .B1(new_n205), .B2(new_n251), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT15), .B(G87), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n284), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n287), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT73), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n442), .B(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n251), .B1(new_n204), .B2(G20), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n291), .A2(new_n445), .B1(new_n251), .B2(new_n290), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G169), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n435), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n437), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n435), .A2(G200), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(new_n444), .A3(new_n446), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(KEYINPUT74), .B1(G190), .B2(new_n436), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT74), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n451), .A2(new_n454), .A3(new_n444), .A4(new_n446), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n450), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g0257(.A1(new_n315), .A2(new_n372), .A3(new_n429), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT5), .B(G41), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n460), .A2(new_n462), .B1(new_n324), .B2(new_n325), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G257), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n460), .A2(G274), .A3(new_n462), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(G244), .B(new_n249), .C1(new_n334), .C2(new_n335), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT4), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT81), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n467), .A2(new_n468), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT81), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n467), .A2(new_n472), .A3(new_n468), .ZN(new_n473));
  OAI211_X1 g0273(.A(G250), .B(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n470), .A2(new_n471), .A3(new_n473), .A4(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n466), .B1(new_n477), .B2(new_n255), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT82), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n474), .B(new_n475), .C1(new_n467), .C2(new_n468), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n472), .B1(new_n467), .B2(new_n468), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n326), .B1(new_n483), .B2(new_n473), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT82), .B1(new_n484), .B2(new_n466), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n480), .A2(new_n485), .A3(G200), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n278), .A2(G77), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT6), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n488), .A2(new_n489), .A3(G107), .ZN(new_n490));
  XNOR2_X1  g0290(.A(G97), .B(G107), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n487), .B1(new_n492), .B2(new_n205), .ZN(new_n493));
  INV_X1    g0293(.A(G107), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n376), .B2(new_n377), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n287), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n289), .A2(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n204), .A2(G33), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n289), .A2(new_n498), .A3(new_n213), .A4(new_n286), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n497), .B1(new_n500), .B2(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n502), .B1(G190), .B2(new_n478), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n486), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n477), .A2(new_n255), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n466), .A2(new_n413), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n505), .A2(new_n506), .B1(new_n496), .B2(new_n501), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n448), .B1(new_n484), .B2(new_n466), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT88), .ZN(new_n511));
  AND2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  NOR2_X1   g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n462), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(new_n326), .A3(G264), .ZN(new_n515));
  INV_X1    g0315(.A(G294), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n245), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G250), .A2(G1698), .ZN(new_n518));
  INV_X1    g0318(.A(G257), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(G1698), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n517), .B1(new_n520), .B2(new_n248), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n465), .B(new_n515), .C1(new_n521), .C2(new_n326), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G169), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT86), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT87), .ZN(new_n526));
  INV_X1    g0326(.A(G179), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n519), .A2(G1698), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(G250), .B2(G1698), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n530), .A2(new_n336), .B1(new_n245), .B2(new_n516), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(new_n255), .B1(new_n463), .B2(G264), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(KEYINPUT87), .A3(G179), .A4(new_n465), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n522), .A2(KEYINPUT86), .A3(G169), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n525), .A2(new_n528), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT23), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n205), .B2(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n494), .A2(KEYINPUT23), .A3(G20), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n205), .A2(G33), .A3(G116), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n205), .B(G87), .C1(new_n334), .C2(new_n335), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT22), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT22), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n248), .A2(new_n544), .A3(new_n205), .A4(G87), .ZN(new_n545));
  AOI211_X1 g0345(.A(KEYINPUT24), .B(new_n541), .C1(new_n543), .C2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n543), .A2(new_n545), .ZN(new_n548));
  INV_X1    g0348(.A(new_n541), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n287), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n290), .A2(KEYINPUT25), .A3(new_n494), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT25), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n289), .B2(G107), .ZN(new_n554));
  AOI22_X1  g0354(.A1(G107), .A2(new_n500), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n511), .B1(new_n535), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n535), .A2(new_n556), .A3(new_n511), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n522), .A2(new_n243), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(G190), .B2(new_n522), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n551), .A3(new_n555), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G244), .B(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n564));
  OAI211_X1 g0364(.A(G238), .B(new_n249), .C1(new_n334), .C2(new_n335), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G116), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n255), .ZN(new_n568));
  OAI21_X1  g0368(.A(G250), .B1(new_n461), .B2(G1), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n255), .A2(new_n569), .B1(new_n461), .B2(new_n257), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G200), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n205), .B1(new_n318), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(G87), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(new_n489), .A3(new_n494), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n205), .B(G68), .C1(new_n334), .C2(new_n335), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n574), .B1(new_n284), .B2(new_n489), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n287), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n440), .A2(new_n290), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n500), .A2(G87), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n570), .B1(new_n567), .B2(new_n255), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G190), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n573), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n440), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n500), .A2(KEYINPUT83), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n499), .B2(new_n440), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n582), .A2(new_n590), .A3(new_n583), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n586), .A2(new_n311), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n593), .B(new_n594), .C1(G169), .C2(new_n586), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n588), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n500), .A2(G116), .ZN(new_n598));
  INV_X1    g0398(.A(G116), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n290), .A2(KEYINPUT84), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT84), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n289), .B2(G116), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n286), .A2(new_n213), .B1(G20), .B2(new_n599), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n475), .B(new_n205), .C1(G33), .C2(new_n489), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n604), .A2(KEYINPUT20), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT20), .B1(new_n604), .B2(new_n605), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n598), .B(new_n603), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n249), .A2(G264), .ZN(new_n609));
  NOR2_X1   g0409(.A1(G257), .A2(G1698), .ZN(new_n610));
  OAI22_X1  g0410(.A1(new_n609), .A2(new_n610), .B1(new_n334), .B2(new_n335), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(new_n255), .C1(G303), .C2(new_n248), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n514), .A2(new_n326), .A3(G270), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n465), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n608), .A2(KEYINPUT21), .A3(G169), .A4(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT85), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n613), .A2(new_n465), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n448), .B1(new_n618), .B2(new_n612), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n619), .A2(KEYINPUT85), .A3(KEYINPUT21), .A4(new_n608), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n608), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n618), .A2(G179), .A3(new_n612), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n622), .A2(new_n623), .B1(new_n625), .B2(new_n608), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n608), .B1(G200), .B2(new_n614), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n305), .B2(new_n614), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n597), .A2(new_n621), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  NOR4_X1   g0429(.A1(new_n459), .A2(new_n510), .A3(new_n563), .A4(new_n629), .ZN(G372));
  INV_X1    g0430(.A(new_n314), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n349), .A2(new_n365), .B1(new_n371), .B2(new_n450), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n424), .A2(new_n425), .ZN(new_n633));
  XNOR2_X1  g0433(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n399), .A2(new_n415), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n399), .B2(new_n415), .ZN(new_n636));
  OAI22_X1  g0436(.A1(new_n632), .A2(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n631), .B1(new_n637), .B2(new_n310), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n486), .A2(new_n503), .B1(new_n508), .B2(new_n507), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n535), .A2(new_n556), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n621), .A3(new_n626), .ZN(new_n641));
  INV_X1    g0441(.A(new_n562), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n596), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n639), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n507), .A2(new_n508), .A3(new_n595), .A4(new_n588), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT89), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n645), .A2(KEYINPUT89), .A3(new_n646), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n595), .B(new_n644), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n638), .B1(new_n459), .B2(new_n652), .ZN(G369));
  NAND2_X1  g0453(.A1(new_n621), .A2(new_n626), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n204), .A2(new_n205), .A3(G13), .ZN(new_n655));
  OAI21_X1  g0455(.A(G213), .B1(new_n655), .B2(KEYINPUT27), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(KEYINPUT27), .B2(new_n655), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT91), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT91), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(new_n608), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n654), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n621), .A2(new_n626), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n628), .ZN(new_n666));
  OAI211_X1 g0466(.A(KEYINPUT92), .B(new_n664), .C1(new_n666), .C2(new_n663), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n664), .A2(KEYINPUT92), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G330), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n535), .A2(new_n511), .A3(new_n556), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n671), .A2(new_n557), .A3(new_n642), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n556), .A2(new_n662), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n535), .A2(new_n556), .A3(new_n662), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n670), .A2(KEYINPUT93), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT93), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n669), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n662), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n654), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n672), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(new_n556), .A3(new_n535), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n208), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n204), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n577), .A2(G116), .ZN(new_n693));
  INV_X1    g0493(.A(new_n690), .ZN(new_n694));
  OAI22_X1  g0494(.A1(new_n692), .A2(new_n693), .B1(new_n211), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n645), .A2(new_n646), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT95), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT95), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n645), .B2(new_n646), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n698), .B(new_n595), .C1(new_n697), .C2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n558), .A2(new_n665), .A3(new_n559), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n702), .A2(new_n639), .A3(new_n643), .ZN(new_n703));
  OAI211_X1 g0503(.A(KEYINPUT29), .B(new_n682), .C1(new_n701), .C2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n652), .A2(new_n662), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(KEYINPUT29), .ZN(new_n706));
  NOR4_X1   g0506(.A1(new_n563), .A2(new_n510), .A3(new_n629), .A4(new_n662), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n662), .A2(KEYINPUT31), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n532), .A2(new_n586), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n624), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT30), .B1(new_n710), .B2(new_n478), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n572), .A2(new_n311), .A3(new_n614), .A4(new_n522), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n478), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT94), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(KEYINPUT30), .A3(new_n478), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n711), .A2(new_n713), .A3(KEYINPUT94), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n708), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  INV_X1    g0519(.A(new_n466), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n505), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n612), .A2(new_n465), .A3(new_n613), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(G179), .A3(new_n532), .A4(new_n586), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n719), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n478), .A2(new_n712), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(new_n725), .A3(new_n715), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n726), .B2(new_n662), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n718), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(G330), .B1(new_n707), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n706), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n696), .B1(new_n731), .B2(G1), .ZN(G364));
  NAND2_X1  g0532(.A1(new_n205), .A2(G13), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT96), .Z(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G45), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n691), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n670), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n667), .A2(new_n668), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n689), .A2(new_n336), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G355), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G116), .B2(new_n208), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n238), .A2(G45), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n689), .A2(new_n248), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n212), .B2(new_n260), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n749), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n213), .B1(G20), .B2(new_n448), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n744), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT97), .Z(new_n757));
  OAI21_X1  g0557(.A(new_n737), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n311), .A2(new_n205), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G190), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n305), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G322), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n759), .A2(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n205), .A2(G179), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n761), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n248), .B1(new_n769), .B2(G329), .ZN(new_n770));
  INV_X1    g0570(.A(G283), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n767), .A2(new_n305), .A3(G200), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n763), .A2(new_n527), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(G303), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n776), .A2(new_n516), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n766), .A2(new_n773), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G326), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n760), .A2(new_n305), .A3(G200), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT33), .B(G317), .Z(new_n784));
  OAI221_X1 g0584(.A(new_n780), .B1(new_n781), .B2(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n783), .A2(new_n276), .B1(new_n489), .B2(new_n776), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT99), .ZN(new_n787));
  INV_X1    g0587(.A(new_n782), .ZN(new_n788));
  INV_X1    g0588(.A(new_n777), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n336), .B1(new_n789), .B2(G87), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n788), .A2(G50), .B1(new_n790), .B2(KEYINPUT98), .ZN(new_n791));
  INV_X1    g0591(.A(new_n762), .ZN(new_n792));
  INV_X1    g0592(.A(new_n772), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n792), .A2(G77), .B1(G107), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n764), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT32), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n768), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n769), .A2(KEYINPUT32), .A3(G159), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n795), .A2(G58), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n791), .A2(new_n794), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n785), .B1(new_n787), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n758), .B1(new_n803), .B2(new_n755), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n738), .A2(new_n741), .B1(new_n746), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  NAND2_X1  g0606(.A1(new_n453), .A2(new_n455), .ZN(new_n807));
  INV_X1    g0607(.A(new_n450), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n447), .A2(new_n662), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT103), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n450), .A2(new_n811), .A3(new_n662), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n437), .A2(new_n447), .A3(new_n662), .A4(new_n449), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(KEYINPUT103), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n662), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n651), .A2(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n456), .A2(new_n809), .B1(new_n812), .B2(new_n814), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n817), .B1(new_n705), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n737), .B1(new_n820), .B2(new_n730), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n730), .B2(new_n820), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n755), .A2(new_n742), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n736), .B1(new_n251), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n788), .A2(G303), .B1(new_n792), .B2(G116), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n771), .B2(new_n783), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT100), .Z(new_n827));
  OAI21_X1  g0627(.A(new_n336), .B1(new_n768), .B2(new_n759), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G97), .B2(new_n775), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n789), .A2(G107), .B1(new_n793), .B2(G87), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n829), .B(new_n830), .C1(new_n516), .C2(new_n764), .ZN(new_n831));
  XOR2_X1   g0631(.A(KEYINPUT101), .B(G143), .Z(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G159), .A2(new_n792), .B1(new_n795), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  INV_X1    g0635(.A(G150), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n782), .C1(new_n836), .C2(new_n783), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT34), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n248), .B1(new_n768), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G68), .B2(new_n793), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G50), .A2(new_n789), .B1(new_n775), .B2(G58), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n839), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n837), .A2(new_n838), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n827), .A2(new_n831), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT102), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n755), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n846), .A2(new_n847), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n824), .B1(new_n743), .B2(new_n819), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n822), .A2(new_n851), .ZN(G384));
  INV_X1    g0652(.A(new_n492), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n214), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  OAI211_X1 g0657(.A(new_n212), .B(G77), .C1(new_n275), .C2(new_n276), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n274), .A2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n204), .B(G13), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(G330), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT40), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT104), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n393), .A2(new_n864), .A3(new_n398), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n864), .B1(new_n393), .B2(new_n398), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n415), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n660), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n865), .B2(new_n866), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n869), .A3(new_n422), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n422), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n401), .A2(new_n402), .A3(new_n868), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n416), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n869), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n429), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n393), .A2(KEYINPUT80), .A3(new_n398), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT80), .B1(new_n393), .B2(new_n398), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n881), .A2(new_n882), .A3(new_n660), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n635), .A2(new_n636), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(new_n633), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n874), .A2(new_n416), .A3(new_n875), .ZN(new_n886));
  INV_X1    g0686(.A(new_n422), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n393), .A2(new_n398), .B1(new_n414), .B2(new_n412), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n872), .B1(new_n889), .B2(new_n875), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n885), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n863), .B1(new_n880), .B2(new_n893), .ZN(new_n894));
  AND4_X1   g0694(.A1(new_n597), .A2(new_n621), .A3(new_n626), .A4(new_n628), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n672), .A2(new_n639), .A3(new_n895), .A4(new_n682), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n727), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n662), .A2(new_n365), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n366), .A2(new_n371), .A3(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n365), .B(new_n662), .C1(new_n370), .C2(new_n349), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n899), .A2(new_n903), .A3(new_n819), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT106), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n818), .B1(new_n896), .B2(new_n898), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT106), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(new_n903), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n894), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n633), .B1(KEYINPUT18), .B2(new_n416), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n869), .B1(new_n910), .B2(new_n428), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n881), .A2(new_n882), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n873), .B1(new_n912), .B2(new_n415), .ZN(new_n913));
  AOI22_X1  g0713(.A1(KEYINPUT37), .A2(new_n870), .B1(new_n913), .B2(new_n875), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n892), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n904), .B1(new_n880), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n909), .B1(KEYINPUT40), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n458), .A2(new_n899), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n862), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n918), .B2(new_n919), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n911), .A2(new_n914), .A3(new_n892), .ZN(new_n923));
  INV_X1    g0723(.A(new_n888), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n422), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT37), .B1(new_n883), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n876), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n927), .B2(new_n885), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n922), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT105), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n366), .B2(new_n662), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n349), .A2(KEYINPUT105), .A3(new_n365), .A4(new_n682), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n915), .A2(KEYINPUT39), .A3(new_n880), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n929), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n808), .A2(new_n662), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n651), .B2(new_n816), .ZN(new_n937));
  INV_X1    g0737(.A(new_n903), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n915), .A2(new_n880), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n939), .A2(new_n940), .B1(new_n884), .B2(new_n660), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n458), .B(new_n704), .C1(new_n705), .C2(KEYINPUT29), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n638), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n921), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n204), .B2(new_n734), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n921), .A2(new_n945), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n861), .B1(new_n947), .B2(new_n948), .ZN(G367));
  OR3_X1    g0749(.A1(new_n660), .A2(new_n585), .A3(new_n661), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT107), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n595), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n950), .A2(KEYINPUT107), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n950), .A2(KEYINPUT107), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(new_n596), .A3(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n558), .A2(new_n559), .B1(new_n486), .B2(new_n503), .ZN(new_n958));
  INV_X1    g0758(.A(new_n509), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n682), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n563), .A2(new_n683), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n662), .A2(new_n502), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n639), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n959), .A2(new_n662), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n961), .A2(KEYINPUT42), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT42), .B1(new_n961), .B2(new_n965), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n957), .B(new_n960), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT108), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n956), .B(KEYINPUT43), .Z(new_n970));
  OAI21_X1  g0770(.A(new_n960), .B1(new_n966), .B2(new_n967), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n968), .A2(KEYINPUT108), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n969), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n963), .A2(new_n964), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n681), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n974), .B(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n690), .B(KEYINPUT41), .Z(new_n978));
  NAND2_X1  g0778(.A1(new_n685), .A2(new_n686), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n979), .A2(KEYINPUT44), .A3(new_n975), .ZN(new_n980));
  AOI21_X1  g0780(.A(KEYINPUT44), .B1(new_n979), .B2(new_n975), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n979), .A2(new_n975), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT45), .B1(new_n687), .B2(new_n965), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n681), .B(new_n982), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n679), .A2(KEYINPUT109), .A3(new_n683), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT109), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n676), .B2(new_n684), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n685), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n670), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n987), .A2(new_n669), .A3(new_n989), .A4(new_n685), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n985), .A2(new_n984), .B1(new_n980), .B2(new_n981), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(new_n680), .A3(new_n677), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n986), .A2(new_n731), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n978), .B1(new_n996), .B2(new_n731), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n735), .A2(G1), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n977), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n757), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n208), .B2(new_n440), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n752), .A2(new_n233), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n737), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n776), .A2(new_n276), .B1(new_n777), .B2(new_n275), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n772), .A2(new_n251), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n248), .B1(new_n768), .B2(new_n835), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n274), .B2(new_n762), .C1(new_n836), .C2(new_n764), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n797), .A2(new_n783), .B1(new_n782), .B2(new_n832), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n789), .A2(G116), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT46), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n771), .B2(new_n762), .C1(new_n778), .C2(new_n764), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n772), .A2(new_n489), .ZN(new_n1013));
  INV_X1    g0813(.A(G317), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n336), .B1(new_n768), .B2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(G107), .C2(new_n775), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n516), .B2(new_n783), .C1(new_n759), .C2(new_n782), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n1008), .A2(new_n1009), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT47), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1003), .B1(new_n1019), .B2(new_n755), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n745), .B2(new_n956), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n999), .A2(new_n1021), .ZN(G387));
  INV_X1    g0822(.A(new_n998), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n991), .B2(new_n992), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT110), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n731), .A2(new_n993), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n694), .B1(new_n731), .B2(new_n993), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n336), .B1(new_n768), .B2(new_n781), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n759), .A2(new_n783), .B1(new_n782), .B2(new_n765), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT111), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n778), .A2(new_n762), .B1(new_n764), .B2(new_n1014), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT48), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(KEYINPUT48), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G294), .A2(new_n789), .B1(new_n775), .B2(G283), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT49), .Z(new_n1040));
  AOI211_X1 g0840(.A(new_n1029), .B(new_n1040), .C1(G116), .C2(new_n793), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n336), .B(new_n1013), .C1(G150), .C2(new_n769), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n789), .A2(G77), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n775), .A2(new_n589), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n274), .A2(new_n764), .B1(new_n762), .B2(new_n276), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n797), .A2(new_n782), .B1(new_n783), .B2(new_n283), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n755), .B1(new_n1041), .B2(new_n1048), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n230), .A2(new_n260), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1050), .A2(new_n751), .B1(new_n693), .B2(new_n747), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n280), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n274), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT50), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n461), .B1(new_n276), .B2(new_n251), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1054), .A2(new_n693), .A3(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1051), .A2(new_n1056), .B1(G107), .B2(new_n208), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n736), .B1(new_n1057), .B2(new_n1000), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1049), .B(new_n1058), .C1(new_n676), .C2(new_n745), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1025), .A2(new_n1028), .A3(new_n1059), .ZN(G393));
  NAND3_X1  g0860(.A1(new_n986), .A2(new_n998), .A3(new_n995), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n975), .A2(new_n744), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT112), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1000), .B1(new_n489), .B2(new_n208), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n751), .A2(new_n241), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n737), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n782), .A2(new_n1014), .B1(new_n764), .B2(new_n759), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT52), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n336), .B1(new_n768), .B2(new_n765), .C1(new_n494), .C2(new_n772), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n776), .A2(new_n599), .B1(new_n777), .B2(new_n771), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G294), .C2(new_n792), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1068), .B(new_n1071), .C1(new_n778), .C2(new_n783), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n782), .A2(new_n836), .B1(new_n764), .B2(new_n797), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT51), .Z(new_n1074));
  OAI221_X1 g0874(.A(new_n248), .B1(new_n772), .B2(new_n576), .C1(new_n768), .C2(new_n832), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n776), .A2(new_n251), .B1(new_n777), .B2(new_n276), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n1052), .C2(new_n792), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n274), .B2(new_n783), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1072), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1066), .B1(new_n1079), .B2(new_n755), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1063), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n996), .A2(new_n690), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n731), .A2(new_n993), .B1(new_n986), .B2(new_n995), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1061), .B(new_n1081), .C1(new_n1082), .C2(new_n1083), .ZN(G390));
  AOI22_X1  g0884(.A1(new_n871), .A2(new_n876), .B1(new_n429), .B2(new_n878), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n928), .B1(KEYINPUT38), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n934), .B1(new_n1086), .B2(KEYINPUT39), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n933), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n937), .B2(new_n938), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT113), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT113), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1088), .B(new_n1091), .C1(new_n937), .C2(new_n938), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1087), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n819), .B(new_n682), .C1(new_n701), .C2(new_n703), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n903), .B1(new_n1095), .B2(new_n936), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1086), .A2(new_n933), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1093), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n899), .A2(new_n903), .A3(new_n819), .A4(G330), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT114), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n906), .A2(KEYINPUT114), .A3(G330), .A4(new_n903), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(G330), .B(new_n819), .C1(new_n707), .C2(new_n729), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1106), .A2(new_n938), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1093), .A2(new_n1107), .A3(new_n1098), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n458), .A2(G330), .A3(new_n899), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n943), .A2(new_n638), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1106), .A2(new_n938), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1102), .A2(new_n1112), .A3(new_n1103), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n937), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n936), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n906), .A2(G330), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n938), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1107), .A2(new_n1116), .A3(new_n1094), .A4(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1111), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1109), .A2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n929), .A2(new_n934), .B1(new_n1089), .B2(KEYINPUT113), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1123), .A2(new_n1092), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1104), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1108), .B(new_n1120), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1122), .A2(new_n690), .A3(new_n1126), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1108), .B(new_n998), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT115), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT115), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1105), .A2(new_n1130), .A3(new_n998), .A4(new_n1108), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1087), .A2(new_n742), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n336), .B1(new_n769), .B2(G125), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n274), .B2(new_n772), .C1(new_n797), .C2(new_n776), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G128), .B2(new_n788), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n835), .B2(new_n783), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n795), .A2(G132), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT54), .B(G143), .Z(new_n1139));
  NAND2_X1  g0939(.A1(new_n792), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT53), .B1(new_n777), .B2(new_n836), .ZN(new_n1141));
  OR3_X1    g0941(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n836), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n788), .A2(G283), .B1(new_n792), .B2(G97), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n494), .B2(new_n783), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT116), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n336), .B1(new_n768), .B2(new_n516), .C1(new_n576), .C2(new_n777), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n776), .A2(new_n251), .B1(new_n772), .B2(new_n276), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(G116), .C2(new_n795), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1144), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n755), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n736), .B(new_n1153), .C1(new_n283), .C2(new_n823), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1133), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1127), .A2(new_n1132), .A3(new_n1155), .ZN(G378));
  XNOR2_X1  g0956(.A(new_n1111), .B(KEYINPUT120), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1126), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(G330), .B1(new_n916), .B2(KEYINPUT40), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n894), .A2(new_n905), .A3(new_n908), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n660), .B1(new_n288), .B2(new_n295), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n315), .B(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1159), .A2(new_n1160), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1163), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1162), .B(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n899), .A2(new_n819), .A3(new_n903), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT38), .B1(new_n877), .B2(new_n879), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1168), .B1(new_n923), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n862), .B1(new_n1170), .B2(new_n863), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1167), .B1(new_n1171), .B2(new_n909), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n942), .B1(new_n1165), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1164), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n935), .A2(new_n941), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(new_n909), .A3(new_n1167), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1158), .A2(new_n1178), .A3(KEYINPUT57), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1126), .A2(new_n1157), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n690), .C1(KEYINPUT57), .C2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT119), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1023), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n736), .B1(new_n274), .B2(new_n823), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n261), .B(new_n336), .C1(new_n768), .C2(new_n771), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1043), .B1(new_n275), .B2(new_n772), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(G68), .C2(new_n775), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n494), .B2(new_n764), .C1(new_n440), .C2(new_n762), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n489), .A2(new_n783), .B1(new_n782), .B2(new_n599), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT117), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G50), .B1(new_n245), .B2(new_n261), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n248), .B2(G41), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n783), .A2(new_n840), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n789), .A2(new_n1139), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n775), .A2(G150), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(G128), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1199), .B1(new_n762), .B2(new_n835), .C1(new_n1200), .C2(new_n764), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1196), .B(new_n1201), .C1(G125), .C2(new_n788), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n793), .A2(G159), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n769), .C2(G124), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  AND4_X1   g1008(.A1(new_n1192), .A2(new_n1193), .A3(new_n1195), .A4(new_n1208), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1184), .B1(new_n1152), .B2(new_n1209), .C1(new_n1167), .C2(new_n743), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT118), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1182), .B1(new_n1183), .B2(new_n1211), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1175), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n998), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT118), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1210), .B(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(KEYINPUT119), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1212), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1181), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1111), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n978), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(new_n1224), .A3(new_n1121), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n938), .A2(new_n742), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n783), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G132), .A2(new_n788), .B1(new_n1227), .B2(new_n1139), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n772), .A2(new_n275), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n248), .B1(new_n768), .B2(new_n1200), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(G159), .C2(new_n789), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1228), .B(new_n1231), .C1(new_n835), .C2(new_n764), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n762), .A2(new_n836), .B1(new_n776), .B2(new_n274), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT121), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G107), .A2(new_n792), .B1(new_n795), .B2(G283), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n248), .B(new_n1005), .C1(G303), .C2(new_n769), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n789), .A2(G97), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1235), .A2(new_n1044), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n599), .A2(new_n783), .B1(new_n782), .B2(new_n516), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1232), .A2(new_n1234), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1240), .A2(new_n755), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n736), .B(new_n1241), .C1(new_n276), .C2(new_n823), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1221), .A2(new_n998), .B1(new_n1226), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1225), .A2(new_n1243), .ZN(G381));
  NAND4_X1  g1044(.A1(new_n1025), .A2(new_n1028), .A3(new_n805), .A4(new_n1059), .ZN(new_n1245));
  OR4_X1    g1045(.A1(G384), .A2(G387), .A3(new_n1245), .A4(G390), .ZN(new_n1246));
  OR4_X1    g1046(.A1(G378), .A2(new_n1246), .A3(G375), .A4(G381), .ZN(G407));
  NAND2_X1  g1047(.A1(new_n661), .A2(G213), .ZN(new_n1248));
  OR3_X1    g1048(.A1(G375), .A2(G378), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(G213), .A3(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT122), .ZN(G409));
  INV_X1    g1051(.A(G390), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n999), .A2(new_n1021), .A3(G390), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT124), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G387), .B2(new_n1252), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1245), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1255), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1259), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1261), .A2(new_n1253), .A3(new_n1256), .A4(new_n1254), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1181), .A2(new_n1219), .A3(G378), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n694), .B1(new_n1109), .B2(new_n1121), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1265), .A2(new_n1126), .B1(new_n1133), .B2(new_n1154), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1158), .A2(new_n1224), .A3(new_n1178), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1215), .A2(new_n1210), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1266), .B(new_n1132), .C1(new_n1267), .C2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1264), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1248), .ZN(new_n1271));
  INV_X1    g1071(.A(G2897), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1248), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1222), .A2(KEYINPUT60), .A3(new_n1111), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n690), .A3(new_n1121), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1222), .B2(new_n1111), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1243), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(G384), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1276), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1223), .A2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1282), .A2(new_n690), .A3(new_n1121), .A4(new_n1274), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1283), .B2(new_n1243), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1273), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1283), .A2(G384), .A3(new_n1243), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1286), .B(new_n1287), .C1(new_n1272), .C2(new_n1248), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1271), .B2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1270), .A2(new_n1248), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT62), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1292), .A2(KEYINPUT62), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1263), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1280), .A2(new_n1284), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1270), .A2(new_n1248), .A3(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT61), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1248), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1264), .B2(new_n1269), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1303), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1302), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1292), .A2(new_n1298), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1297), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1263), .B1(new_n1305), .B2(new_n1299), .ZN(new_n1311));
  AND4_X1   g1111(.A1(new_n1297), .A2(new_n1290), .A3(new_n1309), .A4(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1296), .B1(new_n1310), .B2(new_n1312), .ZN(G405));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1291), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT127), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1291), .A2(new_n1314), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1301), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1316), .A2(new_n1263), .A3(new_n1318), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1291), .A2(new_n1314), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(G375), .A2(new_n1132), .A3(new_n1266), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1264), .B2(new_n1324), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1322), .B(new_n1325), .ZN(G402));
endmodule


