//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1030, new_n1031;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G211gat), .B(G218gat), .Z(new_n210));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n209), .B(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(G148gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G141gat), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G148gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT72), .B(KEYINPUT2), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n214), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT2), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT74), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g025(.A(KEYINPUT74), .B(KEYINPUT2), .C1(new_n222), .C2(new_n223), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n226), .A2(new_n214), .A3(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT73), .B(G141gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n216), .B1(new_n229), .B2(new_n215), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n221), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n213), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G228gat), .A2(G233gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n221), .ZN(new_n238));
  INV_X1    g037(.A(new_n230), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n226), .A2(new_n214), .A3(new_n227), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT75), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n238), .B(KEYINPUT75), .C1(new_n239), .C2(new_n240), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n212), .B(new_n208), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT29), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n243), .B(new_n244), .C1(new_n246), .C2(KEYINPUT3), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n237), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT80), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n208), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(new_n210), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(KEYINPUT29), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n209), .A2(KEYINPUT80), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n210), .A3(new_n250), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n231), .B1(new_n255), .B2(new_n232), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n236), .B1(new_n256), .B2(new_n235), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n248), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G22gat), .ZN(new_n259));
  INV_X1    g058(.A(G22gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n248), .A2(new_n260), .A3(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n259), .A2(KEYINPUT81), .ZN(new_n263));
  XOR2_X1   g062(.A(G78gat), .B(G106gat), .Z(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT79), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT31), .B(G50gat), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n265), .B(new_n266), .Z(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n262), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n268), .B1(new_n259), .B2(KEYINPUT81), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(new_n259), .A3(new_n261), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G15gat), .B(G43gat), .Z(new_n273));
  XNOR2_X1  g072(.A(G71gat), .B(G99gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G227gat), .ZN(new_n276));
  INV_X1    g075(.A(G233gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G113gat), .ZN(new_n280));
  INV_X1    g079(.A(G120gat), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n280), .B2(new_n281), .ZN(new_n283));
  XOR2_X1   g082(.A(G127gat), .B(G134gat), .Z(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT24), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT24), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT66), .B(G190gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT65), .B(G183gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT23), .ZN(new_n295));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(G169gat), .B2(G176gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n293), .A2(new_n300), .A3(KEYINPUT25), .ZN(new_n301));
  NOR2_X1   g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT64), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n299), .B1(new_n306), .B2(new_n290), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n301), .B1(new_n307), .B2(KEYINPUT25), .ZN(new_n308));
  INV_X1    g107(.A(G169gat), .ZN(new_n309));
  INV_X1    g108(.A(G176gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT26), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n296), .B1(new_n311), .B2(KEYINPUT26), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n286), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n316));
  OR2_X1    g115(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT27), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G183gat), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n317), .B(new_n318), .C1(new_n320), .C2(KEYINPUT67), .ZN(new_n321));
  NAND2_X1  g120(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(KEYINPUT67), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT27), .B1(KEYINPUT65), .B2(G183gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n316), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n317), .A2(KEYINPUT28), .A3(new_n318), .ZN(new_n327));
  INV_X1    g126(.A(G183gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT27), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n315), .B1(new_n326), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n308), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n296), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(new_n294), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n338), .A2(new_n312), .B1(G183gat), .B2(G190gat), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n328), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n291), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n324), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(KEYINPUT67), .B2(new_n322), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT28), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n339), .B(new_n334), .C1(new_n344), .C2(new_n331), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n285), .B1(new_n335), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n339), .B1(new_n344), .B2(new_n331), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT25), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n290), .A2(new_n305), .A3(new_n304), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n299), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n348), .A2(KEYINPUT68), .B1(new_n351), .B2(new_n301), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n283), .A2(new_n284), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n283), .A2(new_n284), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n355), .A3(new_n345), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n279), .B1(new_n347), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n275), .B1(new_n357), .B2(KEYINPUT33), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT32), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n347), .A2(new_n356), .ZN(new_n362));
  AOI221_X4 g161(.A(new_n359), .B1(KEYINPUT33), .B2(new_n275), .C1(new_n362), .C2(new_n278), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n356), .A3(new_n279), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT69), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT34), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n361), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n366), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n362), .A2(new_n278), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT33), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n372), .A3(new_n275), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n360), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n368), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI22_X1  g174(.A1(new_n367), .A2(new_n375), .B1(new_n365), .B2(new_n364), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n366), .B1(new_n361), .B2(new_n363), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n373), .A2(new_n374), .A3(new_n368), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n364), .A2(new_n365), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n272), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n308), .A2(new_n348), .ZN(new_n382));
  NAND2_X1  g181(.A1(G226gat), .A2(G233gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n348), .A2(KEYINPUT68), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n345), .A3(new_n308), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n384), .B1(new_n387), .B2(new_n234), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n385), .B1(new_n388), .B2(KEYINPUT71), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT71), .ZN(new_n390));
  AOI211_X1 g189(.A(new_n390), .B(new_n384), .C1(new_n387), .C2(new_n234), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n245), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n382), .A2(new_n234), .A3(new_n383), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n387), .B2(new_n383), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n213), .ZN(new_n395));
  XNOR2_X1  g194(.A(G8gat), .B(G36gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(G64gat), .ZN(new_n397));
  INV_X1    g196(.A(G92gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n392), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT30), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n392), .A2(KEYINPUT30), .A3(new_n395), .A4(new_n399), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n392), .A2(new_n395), .ZN(new_n404));
  INV_X1    g203(.A(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n243), .A2(new_n244), .A3(new_n285), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n231), .A2(new_n355), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n408), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n243), .A2(KEYINPUT3), .A3(new_n244), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n285), .A3(new_n233), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(new_n241), .B2(new_n285), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n413), .B1(new_n241), .B2(new_n285), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n355), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n418), .A2(new_n420), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n410), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n413), .A2(KEYINPUT5), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n426), .A2(new_n416), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G1gat), .B(G29gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT0), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(G57gat), .ZN(new_n433));
  INV_X1    g232(.A(G85gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n423), .A2(new_n429), .A3(new_n435), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n437), .A2(KEYINPUT78), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n430), .A2(KEYINPUT6), .A3(new_n436), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT78), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n407), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n202), .B1(new_n381), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n402), .A2(new_n403), .A3(new_n406), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n270), .B(new_n262), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n379), .B1(new_n377), .B2(new_n378), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n448), .B(new_n449), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n443), .A2(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n202), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n447), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n453), .ZN(new_n457));
  INV_X1    g256(.A(new_n404), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n399), .B1(new_n458), .B2(KEYINPUT38), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n392), .A2(new_n460), .A3(new_n395), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT38), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n392), .B2(new_n395), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n213), .B1(new_n389), .B2(new_n391), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n460), .B1(new_n394), .B2(new_n245), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n399), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT38), .B1(new_n467), .B2(new_n461), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n457), .B(new_n459), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n426), .A2(new_n416), .A3(new_n427), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT82), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n413), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n472), .B1(new_n471), .B2(new_n413), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n475), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n411), .A2(new_n413), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(new_n470), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n473), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(new_n480), .A3(new_n435), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT40), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n476), .A2(new_n480), .A3(KEYINPUT40), .A4(new_n435), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n407), .A3(new_n437), .A4(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n469), .A2(new_n485), .A3(new_n449), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n450), .B2(new_n451), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n376), .A2(KEYINPUT36), .A3(new_n380), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n488), .B(new_n489), .C1(new_n446), .C2(new_n449), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n456), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT14), .ZN(new_n495));
  INV_X1    g294(.A(G29gat), .ZN(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G50gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(G43gat), .ZN(new_n502));
  INV_X1    g301(.A(G43gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G50gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g304(.A1(G29gat), .A2(G36gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n500), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n501), .B2(G43gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n503), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n511));
  AND2_X1   g310(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n510), .B(new_n511), .C1(new_n514), .C2(G50gat), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n507), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT85), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(KEYINPUT85), .A3(new_n497), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n499), .A2(KEYINPUT84), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT84), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n522), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n518), .A2(new_n520), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n505), .B1(new_n524), .B2(new_n506), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n494), .B1(new_n516), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n528));
  AOI21_X1  g327(.A(G50gat), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n511), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n508), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT15), .B1(new_n501), .B2(G43gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n503), .A2(G50gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n506), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n496), .A2(new_n497), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n535), .A2(KEYINPUT14), .B1(new_n519), .B2(new_n497), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n506), .ZN(new_n539));
  NOR4_X1   g338(.A1(new_n517), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT85), .B1(new_n519), .B2(new_n497), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n521), .A2(new_n523), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n538), .B(KEYINPUT17), .C1(new_n544), .C2(new_n505), .ZN(new_n545));
  INV_X1    g344(.A(G8gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n260), .A2(G15gat), .ZN(new_n547));
  INV_X1    g346(.A(G15gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G22gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n549), .A3(KEYINPUT88), .ZN(new_n550));
  INV_X1    g349(.A(G1gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(KEYINPUT88), .A3(G1gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT16), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AND4_X1   g355(.A1(new_n546), .A2(new_n552), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n550), .A2(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n546), .B1(new_n558), .B2(new_n554), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n526), .A2(new_n545), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT89), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n557), .B2(new_n559), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n538), .B1(new_n544), .B2(new_n505), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G8gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n558), .A2(new_n546), .A3(new_n554), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(KEYINPUT89), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n563), .A2(KEYINPUT90), .A3(new_n568), .A4(new_n564), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n493), .B(new_n561), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT91), .B1(new_n573), .B2(KEYINPUT18), .ZN(new_n574));
  XNOR2_X1  g373(.A(G169gat), .B(G197gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT12), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n571), .A2(new_n572), .ZN(new_n582));
  INV_X1    g381(.A(new_n561), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT18), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n493), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n564), .B1(new_n563), .B2(new_n568), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n571), .B2(new_n572), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n492), .B(KEYINPUT13), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n561), .B1(new_n571), .B2(new_n572), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT18), .B1(new_n592), .B2(new_n492), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n574), .B(new_n581), .C1(new_n591), .C2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n587), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n582), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n596), .A2(new_n589), .B1(new_n592), .B2(new_n585), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n492), .A3(new_n583), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n584), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n597), .B(new_n599), .C1(KEYINPUT91), .C2(new_n580), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n491), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n603));
  XOR2_X1   g402(.A(G99gat), .B(G106gat), .Z(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G85gat), .A2(G92gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT7), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT7), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(G85gat), .A3(G92gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n612), .B1(new_n434), .B2(new_n398), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n611), .B1(new_n610), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n605), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n613), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT95), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n610), .A2(new_n613), .A3(new_n611), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n604), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n603), .B1(new_n621), .B2(new_n564), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n620), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n526), .A2(new_n545), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT96), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT98), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n630), .A3(new_n627), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(new_n625), .B2(new_n627), .ZN(new_n637));
  INV_X1    g436(.A(new_n627), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n622), .A2(KEYINPUT97), .A3(new_n624), .A4(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n635), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n632), .A2(new_n640), .A3(KEYINPUT99), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT99), .B1(new_n632), .B2(new_n640), .ZN(new_n642));
  INV_X1    g441(.A(new_n635), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n637), .A2(new_n639), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n628), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n641), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(G57gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(G64gat), .ZN(new_n648));
  INV_X1    g447(.A(G64gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(G57gat), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n648), .B1(KEYINPUT92), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT92), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n649), .B2(G57gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G71gat), .A2(G78gat), .ZN(new_n655));
  OR2_X1    g454(.A1(G71gat), .A2(G78gat), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT9), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT9), .B1(new_n650), .B2(new_n648), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n656), .A2(new_n655), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n654), .A2(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n563), .A2(new_n568), .B1(KEYINPUT21), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(new_n328), .ZN(new_n663));
  XNOR2_X1  g462(.A(G127gat), .B(G155gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT20), .ZN(new_n665));
  NAND2_X1  g464(.A1(G231gat), .A2(G233gat), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT93), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n665), .B(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n663), .A2(new_n668), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n661), .A2(KEYINPUT21), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G211gat), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n669), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n674), .B1(new_n669), .B2(new_n670), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(G230gat), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n277), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n616), .A2(new_n620), .A3(new_n661), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n661), .B1(new_n616), .B2(new_n620), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n681), .A2(new_n682), .A3(KEYINPUT10), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n616), .A2(new_n620), .A3(new_n661), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT10), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n680), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n661), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n623), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n680), .B1(new_n689), .B2(new_n684), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(G120gat), .B(G148gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G176gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G204gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n687), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n689), .A2(new_n685), .A3(new_n684), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n681), .A2(KEYINPUT10), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n679), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n694), .B1(new_n699), .B2(new_n690), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n696), .A2(new_n700), .A3(KEYINPUT100), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n702), .B(new_n694), .C1(new_n699), .C2(new_n690), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n646), .A2(new_n677), .A3(new_n704), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n705), .A2(KEYINPUT101), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(KEYINPUT101), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n602), .A2(KEYINPUT102), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT102), .B1(new_n602), .B2(new_n708), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n445), .A2(new_n440), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(new_n551), .ZN(G1324gat));
  OAI21_X1  g514(.A(new_n407), .B1(new_n709), .B2(new_n710), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT16), .B(G8gat), .Z(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT103), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n716), .A2(G8gat), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n722));
  OAI211_X1 g521(.A(KEYINPUT103), .B(new_n722), .C1(new_n716), .C2(new_n718), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(G1325gat));
  NAND2_X1  g523(.A1(new_n488), .A2(new_n489), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G15gat), .B1(new_n711), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n450), .A2(new_n451), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n548), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n711), .B2(new_n730), .ZN(G1326gat));
  OAI21_X1  g530(.A(new_n272), .B1(new_n709), .B2(new_n710), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT43), .B(G22gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1327gat));
  NOR2_X1   g533(.A1(new_n646), .A2(new_n677), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n704), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n602), .A2(new_n496), .A3(new_n712), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT45), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n447), .A2(new_n455), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT105), .B1(new_n486), .B2(new_n490), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n469), .A2(new_n485), .A3(new_n449), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n272), .B1(new_n712), .B2(new_n407), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n726), .A2(new_n744), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n742), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n741), .B1(new_n748), .B2(new_n646), .ZN(new_n749));
  INV_X1    g548(.A(new_n646), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n491), .A2(KEYINPUT44), .A3(new_n750), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n704), .B(KEYINPUT104), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n594), .A2(new_n600), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n753), .A2(new_n754), .A3(new_n677), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n752), .A2(new_n712), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT106), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G29gat), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n756), .A2(KEYINPUT106), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n740), .B1(new_n758), .B2(new_n759), .ZN(G1328gat));
  NAND4_X1  g559(.A1(new_n602), .A2(new_n497), .A3(new_n407), .A4(new_n738), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(KEYINPUT107), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n762), .A2(KEYINPUT107), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n752), .A2(new_n407), .A3(new_n755), .ZN(new_n766));
  OAI221_X1 g565(.A(new_n765), .B1(new_n763), .B2(new_n761), .C1(new_n766), .C2(new_n497), .ZN(G1329gat));
  NAND4_X1  g566(.A1(new_n749), .A2(new_n751), .A3(new_n725), .A4(new_n755), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n513), .B2(new_n512), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n602), .A2(new_n729), .A3(new_n514), .A4(new_n738), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT47), .Z(G1330gat));
  NAND4_X1  g571(.A1(new_n602), .A2(new_n501), .A3(new_n272), .A4(new_n738), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n749), .A2(new_n751), .A3(new_n272), .A4(new_n755), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G50gat), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n774), .A2(new_n775), .ZN(new_n778));
  OAI211_X1 g577(.A(KEYINPUT48), .B(new_n773), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n774), .A2(G50gat), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n773), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(KEYINPUT48), .B2(new_n781), .ZN(G1331gat));
  NAND2_X1  g581(.A1(new_n743), .A2(new_n747), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n601), .B1(new_n783), .B2(new_n456), .ZN(new_n784));
  INV_X1    g583(.A(new_n677), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n750), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n786), .A3(new_n753), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n713), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(new_n647), .ZN(G1332gat));
  NOR2_X1   g588(.A1(new_n787), .A2(new_n448), .ZN(new_n790));
  NOR2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  AND2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n790), .B2(new_n791), .ZN(G1333gat));
  INV_X1    g593(.A(new_n787), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(G71gat), .A3(new_n725), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n728), .B(KEYINPUT109), .Z(new_n797));
  NOR2_X1   g596(.A1(new_n787), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n798), .B2(G71gat), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g599(.A1(new_n795), .A2(new_n272), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g601(.A1(new_n704), .A2(G85gat), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n783), .A2(new_n456), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(new_n754), .A3(new_n735), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n784), .A2(KEYINPUT51), .A3(new_n735), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(KEYINPUT110), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(KEYINPUT110), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n712), .B(new_n803), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n677), .A2(new_n601), .A3(new_n704), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n752), .A2(new_n712), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n434), .B2(new_n814), .ZN(G1336gat));
  NAND3_X1  g614(.A1(new_n752), .A2(new_n407), .A3(new_n813), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G92gat), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n809), .A2(new_n398), .A3(new_n407), .A4(new_n753), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT52), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(G1337gat));
  INV_X1    g622(.A(G99gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n752), .A2(new_n725), .A3(new_n813), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n825), .B2(KEYINPUT111), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n826), .B1(KEYINPUT111), .B2(new_n825), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n728), .A2(G99gat), .A3(new_n704), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n810), .B2(new_n811), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(G1338gat));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n449), .A2(G106gat), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n809), .A2(new_n831), .A3(new_n753), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT51), .B1(new_n784), .B2(new_n735), .ZN(new_n834));
  NOR4_X1   g633(.A1(new_n748), .A2(new_n806), .A3(new_n601), .A4(new_n736), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n753), .B(new_n832), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT112), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n749), .A2(new_n751), .A3(new_n272), .A4(new_n813), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G106gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n833), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT53), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT53), .B1(new_n838), .B2(G106gat), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n836), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n836), .A2(new_n843), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n841), .A2(new_n846), .ZN(G1339gat));
  NOR2_X1   g646(.A1(new_n705), .A2(new_n601), .ZN(new_n848));
  INV_X1    g647(.A(new_n696), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n697), .A2(new_n698), .A3(new_n679), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n687), .A2(KEYINPUT54), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n695), .B1(new_n699), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n849), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n851), .A2(new_n853), .A3(KEYINPUT55), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT114), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n851), .A2(new_n853), .A3(new_n859), .A4(KEYINPUT55), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n596), .A2(new_n589), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n599), .A2(new_n862), .A3(new_n586), .A4(new_n580), .ZN(new_n863));
  INV_X1    g662(.A(new_n579), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n592), .A2(new_n492), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n587), .B(new_n589), .C1(new_n571), .C2(new_n572), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n646), .A2(new_n861), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n863), .A2(new_n703), .A3(new_n701), .A4(new_n867), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT115), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n737), .A2(new_n872), .A3(new_n867), .A4(new_n863), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n871), .B(new_n873), .C1(new_n754), .C2(new_n861), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n869), .B1(new_n874), .B2(new_n646), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n677), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n856), .A2(new_n860), .A3(new_n858), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n878), .A2(new_n601), .B1(KEYINPUT115), .B2(new_n870), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n750), .B1(new_n879), .B2(new_n873), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT116), .B1(new_n880), .B2(new_n869), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n848), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(new_n713), .A3(new_n452), .ZN(new_n883));
  AOI21_X1  g682(.A(G113gat), .B1(new_n883), .B2(new_n601), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n713), .A2(new_n407), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR4_X1   g685(.A1(new_n882), .A2(new_n272), .A3(new_n728), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n754), .A2(new_n280), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(G1340gat));
  AOI21_X1  g688(.A(G120gat), .B1(new_n883), .B2(new_n737), .ZN(new_n890));
  INV_X1    g689(.A(new_n753), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n281), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n887), .B2(new_n892), .ZN(G1341gat));
  INV_X1    g692(.A(G127gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n883), .A2(new_n894), .A3(new_n677), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n887), .A2(new_n677), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n894), .ZN(G1342gat));
  AND2_X1   g696(.A1(new_n887), .A2(new_n750), .ZN(new_n898));
  INV_X1    g697(.A(G134gat), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n883), .A2(new_n899), .A3(new_n750), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(KEYINPUT56), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(KEYINPUT56), .B2(new_n901), .ZN(G1343gat));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n882), .B2(new_n449), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT117), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n907), .B(new_n904), .C1(new_n882), .C2(new_n449), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n449), .A2(new_n904), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT118), .B(new_n870), .C1(new_n754), .C2(new_n861), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n878), .A2(new_n601), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT118), .B1(new_n912), .B2(new_n870), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n646), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n869), .B1(new_n914), .B2(KEYINPUT119), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n916), .B(new_n646), .C1(new_n911), .C2(new_n913), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n677), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n909), .B1(new_n918), .B2(new_n848), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n906), .A2(new_n908), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n886), .A2(new_n725), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n601), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n229), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n726), .A2(new_n272), .ZN(new_n924));
  NOR4_X1   g723(.A1(new_n882), .A2(new_n713), .A3(new_n407), .A4(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n217), .A3(new_n601), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT58), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n928), .B1(new_n926), .B2(KEYINPUT120), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n923), .B(new_n926), .C1(KEYINPUT120), .C2(new_n928), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1344gat));
  OAI21_X1  g731(.A(KEYINPUT57), .B1(new_n882), .B2(new_n449), .ZN(new_n933));
  INV_X1    g732(.A(new_n869), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n677), .B1(new_n914), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n601), .B1(new_n706), .B2(new_n707), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n904), .B(new_n272), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(new_n737), .A3(new_n921), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT59), .B1(new_n939), .B2(new_n215), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n215), .A2(KEYINPUT59), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n920), .A2(new_n921), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n704), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n925), .A2(new_n215), .A3(new_n737), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1345gat));
  OAI21_X1  g745(.A(G155gat), .B1(new_n942), .B2(new_n785), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n925), .A2(new_n222), .A3(new_n677), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1346gat));
  NAND3_X1  g748(.A1(new_n920), .A2(new_n750), .A3(new_n921), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G162gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n925), .A2(new_n223), .A3(new_n750), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT121), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT121), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n955), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1347gat));
  INV_X1    g756(.A(new_n848), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n874), .A2(new_n646), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n876), .A3(new_n934), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(new_n785), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n875), .A2(new_n876), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(new_n964), .A3(new_n713), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT122), .B1(new_n882), .B2(new_n712), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n381), .A2(new_n407), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(G169gat), .B1(new_n970), .B2(new_n601), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n882), .A2(new_n272), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n713), .A2(new_n407), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n797), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n972), .A2(KEYINPUT123), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT123), .B1(new_n972), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n754), .A2(new_n309), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n971), .B1(new_n977), .B2(new_n978), .ZN(G1348gat));
  NAND3_X1  g778(.A1(new_n970), .A2(new_n310), .A3(new_n737), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n975), .A2(new_n976), .A3(new_n891), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n981), .B2(new_n310), .ZN(G1349gat));
  NAND4_X1  g781(.A1(new_n970), .A2(new_n320), .A3(new_n329), .A4(new_n677), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT60), .ZN(new_n984));
  INV_X1    g783(.A(new_n292), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n975), .A2(new_n976), .A3(new_n785), .ZN(new_n986));
  OAI211_X1 g785(.A(new_n983), .B(new_n984), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n986), .A2(new_n985), .ZN(new_n988));
  NOR4_X1   g787(.A1(new_n968), .A2(new_n330), .A3(new_n785), .A4(new_n969), .ZN(new_n989));
  OAI21_X1  g788(.A(KEYINPUT60), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n987), .A2(new_n990), .ZN(G1350gat));
  INV_X1    g790(.A(G190gat), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n992), .B1(new_n977), .B2(new_n750), .ZN(new_n993));
  OR2_X1    g792(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n994));
  NAND2_X1  g793(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n970), .A2(new_n317), .A3(new_n318), .A4(new_n750), .ZN(new_n997));
  OAI211_X1 g796(.A(new_n996), .B(new_n997), .C1(new_n993), .C2(new_n994), .ZN(G1351gat));
  NAND3_X1  g797(.A1(new_n726), .A2(new_n407), .A3(new_n272), .ZN(new_n999));
  XOR2_X1   g798(.A(new_n999), .B(KEYINPUT125), .Z(new_n1000));
  AND2_X1   g799(.A1(new_n967), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g800(.A(G197gat), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n1001), .A2(new_n1002), .A3(new_n601), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n973), .A2(new_n725), .ZN(new_n1004));
  AND2_X1   g803(.A1(new_n938), .A2(new_n1004), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n1005), .A2(new_n601), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1003), .B1(new_n1006), .B2(new_n1002), .ZN(G1352gat));
  INV_X1    g806(.A(KEYINPUT62), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n704), .A2(G204gat), .ZN(new_n1009));
  NAND4_X1  g808(.A1(new_n967), .A2(new_n1008), .A3(new_n1000), .A4(new_n1009), .ZN(new_n1010));
  NAND4_X1  g809(.A1(new_n933), .A2(new_n753), .A3(new_n937), .A4(new_n1004), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1011), .A2(G204gat), .ZN(new_n1012));
  AND2_X1   g811(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n964), .B1(new_n963), .B2(new_n713), .ZN(new_n1014));
  NOR3_X1   g813(.A1(new_n882), .A2(KEYINPUT122), .A3(new_n712), .ZN(new_n1015));
  OAI211_X1 g814(.A(new_n1000), .B(new_n1009), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1017));
  AND3_X1   g816(.A1(new_n1016), .A2(new_n1017), .A3(KEYINPUT62), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n1017), .B1(new_n1016), .B2(KEYINPUT62), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1013), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1020), .A2(KEYINPUT127), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT127), .ZN(new_n1022));
  OAI211_X1 g821(.A(new_n1013), .B(new_n1022), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1021), .A2(new_n1023), .ZN(G1353gat));
  NAND3_X1  g823(.A1(new_n1001), .A2(new_n205), .A3(new_n677), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1005), .A2(new_n677), .ZN(new_n1026));
  AND3_X1   g825(.A1(new_n1026), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1027));
  AOI21_X1  g826(.A(KEYINPUT63), .B1(new_n1026), .B2(G211gat), .ZN(new_n1028));
  OAI21_X1  g827(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(G1354gat));
  NAND3_X1  g828(.A1(new_n1001), .A2(new_n206), .A3(new_n750), .ZN(new_n1030));
  AND2_X1   g829(.A1(new_n1005), .A2(new_n750), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n1030), .B1(new_n1031), .B2(new_n206), .ZN(G1355gat));
endmodule


