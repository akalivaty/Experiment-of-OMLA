//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR3_X1   g0010(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT64), .Z(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT67), .B(G238), .ZN(new_n215));
  AOI22_X1  g0015(.A1(new_n215), .A2(G68), .B1(G77), .B2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n206), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G116), .ZN(new_n221));
  INV_X1    g0021(.A(G270), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n205), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g0025(.A1(G50), .A2(G226), .ZN(new_n226));
  NOR4_X1   g0026(.A1(new_n220), .A2(new_n223), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G87), .A2(G250), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n227), .A2(new_n228), .B1(G1), .B2(G20), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT1), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n214), .B(new_n230), .C1(new_n234), .C2(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G226), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n222), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT69), .B(G264), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n242), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT70), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT21), .ZN(new_n256));
  INV_X1    g0056(.A(G45), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT5), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  OAI211_X1 g0066(.A(G1), .B(G13), .C1(new_n266), .C2(new_n259), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n265), .B1(new_n222), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n266), .A2(KEYINPUT83), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT83), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(new_n277), .B2(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G264), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT90), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n271), .B1(new_n274), .B2(new_n276), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT90), .ZN(new_n283));
  NOR4_X1   g0083(.A1(new_n282), .A2(new_n283), .A3(new_n273), .A4(new_n279), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT83), .B(G33), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n286), .B(new_n272), .C1(new_n287), .C2(new_n271), .ZN(new_n288));
  INV_X1    g0088(.A(G303), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n272), .A2(new_n290), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n288), .A2(new_n224), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT91), .B1(new_n285), .B2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n272), .B(new_n280), .C1(new_n287), .C2(new_n271), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n283), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n297), .A2(KEYINPUT90), .A3(new_n272), .A4(new_n280), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT91), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n299), .A2(new_n292), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n270), .B1(new_n294), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT92), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n285), .A2(new_n293), .A3(KEYINPUT91), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n300), .B1(new_n299), .B2(new_n292), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT92), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(new_n270), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n269), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n232), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n209), .A2(G20), .ZN(new_n312));
  INV_X1    g0112(.A(G13), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI211_X1 g0114(.A(new_n311), .B(new_n314), .C1(new_n209), .C2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G116), .ZN(new_n316));
  INV_X1    g0116(.A(new_n314), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G283), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n231), .B(new_n318), .C1(G33), .C2(new_n205), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n319), .B(new_n311), .C1(new_n210), .C2(G116), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT20), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n320), .A2(new_n321), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n316), .B1(G116), .B2(new_n317), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G169), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n256), .B1(new_n309), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n309), .A2(G179), .A3(new_n324), .ZN(new_n327));
  INV_X1    g0127(.A(new_n269), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n307), .B1(new_n306), .B2(new_n270), .ZN(new_n329));
  AOI211_X1 g0129(.A(KEYINPUT92), .B(new_n267), .C1(new_n304), .C2(new_n305), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n325), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(KEYINPUT21), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n326), .A2(new_n327), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT72), .ZN(new_n336));
  AOI21_X1  g0136(.A(G1), .B1(new_n259), .B2(new_n257), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT71), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n264), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n267), .B1(new_n337), .B2(new_n338), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n341), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(KEYINPUT72), .A3(new_n339), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n270), .A2(new_n337), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G238), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n218), .A2(G1698), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n291), .B(new_n351), .C1(G226), .C2(G1698), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n266), .B2(new_n205), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT81), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n352), .B(KEYINPUT81), .C1(new_n266), .C2(new_n205), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n270), .A3(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n349), .A2(new_n350), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n350), .B1(new_n349), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g0159(.A(G200), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n349), .A2(new_n357), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT13), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n349), .A2(new_n350), .A3(new_n357), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(G190), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(G20), .A2(G33), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G50), .ZN(new_n366));
  AND2_X1   g0166(.A1(KEYINPUT65), .A2(G20), .ZN(new_n367));
  NOR2_X1   g0167(.A1(KEYINPUT65), .A2(G20), .ZN(new_n368));
  OAI21_X1  g0168(.A(G33), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G77), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n366), .B1(new_n210), .B2(G68), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n311), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n372), .A2(KEYINPUT11), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(KEYINPUT11), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n317), .A2(KEYINPUT12), .A3(G68), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT12), .ZN(new_n377));
  INV_X1    g0177(.A(G68), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n377), .B1(new_n314), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n312), .A2(new_n232), .A3(new_n310), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n376), .A2(new_n379), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n360), .A2(new_n364), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(G169), .B1(new_n358), .B2(new_n359), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT14), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT14), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n386), .B(G169), .C1(new_n358), .C2(new_n359), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n362), .A2(G179), .A3(new_n363), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n382), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n383), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n391), .A2(KEYINPUT82), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n390), .ZN(new_n393));
  INV_X1    g0193(.A(new_n383), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(KEYINPUT82), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G244), .ZN(new_n396));
  INV_X1    g0196(.A(new_n346), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n345), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT75), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n291), .A2(G1698), .A3(new_n215), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n206), .B2(new_n291), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n272), .A2(new_n290), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n403), .A2(new_n218), .A3(G1698), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n270), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n398), .A2(new_n399), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n400), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n407), .A2(G179), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT8), .B(G58), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT76), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n365), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT15), .B(G87), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n413), .A2(KEYINPUT77), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(KEYINPUT77), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n411), .B1(new_n370), .B2(new_n231), .C1(new_n416), .C2(new_n369), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n311), .B1(new_n370), .B2(new_n314), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n380), .A2(new_n370), .ZN(new_n419));
  XOR2_X1   g0219(.A(new_n419), .B(KEYINPUT78), .Z(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G169), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n407), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n408), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n392), .A2(new_n395), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT79), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n317), .A2(G50), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n380), .A2(new_n202), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n365), .A2(G150), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT8), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G58), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(G58), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(KEYINPUT73), .ZN(new_n434));
  OR3_X1    g0234(.A1(new_n217), .A2(KEYINPUT73), .A3(KEYINPUT8), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(KEYINPUT74), .B(new_n430), .C1(new_n436), .C2(new_n369), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n203), .A2(G20), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT74), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n369), .B1(new_n434), .B2(new_n435), .ZN(new_n440));
  INV_X1    g0240(.A(new_n430), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n437), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  AOI211_X1 g0243(.A(new_n428), .B(new_n429), .C1(new_n443), .C2(new_n311), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n427), .B1(new_n444), .B2(KEYINPUT9), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n311), .ZN(new_n446));
  INV_X1    g0246(.A(new_n428), .ZN(new_n447));
  INV_X1    g0247(.A(new_n429), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT9), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(KEYINPUT79), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT80), .B1(new_n449), .B2(new_n450), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT80), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n444), .A2(new_n454), .A3(KEYINPUT9), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n346), .A2(G226), .ZN(new_n457));
  INV_X1    g0257(.A(G223), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G1698), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(G222), .B2(G1698), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n267), .B1(new_n291), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(G77), .B2(new_n291), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n345), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G200), .ZN(new_n464));
  INV_X1    g0264(.A(G190), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(new_n463), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n452), .A2(new_n456), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT10), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n445), .B2(new_n451), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT10), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n456), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n463), .A2(G179), .ZN(new_n474));
  AOI211_X1 g0274(.A(new_n474), .B(new_n444), .C1(new_n423), .C2(new_n463), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n422), .B1(new_n407), .B2(G200), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n465), .B2(new_n407), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT16), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n274), .A2(new_n276), .A3(new_n271), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n290), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT7), .B1(new_n403), .B2(new_n210), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n378), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(G58), .A2(G68), .ZN(new_n487));
  OAI21_X1  g0287(.A(G20), .B1(new_n487), .B2(new_n201), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n365), .A2(G159), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT84), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(KEYINPUT84), .A3(new_n489), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n480), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT85), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT7), .B1(new_n278), .B2(G20), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT7), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n498), .B(new_n231), .C1(new_n282), .C2(new_n273), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(G68), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n492), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n490), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(KEYINPUT16), .A3(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(KEYINPUT85), .B(new_n480), .C1(new_n486), .C2(new_n493), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n496), .A2(new_n311), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n342), .A2(new_n344), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n458), .A2(new_n286), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n278), .B(new_n507), .C1(G226), .C2(new_n286), .ZN(new_n508));
  INV_X1    g0308(.A(G87), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n266), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n267), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n337), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G232), .A3(new_n267), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT86), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n506), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G190), .ZN(new_n518));
  INV_X1    g0318(.A(new_n436), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n380), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n314), .B2(new_n519), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n508), .A2(new_n511), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n270), .ZN(new_n523));
  INV_X1    g0323(.A(new_n516), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n345), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G200), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n505), .A2(new_n518), .A3(new_n521), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n521), .ZN(new_n530));
  INV_X1    g0330(.A(new_n504), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n367), .A2(new_n368), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n481), .B2(new_n290), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n484), .B1(new_n533), .B2(KEYINPUT7), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n502), .B1(new_n534), .B2(new_n378), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT85), .B1(new_n535), .B2(new_n480), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n503), .A2(new_n311), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n530), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n540), .A2(KEYINPUT17), .A3(new_n518), .A4(new_n526), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n505), .A2(new_n521), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n523), .A2(new_n524), .A3(G179), .A4(new_n345), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n517), .B2(new_n423), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n542), .A2(KEYINPUT18), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT18), .B1(new_n542), .B2(new_n544), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n529), .B(new_n541), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n426), .A2(new_n479), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n331), .A2(G200), .ZN(new_n549));
  INV_X1    g0349(.A(new_n324), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n549), .B(new_n550), .C1(new_n465), .C2(new_n331), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n265), .B1(new_n224), .B2(new_n268), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT88), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n291), .A2(KEYINPUT4), .A3(G244), .A4(new_n286), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n291), .A2(G250), .A3(G1698), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n318), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT4), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n278), .A2(G244), .A3(new_n286), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n554), .B1(new_n267), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n423), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n365), .A2(G77), .ZN(new_n563));
  XNOR2_X1  g0363(.A(KEYINPUT87), .B(KEYINPUT6), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G97), .A2(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n207), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n205), .A2(G107), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  OAI221_X1 g0368(.A(new_n563), .B1(new_n568), .B2(new_n231), .C1(new_n534), .C2(new_n206), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n569), .A2(new_n311), .B1(new_n205), .B2(new_n314), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n315), .A2(G97), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G179), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n554), .B(new_n573), .C1(new_n267), .C2(new_n560), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n562), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n554), .B(G190), .C1(new_n267), .C2(new_n560), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n552), .B(KEYINPUT88), .ZN(new_n577));
  INV_X1    g0377(.A(new_n557), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n559), .A2(new_n558), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n267), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(G200), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n576), .A2(new_n581), .A3(new_n571), .A4(new_n570), .ZN(new_n582));
  XNOR2_X1  g0382(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n583), .A2(new_n266), .A3(new_n205), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n584), .A2(new_n532), .B1(G87), .B2(new_n207), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n583), .B1(new_n369), .B2(new_n205), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n278), .A2(G68), .A3(new_n231), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n311), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n416), .A2(new_n314), .ZN(new_n590));
  INV_X1    g0390(.A(new_n315), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(new_n416), .ZN(new_n592));
  INV_X1    g0392(.A(new_n258), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n267), .A2(new_n593), .A3(G250), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n277), .A2(new_n221), .ZN(new_n595));
  NOR2_X1   g0395(.A1(G238), .A2(G1698), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n596), .B1(new_n396), .B2(G1698), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n595), .B1(new_n278), .B2(new_n597), .ZN(new_n598));
  OAI221_X1 g0398(.A(new_n594), .B1(new_n264), .B2(new_n593), .C1(new_n598), .C2(new_n267), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n599), .A2(G179), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n423), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n592), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n315), .A2(G87), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n589), .A2(new_n590), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(G200), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n604), .B(new_n605), .C1(new_n465), .C2(new_n599), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n575), .A2(new_n582), .A3(new_n602), .A4(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n210), .B1(new_n595), .B2(KEYINPUT23), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT22), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n231), .A2(G87), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n403), .ZN(new_n611));
  NAND2_X1  g0411(.A1(KEYINPUT23), .A2(G107), .ZN(new_n612));
  OR3_X1    g0412(.A1(new_n231), .A2(KEYINPUT23), .A3(G107), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n608), .A2(new_n611), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n278), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n615), .A2(new_n609), .A3(new_n610), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT24), .ZN(new_n617));
  OR3_X1    g0417(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n614), .B2(new_n616), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n311), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n314), .A2(new_n206), .ZN(new_n621));
  XOR2_X1   g0421(.A(new_n621), .B(KEYINPUT25), .Z(new_n622));
  OAI211_X1 g0422(.A(new_n620), .B(new_n622), .C1(new_n206), .C2(new_n591), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n278), .B1(G250), .B2(G1698), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n286), .A2(G257), .ZN(new_n625));
  INV_X1    g0425(.A(G294), .ZN(new_n626));
  OAI22_X1  g0426(.A1(new_n624), .A2(new_n625), .B1(new_n626), .B2(new_n277), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n270), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n263), .A2(G264), .A3(new_n267), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n628), .A2(new_n265), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(KEYINPUT93), .A3(G179), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT93), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n628), .A2(G179), .A3(new_n265), .A4(new_n629), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n632), .B(new_n633), .C1(new_n630), .C2(new_n423), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n623), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n630), .A2(G190), .ZN(new_n636));
  INV_X1    g0436(.A(G200), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n623), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n607), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n335), .A2(new_n548), .A3(new_n551), .A4(new_n640), .ZN(G372));
  NAND3_X1  g0441(.A1(new_n623), .A2(new_n631), .A3(new_n634), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n326), .A2(new_n327), .A3(new_n333), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n607), .A2(new_n639), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n606), .A2(new_n602), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n575), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n647), .A2(new_n575), .A3(KEYINPUT26), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n645), .A2(new_n602), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n548), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n383), .B1(new_n393), .B2(new_n425), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(new_n529), .A3(new_n541), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n545), .A2(new_n546), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n475), .B1(new_n658), .B2(new_n473), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n654), .A2(new_n659), .ZN(G369));
  INV_X1    g0460(.A(new_n551), .ZN(new_n661));
  OR3_X1    g0461(.A1(new_n661), .A2(KEYINPUT95), .A3(new_n334), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n532), .A2(new_n313), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n209), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT94), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT27), .ZN(new_n666));
  OAI21_X1  g0466(.A(G213), .B1(new_n664), .B2(KEYINPUT27), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n664), .B2(KEYINPUT27), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n324), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT95), .B1(new_n661), .B2(new_n334), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n662), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n334), .A2(new_n673), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n642), .A2(new_n672), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n623), .A2(new_n672), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n639), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n677), .B1(new_n679), .B2(new_n642), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n675), .A2(G330), .A3(new_n676), .A4(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n335), .A2(new_n672), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n635), .A2(new_n639), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n677), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT96), .ZN(G399));
  INV_X1    g0489(.A(new_n211), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT97), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT97), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n695), .B(new_n696), .C1(new_n235), .C2(new_n692), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(new_n672), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n653), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT29), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  OAI211_X1 g0503(.A(G179), .B(new_n328), .C1(new_n329), .C2(new_n330), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n628), .A2(new_n629), .ZN(new_n705));
  OR3_X1    g0505(.A1(new_n561), .A2(new_n599), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n561), .A2(new_n599), .A3(new_n705), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n309), .A2(KEYINPUT30), .A3(G179), .A4(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n331), .A2(new_n573), .A3(new_n561), .A4(new_n599), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n707), .B(new_n709), .C1(new_n710), .C2(new_n630), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT31), .B1(new_n711), .B2(new_n672), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n640), .A2(new_n335), .A3(new_n551), .A4(new_n699), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n702), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n701), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n698), .B1(new_n717), .B2(G1), .ZN(G364));
  NAND2_X1  g0518(.A1(new_n675), .A2(new_n676), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n209), .B1(new_n663), .B2(G45), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n691), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n236), .A2(new_n257), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n278), .A2(new_n690), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n727), .B(new_n728), .C1(new_n251), .C2(new_n257), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n291), .A2(G355), .A3(new_n211), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n729), .B(new_n730), .C1(G116), .C2(new_n211), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n232), .B1(G20), .B2(new_n423), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n722), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n532), .A2(new_n465), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n573), .A2(G200), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n465), .A2(G179), .A3(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n231), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n739), .A2(G77), .B1(G97), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n637), .A2(G179), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G20), .A3(G190), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n291), .B1(new_n745), .B2(new_n509), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n573), .A2(new_n637), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n532), .A2(G190), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n746), .B1(new_n749), .B2(G50), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n736), .A2(new_n747), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n743), .B(new_n750), .C1(new_n378), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n736), .A2(new_n573), .A3(new_n637), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT98), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT98), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G159), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT32), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n736), .A2(new_n744), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT99), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G107), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n532), .A2(G190), .A3(new_n737), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n752), .B(new_n763), .C1(G58), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n745), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n761), .A2(G283), .B1(G303), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n291), .B1(new_n765), .B2(G322), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n768), .B(new_n769), .C1(new_n626), .C2(new_n741), .ZN(new_n770));
  INV_X1    g0570(.A(new_n756), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n771), .A2(G329), .B1(G326), .B2(new_n749), .ZN(new_n772));
  XOR2_X1   g0572(.A(KEYINPUT33), .B(G317), .Z(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n751), .B2(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n770), .B(new_n774), .C1(G311), .C2(new_n739), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n732), .B1(new_n766), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n723), .A2(new_n726), .A3(new_n734), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n719), .A2(new_n702), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n675), .A2(G330), .A3(new_n676), .ZN(new_n779));
  INV_X1    g0579(.A(new_n726), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  NAND2_X1  g0583(.A1(new_n422), .A2(new_n672), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n478), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n425), .ZN(new_n786));
  AND4_X1   g0586(.A1(new_n422), .A2(new_n408), .A3(new_n424), .A4(new_n699), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n700), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n787), .B1(new_n425), .B2(new_n785), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n653), .A2(new_n699), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(new_n716), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n780), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n741), .A2(new_n205), .B1(new_n206), .B2(new_n745), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n739), .A2(G116), .B1(new_n749), .B2(G303), .ZN(new_n797));
  INV_X1    g0597(.A(new_n751), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT100), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(KEYINPUT100), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT101), .B(G283), .Z(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n797), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT102), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n771), .A2(G311), .B1(new_n761), .B2(G87), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n806), .A2(new_n403), .A3(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n796), .B(new_n808), .C1(G294), .C2(new_n765), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n798), .A2(G150), .B1(new_n749), .B2(G137), .ZN(new_n810));
  INV_X1    g0610(.A(G143), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n810), .B1(new_n811), .B2(new_n764), .C1(new_n757), .C2(new_n738), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT34), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n812), .A2(new_n813), .B1(G50), .B2(new_n767), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT103), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n615), .B1(new_n771), .B2(G132), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n815), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n761), .A2(G68), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(new_n813), .C2(new_n812), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n817), .B(new_n820), .C1(G58), .C2(new_n742), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n732), .B1(new_n809), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n789), .A2(new_n720), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n732), .A2(new_n720), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n370), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n822), .A2(new_n726), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n795), .A2(new_n826), .ZN(G384));
  NOR2_X1   g0627(.A1(new_n393), .A2(new_n672), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT16), .B1(new_n500), .B2(new_n502), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n521), .B1(new_n538), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n547), .A2(new_n669), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n542), .B1(new_n544), .B2(new_n669), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT37), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(new_n834), .A3(new_n527), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n543), .B(new_n670), .C1(new_n517), .C2(new_n423), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n831), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n527), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT105), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n835), .A2(new_n839), .A3(KEYINPUT105), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n832), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n835), .A2(new_n839), .A3(KEYINPUT105), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT105), .B1(new_n835), .B2(new_n839), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n849), .A2(KEYINPUT38), .A3(new_n832), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT39), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n540), .A2(new_n670), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n547), .A2(KEYINPUT106), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT106), .B1(new_n547), .B2(new_n854), .ZN(new_n856));
  INV_X1    g0656(.A(new_n835), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n834), .B1(new_n833), .B2(new_n527), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n855), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n853), .B(new_n850), .C1(new_n860), .C2(KEYINPUT38), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n829), .B1(new_n852), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n699), .A2(new_n382), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n863), .B(new_n383), .C1(new_n389), .C2(new_n390), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n393), .A2(new_n699), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n792), .B2(new_n788), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n867), .A2(new_n851), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n657), .A2(new_n669), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n862), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n701), .A2(new_n548), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n659), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n870), .B(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT40), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n850), .B1(new_n860), .B2(KEYINPUT38), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n791), .B1(new_n864), .B2(new_n865), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n714), .B2(new_n715), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n874), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n865), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n391), .B1(new_n382), .B2(new_n699), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n789), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n711), .A2(new_n672), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT31), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(new_n715), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n881), .A2(new_n886), .A3(new_n874), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n849), .B2(new_n832), .ZN(new_n888));
  AND4_X1   g0688(.A1(KEYINPUT38), .A2(new_n832), .A3(new_n842), .A4(new_n843), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(G330), .B1(new_n878), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n548), .A2(new_n716), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n856), .ZN(new_n895));
  INV_X1    g0695(.A(new_n859), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n547), .A2(KEYINPUT106), .A3(new_n854), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n889), .B1(new_n845), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n881), .A2(new_n886), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT40), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n877), .A2(new_n874), .A3(new_n851), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n548), .A3(new_n886), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n894), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n873), .B(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n209), .B2(new_n663), .ZN(new_n907));
  OAI21_X1  g0707(.A(G77), .B1(new_n217), .B2(new_n378), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n908), .A2(new_n235), .B1(G50), .B2(new_n378), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(G1), .A3(new_n313), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n568), .B(KEYINPUT35), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(G116), .A3(new_n234), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT104), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT36), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n907), .A2(new_n910), .A3(new_n914), .ZN(G367));
  NAND2_X1  g0715(.A1(new_n572), .A2(new_n672), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n575), .A2(new_n582), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n686), .A2(KEYINPUT42), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n687), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n649), .A2(new_n699), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n683), .A2(new_n918), .A3(new_n684), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT42), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n699), .A2(new_n604), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n925), .A2(new_n602), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n648), .A2(new_n925), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n924), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n686), .B1(new_n685), .B2(KEYINPUT42), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(new_n918), .B1(KEYINPUT42), .B2(new_n922), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n935), .A2(new_n930), .A3(new_n929), .A4(new_n921), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n649), .A2(new_n672), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n917), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n681), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT108), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n933), .A2(new_n936), .A3(KEYINPUT108), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n933), .A2(new_n936), .ZN(new_n946));
  INV_X1    g0746(.A(new_n940), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT107), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n943), .A2(new_n948), .A3(new_n949), .A4(new_n944), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n685), .A2(new_n686), .A3(new_n938), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT45), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n685), .A2(KEYINPUT45), .A3(new_n686), .A4(new_n938), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n938), .B1(new_n685), .B2(new_n686), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n959), .A2(KEYINPUT44), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(KEYINPUT44), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n958), .B(new_n681), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n959), .B(KEYINPUT44), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n681), .B1(new_n964), .B2(new_n958), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n683), .A2(new_n680), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n779), .A2(new_n685), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n685), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n969), .A2(G330), .A3(new_n676), .A4(new_n675), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n717), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT110), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(new_n717), .A3(KEYINPUT110), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n966), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n717), .ZN(new_n977));
  XNOR2_X1  g0777(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n691), .B(new_n978), .Z(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n953), .B1(new_n981), .B2(new_n724), .ZN(new_n982));
  INV_X1    g0782(.A(new_n760), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n801), .A2(G159), .B1(G77), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n984), .B(new_n291), .C1(new_n202), .C2(new_n738), .ZN(new_n985));
  INV_X1    g0785(.A(G150), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n764), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n748), .A2(new_n811), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n745), .A2(new_n217), .ZN(new_n989));
  NOR4_X1   g0789(.A1(new_n985), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(G137), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n990), .B1(new_n378), .B2(new_n741), .C1(new_n991), .C2(new_n756), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT114), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n767), .A2(G116), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT46), .Z(new_n995));
  XNOR2_X1  g0795(.A(KEYINPUT111), .B(G311), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n749), .A2(new_n996), .B1(new_n742), .B2(G107), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT112), .B(G317), .Z(new_n998));
  AOI21_X1  g0798(.A(new_n278), .B1(new_n771), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n205), .B2(new_n760), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n997), .B1(new_n626), .B2(new_n802), .C1(new_n1000), .C2(KEYINPUT113), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n995), .B(new_n1001), .C1(KEYINPUT113), .C2(new_n1000), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n289), .B2(new_n764), .C1(new_n738), .C2(new_n804), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n993), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT47), .Z(new_n1005));
  INV_X1    g0805(.A(new_n732), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n728), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n733), .B1(new_n211), .B2(new_n416), .C1(new_n246), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n722), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n726), .B(new_n1009), .C1(new_n928), .C2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n982), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(G387));
  NOR2_X1   g0814(.A1(new_n680), .A2(new_n1010), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n801), .A2(new_n996), .B1(new_n765), .B2(new_n998), .ZN(new_n1016));
  INV_X1    g0816(.A(G322), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n289), .B2(new_n738), .C1(new_n1017), .C2(new_n748), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT48), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n742), .A2(new_n803), .B1(new_n767), .B2(G294), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT116), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1020), .A2(KEYINPUT116), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT49), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n278), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n983), .A2(G116), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n771), .A2(G326), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n416), .A2(new_n741), .B1(new_n757), .B2(new_n748), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n761), .A2(G97), .B1(G77), .B2(new_n767), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1031), .B(new_n278), .C1(new_n986), .C2(new_n756), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT115), .Z(new_n1033));
  AOI211_X1 g0833(.A(new_n1030), .B(new_n1033), .C1(G50), .C2(new_n765), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n378), .B2(new_n738), .C1(new_n436), .C2(new_n751), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1006), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n410), .A2(new_n202), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT50), .Z(new_n1038));
  AOI21_X1  g0838(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n693), .A3(new_n1039), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n693), .A2(new_n690), .A3(new_n403), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1008), .B1(new_n242), .B2(G45), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n690), .A2(new_n206), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1015), .B(new_n1036), .C1(new_n733), .C2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1046), .A2(new_n726), .B1(new_n725), .B2(new_n971), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n971), .A2(new_n717), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n691), .A3(new_n972), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(G393));
  OAI21_X1  g0850(.A(new_n972), .B1(new_n963), .B2(new_n965), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n976), .A2(new_n691), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT117), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n986), .A2(new_n748), .B1(new_n764), .B2(new_n757), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT51), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n278), .B1(new_n378), .B2(new_n745), .C1(new_n802), .C2(new_n202), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G77), .B2(new_n742), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n761), .A2(G87), .B1(new_n410), .B2(new_n739), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n771), .A2(G143), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1060));
  AND4_X1   g0860(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G311), .A2(new_n765), .B1(new_n749), .B2(G317), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT52), .Z(new_n1063));
  OAI211_X1 g0863(.A(new_n1063), .B(new_n403), .C1(new_n1017), .C2(new_n756), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n742), .A2(G116), .B1(new_n767), .B2(new_n803), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n762), .B(new_n1065), .C1(new_n802), .C2(new_n289), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(G294), .C2(new_n739), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n732), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n733), .B1(new_n205), .B2(new_n211), .C1(new_n1008), .C2(new_n254), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n780), .B1(new_n939), .B2(new_n722), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n966), .B2(new_n725), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1052), .A2(new_n1053), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1053), .B1(new_n1052), .B2(new_n1072), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(G390));
  INV_X1    g0877(.A(KEYINPUT119), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n886), .A2(G330), .A3(new_n791), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n866), .A2(new_n1079), .B1(new_n716), .B2(new_n881), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n792), .A2(new_n788), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1078), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT118), .B1(new_n792), .B2(new_n788), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n792), .A2(KEYINPUT118), .A3(new_n788), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1080), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1079), .A2(new_n866), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n881), .A2(new_n886), .A3(G330), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1089), .A2(KEYINPUT119), .A3(new_n1081), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1083), .A2(new_n1086), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n871), .A2(new_n893), .A3(new_n659), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n852), .B(new_n861), .C1(new_n867), .C2(new_n828), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1085), .A2(new_n1084), .A3(new_n866), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n875), .A2(new_n829), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1088), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1095), .B(new_n1088), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1094), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1091), .A2(new_n1100), .A3(new_n1093), .A4(new_n1101), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n691), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1100), .A2(new_n725), .A3(new_n1101), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(KEYINPUT120), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT120), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1100), .A2(new_n1108), .A3(new_n725), .A4(new_n1101), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n852), .A2(new_n720), .A3(new_n861), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n819), .B1(new_n221), .B2(new_n764), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G283), .B2(new_n749), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n370), .B2(new_n741), .C1(new_n626), .C2(new_n756), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n738), .A2(new_n205), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n802), .A2(new_n206), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n403), .B1(new_n745), .B2(new_n509), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT121), .Z(new_n1118));
  NOR4_X1   g0918(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n801), .A2(G137), .B1(G50), .B2(new_n983), .ZN(new_n1120));
  XOR2_X1   g0920(.A(KEYINPUT54), .B(G143), .Z(new_n1121));
  NAND2_X1  g0921(.A1(new_n739), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n291), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n767), .A2(G150), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(KEYINPUT53), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n771), .A2(G125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(KEYINPUT53), .A2(new_n1124), .B1(new_n742), .B2(G159), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n749), .A2(G128), .ZN(new_n1128));
  INV_X1    g0928(.A(G132), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1127), .B(new_n1128), .C1(new_n1129), .C2(new_n764), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n732), .B1(new_n1119), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n436), .A2(new_n824), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1111), .A2(new_n726), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1105), .A2(new_n1110), .A3(new_n1134), .ZN(G378));
  INV_X1    g0935(.A(KEYINPUT125), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1092), .B(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n870), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT124), .B(KEYINPUT56), .Z(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT55), .B1(new_n473), .B2(new_n476), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT55), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1142), .B(new_n475), .C1(new_n469), .C2(new_n472), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n444), .A2(new_n670), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1144), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n472), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n471), .B1(new_n470), .B2(new_n456), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n476), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1142), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n473), .A2(KEYINPUT55), .A3(new_n476), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1146), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1140), .B1(new_n1145), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1144), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1150), .A2(new_n1146), .A3(new_n1151), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n1155), .A3(new_n1139), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n903), .B2(G330), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(G330), .C1(new_n878), .C2(new_n891), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1138), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n892), .A2(new_n1156), .A3(new_n1153), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n870), .A3(new_n1159), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1104), .A2(new_n1137), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n691), .B1(new_n1164), .B2(KEYINPUT57), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1104), .A2(new_n1137), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1166), .A2(KEYINPUT57), .A3(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1153), .A2(new_n720), .A3(new_n1156), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n739), .A2(G137), .B1(new_n749), .B2(G125), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n798), .A2(G132), .B1(new_n767), .B2(new_n1121), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n742), .A2(G150), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n765), .A2(G128), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT59), .Z(new_n1176));
  NAND2_X1  g0976(.A1(new_n771), .A2(G124), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n266), .A2(new_n259), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT122), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n983), .B2(G159), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1176), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1179), .B(new_n202), .C1(new_n278), .C2(G41), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n416), .A2(new_n738), .B1(new_n751), .B2(new_n205), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT123), .Z(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n370), .B2(new_n745), .C1(new_n206), .C2(new_n764), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n741), .A2(new_n378), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n760), .A2(new_n217), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n771), .A2(G283), .B1(G116), .B2(new_n749), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n259), .A3(new_n615), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1181), .B(new_n1182), .C1(new_n1190), .C2(KEYINPUT58), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1190), .A2(KEYINPUT58), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n732), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n824), .A2(new_n202), .ZN(new_n1194));
  AND4_X1   g0994(.A1(new_n726), .A2(new_n1170), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n1167), .B2(new_n725), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1169), .A2(new_n1196), .ZN(G375));
  NAND4_X1  g0997(.A1(new_n1083), .A2(new_n1086), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1094), .A2(new_n980), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n866), .A2(new_n720), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n824), .A2(new_n378), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n801), .A2(G116), .B1(G283), .B2(new_n765), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n205), .B2(new_n745), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n291), .B(new_n1204), .C1(G294), .C2(new_n749), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n761), .A2(G77), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n771), .A2(G303), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n416), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1208), .A2(new_n742), .B1(G107), .B2(new_n739), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n745), .A2(new_n757), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1187), .B1(new_n801), .B2(new_n1121), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n615), .B1(new_n771), .B2(G128), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n765), .A2(G137), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n748), .A2(new_n1129), .B1(new_n741), .B2(new_n202), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n739), .B2(G150), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1210), .B1(new_n1211), .B2(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n780), .B(new_n1202), .C1(new_n732), .C2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1091), .B2(new_n725), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1199), .A2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT126), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(G381));
  INV_X1    g1023(.A(KEYINPUT127), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(G375), .B(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(G384), .ZN(new_n1226));
  INV_X1    g1026(.A(G378), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1075), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n979), .B1(new_n976), .B2(new_n717), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n952), .B(new_n951), .C1(new_n1230), .C2(new_n725), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1012), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1229), .A2(new_n1231), .A3(new_n1232), .A4(new_n1073), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G396), .A2(G381), .A3(G393), .A4(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1228), .A2(new_n1234), .ZN(G407));
  NAND3_X1  g1035(.A1(new_n1225), .A2(new_n671), .A3(new_n1227), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G213), .B(new_n1236), .C1(new_n1228), .C2(new_n1234), .ZN(G409));
  OAI22_X1  g1037(.A1(new_n982), .A2(new_n1012), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(G393), .B(new_n782), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1238), .A2(new_n1233), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1238), .B2(new_n1233), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G378), .B(new_n1196), .C1(new_n1165), .C2(new_n1168), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1164), .A2(new_n980), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1196), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1227), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(G213), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(G343), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(G2897), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT119), .B1(new_n1089), .B2(new_n1081), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1078), .B(new_n1082), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1256), .A2(KEYINPUT60), .A3(new_n1092), .A4(new_n1086), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT60), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1198), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1257), .A2(new_n1259), .A3(new_n691), .A4(new_n1094), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(G384), .A3(new_n1220), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G384), .B1(new_n1260), .B2(new_n1220), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1253), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1263), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n1261), .A3(new_n1252), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1251), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1261), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1247), .A2(new_n1250), .A3(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT62), .B1(new_n1268), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1249), .B(new_n1269), .C1(new_n1243), .C2(new_n1246), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1242), .B1(new_n1272), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(new_n1250), .B2(new_n1247), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT63), .B1(new_n1279), .B2(new_n1274), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1242), .A2(KEYINPUT61), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1271), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(new_n1281), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1277), .A2(new_n1284), .ZN(G405));
  AOI21_X1  g1085(.A(G378), .B1(new_n1169), .B2(new_n1196), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1243), .ZN(new_n1287));
  OR3_X1    g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1270), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1270), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1288), .A2(new_n1242), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1242), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(G402));
endmodule


