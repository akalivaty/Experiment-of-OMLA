//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT90), .ZN(new_n207));
  AOI21_X1  g006(.A(G8gat), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n202), .A2(new_n204), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n206), .A2(G8gat), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n211), .A2(KEYINPUT89), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(KEYINPUT89), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(KEYINPUT87), .B(G29gat), .Z(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G36gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT14), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT14), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G43gat), .B(G50gat), .Z(new_n224));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT88), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n225), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n219), .A2(new_n221), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT88), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n229), .A2(new_n217), .A3(new_n230), .A4(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n227), .B1(new_n233), .B2(new_n226), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT17), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n227), .B(new_n236), .C1(new_n233), .C2(new_n226), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT91), .B1(new_n214), .B2(new_n234), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT91), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n215), .A2(new_n238), .A3(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n242), .A2(KEYINPUT18), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n243), .B(new_n245), .C1(new_n240), .C2(new_n241), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT18), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n214), .B(new_n234), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n243), .B(KEYINPUT13), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G197gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT11), .ZN(new_n256));
  INV_X1    g055(.A(G169gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n246), .A2(new_n249), .A3(new_n259), .A4(new_n252), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G230gat), .A2(G233gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(G85gat), .A2(G92gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT7), .ZN(new_n266));
  NAND2_X1  g065(.A1(G99gat), .A2(G106gat), .ZN(new_n267));
  INV_X1    g066(.A(G85gat), .ZN(new_n268));
  INV_X1    g067(.A(G92gat), .ZN(new_n269));
  AOI22_X1  g068(.A1(KEYINPUT8), .A2(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G99gat), .B(G106gat), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n271), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G71gat), .A2(G78gat), .ZN(new_n275));
  OR2_X1    g074(.A1(G71gat), .A2(G78gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT9), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G57gat), .B(G64gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(KEYINPUT92), .ZN(new_n280));
  INV_X1    g079(.A(G64gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G57gat), .ZN(new_n282));
  INV_X1    g081(.A(G57gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G64gat), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n282), .A2(new_n284), .A3(KEYINPUT92), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n278), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n275), .B(new_n276), .C1(new_n279), .C2(new_n277), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n286), .A2(KEYINPUT98), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT98), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n274), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n271), .B(new_n272), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT98), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(new_n287), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n264), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n295), .B(KEYINPUT100), .Z(new_n296));
  XNOR2_X1  g095(.A(G120gat), .B(G148gat), .ZN(new_n297));
  INV_X1    g096(.A(G176gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G204gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n264), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT10), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n291), .A2(new_n304), .A3(new_n293), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n294), .A3(new_n304), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT99), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n290), .A2(new_n294), .A3(KEYINPUT99), .A4(new_n304), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n305), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n296), .B(new_n302), .C1(new_n303), .C2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT101), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n310), .A2(new_n303), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n314), .A2(KEYINPUT101), .A3(new_n302), .A4(new_n296), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n264), .B(KEYINPUT102), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n296), .B1(new_n310), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n301), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n263), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n325));
  INV_X1    g124(.A(G120gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n325), .B1(new_n326), .B2(G113gat), .ZN(new_n327));
  INV_X1    g126(.A(G113gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n327), .B(new_n329), .C1(new_n328), .C2(G120gat), .ZN(new_n330));
  INV_X1    g129(.A(G127gat), .ZN(new_n331));
  INV_X1    g130(.A(G134gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G127gat), .A2(G134gat), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT1), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT1), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n328), .A2(G120gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n326), .A2(G113gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n333), .A2(new_n334), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G141gat), .B(G148gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(G155gat), .B2(G162gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n346), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G141gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G148gat), .ZN(new_n352));
  INV_X1    g151(.A(G148gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G141gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G155gat), .B(G162gat), .ZN(new_n356));
  INV_X1    g155(.A(G155gat), .ZN(new_n357));
  INV_X1    g156(.A(G162gat), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT2), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n355), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n350), .A2(new_n360), .ZN(new_n361));
  OR3_X1    g160(.A1(new_n343), .A2(KEYINPUT4), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n361), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n330), .A2(new_n335), .B1(new_n340), .B2(new_n341), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT4), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n355), .A2(new_n356), .A3(new_n359), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n356), .B1(new_n359), .B2(new_n355), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n350), .A2(new_n360), .A3(KEYINPUT75), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n368), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n343), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n350), .A2(new_n360), .A3(KEYINPUT75), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT75), .B1(new_n350), .B2(new_n360), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n375), .B(KEYINPUT3), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n368), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n324), .B(new_n367), .C1(new_n376), .C2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n343), .B1(new_n377), .B2(new_n378), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n365), .ZN(new_n385));
  INV_X1    g184(.A(new_n324), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI211_X1 g187(.A(KEYINPUT77), .B(new_n324), .C1(new_n384), .C2(new_n365), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n382), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n382), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(KEYINPUT5), .A3(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n387), .A2(new_n389), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT5), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n392), .B(new_n382), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G57gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(new_n268), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT6), .ZN(new_n404));
  INV_X1    g203(.A(new_n402), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n394), .A2(new_n397), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n394), .A2(KEYINPUT6), .A3(new_n397), .A4(new_n405), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT80), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n403), .A2(KEYINPUT79), .A3(new_n404), .A4(new_n406), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G8gat), .B(G36gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(new_n281), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(new_n269), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G197gat), .B(G204gat), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT73), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(G211gat), .A2(G218gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(G211gat), .A2(G218gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G211gat), .B(G218gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(new_n422), .A3(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G226gat), .ZN(new_n431));
  INV_X1    g230(.A(G233gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(KEYINPUT29), .ZN(new_n434));
  NOR2_X1   g233(.A1(G183gat), .A2(G190gat), .ZN(new_n435));
  AND2_X1   g234(.A1(G183gat), .A2(G190gat), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(KEYINPUT24), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT65), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n436), .B2(KEYINPUT24), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT65), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n257), .A2(new_n298), .A3(KEYINPUT23), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT23), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(G169gat), .B2(G176gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(G169gat), .A2(G176gat), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  OR2_X1    g250(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n452));
  NAND2_X1  g251(.A1(G183gat), .A2(G190gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n447), .B1(new_n437), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n449), .A2(new_n451), .B1(new_n456), .B2(KEYINPUT25), .ZN(new_n457));
  INV_X1    g256(.A(G190gat), .ZN(new_n458));
  AND2_X1   g257(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT28), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT28), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n463), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT26), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(new_n257), .A3(new_n298), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n446), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n453), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(KEYINPUT67), .A3(new_n453), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT74), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n457), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n437), .A2(new_n455), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n477), .A2(new_n448), .A3(KEYINPUT25), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n440), .B(new_n438), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n447), .B1(new_n479), .B2(new_n437), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n478), .B1(new_n480), .B2(new_n450), .ZN(new_n481));
  INV_X1    g280(.A(new_n473), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT67), .B1(new_n469), .B2(new_n453), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n462), .B(new_n464), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT74), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n434), .B1(new_n476), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(new_n484), .A3(new_n433), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n430), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n475), .B1(new_n457), .B2(new_n474), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n481), .A2(new_n484), .A3(KEYINPUT74), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n433), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n434), .B1(new_n457), .B2(new_n474), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n491), .A2(new_n430), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n417), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(new_n430), .A3(new_n492), .ZN(new_n495));
  INV_X1    g294(.A(new_n487), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n489), .A2(new_n490), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(new_n434), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n495), .B(new_n416), .C1(new_n498), .C2(new_n430), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(new_n499), .A3(KEYINPUT30), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT30), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(new_n417), .C1(new_n488), .C2(new_n493), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n413), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT29), .B1(new_n363), .B2(new_n368), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(new_n430), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G228gat), .A2(G233gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT29), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT3), .B1(new_n430), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n377), .A2(new_n378), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n507), .B(new_n509), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(G197gat), .A2(G204gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(G197gat), .A2(G204gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n428), .B1(new_n516), .B2(new_n419), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n426), .A2(new_n418), .A3(new_n420), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n518), .A3(new_n510), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT81), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT81), .A4(new_n510), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n368), .A3(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n523), .A2(KEYINPUT82), .A3(new_n361), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT82), .B1(new_n523), .B2(new_n361), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n524), .A2(new_n525), .A3(new_n506), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n513), .B1(new_n526), .B2(new_n509), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT83), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(G22gat), .ZN(new_n529));
  XOR2_X1   g328(.A(G78gat), .B(G106gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT31), .ZN(new_n531));
  INV_X1    g330(.A(G50gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n523), .A2(new_n361), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT82), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n523), .A2(KEYINPUT82), .A3(new_n361), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n507), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n508), .ZN(new_n539));
  INV_X1    g338(.A(G22gat), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n539), .A2(new_n540), .A3(new_n513), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n539), .B2(new_n513), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n529), .B(new_n533), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n527), .A2(G22gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n540), .A3(new_n513), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n533), .A2(KEYINPUT83), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT84), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT84), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n543), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n504), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n364), .B1(new_n457), .B2(new_n474), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n481), .A2(new_n484), .A3(new_n343), .ZN(new_n556));
  INV_X1    g355(.A(G227gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(new_n432), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G15gat), .B(G43gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G71gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G99gat), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT33), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(KEYINPUT32), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT69), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n559), .A2(KEYINPUT32), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n562), .B1(new_n559), .B2(new_n563), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT69), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n556), .ZN(new_n573));
  INV_X1    g372(.A(new_n558), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT70), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT71), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n558), .B1(new_n555), .B2(new_n556), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT71), .B1(new_n579), .B2(KEYINPUT70), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT34), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT34), .B1(new_n578), .B2(new_n580), .ZN(new_n582));
  OAI22_X1  g381(.A1(new_n569), .A2(new_n572), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n567), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(KEYINPUT69), .A3(new_n565), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT34), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n577), .B1(new_n575), .B2(new_n576), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n579), .A2(KEYINPUT70), .A3(KEYINPUT71), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT34), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n585), .A2(new_n589), .A3(new_n571), .A4(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n583), .A2(KEYINPUT72), .A3(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n581), .A2(new_n582), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT72), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n585), .A4(new_n571), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(KEYINPUT36), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n583), .A2(new_n597), .A3(new_n591), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n599), .B1(new_n488), .B2(new_n493), .ZN(new_n600));
  OAI211_X1 g399(.A(KEYINPUT37), .B(new_n495), .C1(new_n498), .C2(new_n430), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(new_n601), .A3(new_n416), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT38), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n599), .B1(new_n498), .B2(new_n430), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n491), .A2(new_n492), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n604), .B1(new_n430), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n606), .A2(new_n607), .A3(new_n416), .A4(new_n600), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n603), .A2(new_n494), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n411), .A3(new_n407), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT40), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n367), .B1(new_n376), .B2(new_n381), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n612), .A2(new_n386), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT39), .B1(new_n385), .B2(new_n386), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(KEYINPUT86), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n614), .A2(KEYINPUT86), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n612), .A2(new_n386), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n402), .B1(new_n618), .B2(KEYINPUT39), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n611), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n620), .A2(new_n406), .ZN(new_n621));
  OR3_X1    g420(.A1(new_n617), .A2(new_n611), .A3(new_n619), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n500), .A2(KEYINPUT85), .A3(new_n502), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT85), .B1(new_n500), .B2(new_n502), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n552), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n554), .A2(new_n596), .A3(new_n598), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n592), .A2(new_n595), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n413), .A2(new_n552), .A3(new_n628), .A4(new_n503), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT35), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT80), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n410), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n410), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n407), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT35), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n623), .A2(new_n624), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n583), .A2(new_n591), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n549), .B2(new_n551), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n630), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n323), .B1(new_n627), .B2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT95), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n274), .B1(new_n235), .B2(new_n237), .ZN(new_n646));
  NAND2_X1  g445(.A1(G232gat), .A2(G233gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT94), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n234), .A2(new_n274), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n645), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  NOR4_X1   g453(.A1(new_n646), .A2(new_n654), .A3(KEYINPUT95), .A4(new_n650), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n644), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n238), .A2(new_n291), .ZN(new_n657));
  INV_X1    g456(.A(new_n650), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n652), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT95), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n651), .A2(new_n645), .A3(new_n652), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n643), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n656), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT97), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n656), .A2(new_n662), .A3(new_n663), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n656), .A2(new_n662), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT96), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n648), .A2(new_n649), .ZN(new_n671));
  XOR2_X1   g470(.A(G134gat), .B(G162gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n665), .A2(new_n670), .A3(new_n673), .A4(new_n667), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n293), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT21), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n215), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n681), .B2(new_n215), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n684));
  XNOR2_X1  g483(.A(G155gat), .B(G183gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n683), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(G231gat), .A2(G233gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(new_n331), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G211gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n687), .B(new_n690), .Z(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n642), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n413), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT103), .B(G1gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1324gat));
  INV_X1    g496(.A(G8gat), .ZN(new_n698));
  INV_X1    g497(.A(new_n694), .ZN(new_n699));
  INV_X1    g498(.A(new_n636), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n702));
  AND2_X1   g501(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n703));
  NOR4_X1   g502(.A1(new_n694), .A2(new_n636), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT42), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(KEYINPUT42), .B2(new_n704), .ZN(G1325gat));
  AND3_X1   g505(.A1(new_n596), .A2(KEYINPUT104), .A3(new_n598), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT104), .B1(new_n596), .B2(new_n598), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n699), .A2(G15gat), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n638), .ZN(new_n712));
  AOI21_X1  g511(.A(G15gat), .B1(new_n699), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n711), .A2(new_n713), .ZN(G1326gat));
  NOR2_X1   g513(.A1(new_n694), .A2(new_n552), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT43), .B(G22gat), .Z(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  NAND2_X1  g516(.A1(new_n642), .A2(new_n692), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n675), .A2(new_n676), .ZN(new_n719));
  NOR4_X1   g518(.A1(new_n718), .A2(new_n413), .A3(new_n216), .A4(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT45), .Z(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n610), .A2(new_n552), .A3(new_n625), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n552), .B1(new_n413), .B2(new_n503), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n725), .A2(new_n709), .B1(new_n630), .B2(new_n640), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n722), .B1(new_n726), .B2(new_n719), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n691), .B(KEYINPUT105), .Z(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n323), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n596), .A2(new_n598), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n723), .A2(new_n724), .A3(new_n730), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n629), .A2(KEYINPUT35), .B1(new_n637), .B2(new_n639), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT44), .B(new_n677), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n727), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n216), .B1(new_n734), .B2(new_n413), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n721), .A2(new_n735), .ZN(G1328gat));
  NOR4_X1   g535(.A1(new_n718), .A2(G36gat), .A3(new_n719), .A4(new_n636), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G36gat), .B1(new_n734), .B2(new_n636), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n738), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(G1329gat));
  OAI21_X1  g541(.A(G43gat), .B1(new_n734), .B2(new_n709), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n638), .A2(G43gat), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n642), .A2(new_n692), .A3(new_n677), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748));
  OR3_X1    g547(.A1(new_n734), .A2(new_n748), .A3(new_n552), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n734), .B2(new_n552), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(G50gat), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n718), .A2(new_n719), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(new_n532), .A3(new_n553), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(KEYINPUT48), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G50gat), .B1(new_n734), .B2(new_n552), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(new_n753), .A3(KEYINPUT106), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n756), .B(new_n757), .C1(KEYINPUT106), .C2(new_n755), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n754), .A2(new_n758), .ZN(G1331gat));
  NAND2_X1  g558(.A1(new_n261), .A2(new_n262), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n677), .A2(new_n692), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n321), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT108), .ZN(new_n763));
  INV_X1    g562(.A(new_n726), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(new_n413), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(new_n283), .ZN(G1332gat));
  NOR2_X1   g566(.A1(new_n765), .A2(new_n636), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  AND2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(G1333gat));
  OAI21_X1  g571(.A(G71gat), .B1(new_n765), .B2(new_n709), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n638), .A2(G71gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n765), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g575(.A1(new_n765), .A2(new_n552), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT109), .B(G78gat), .Z(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1335gat));
  NAND2_X1  g578(.A1(new_n692), .A2(new_n263), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT110), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n726), .A2(new_n719), .A3(new_n781), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n782), .A2(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(KEYINPUT51), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n321), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n413), .A2(new_n786), .A3(G85gat), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT112), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n781), .A2(new_n786), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n709), .A2(new_n554), .A3(new_n626), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n719), .B1(new_n791), .B2(new_n641), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n733), .B(new_n790), .C1(new_n792), .C2(KEYINPUT44), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n727), .A2(KEYINPUT111), .A3(new_n733), .A4(new_n790), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n413), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n789), .B1(new_n797), .B2(new_n268), .ZN(G1336gat));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n796), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n269), .B1(new_n799), .B2(new_n700), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n786), .A2(new_n636), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g601(.A(G92gat), .B(new_n802), .C1(new_n783), .C2(new_n784), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT52), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n785), .A2(new_n269), .A3(new_n801), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  OAI21_X1  g605(.A(G92gat), .B1(new_n793), .B2(new_n636), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n808), .ZN(G1337gat));
  NAND2_X1  g608(.A1(new_n799), .A2(new_n710), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n799), .A2(KEYINPUT113), .A3(new_n710), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(G99gat), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(G99gat), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n785), .A2(new_n815), .A3(new_n712), .A4(new_n321), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1338gat));
  INV_X1    g616(.A(G106gat), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n799), .B2(new_n553), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n786), .A2(G106gat), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n552), .B(new_n821), .C1(new_n783), .C2(new_n784), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT53), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n785), .A2(new_n553), .A3(new_n820), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  OAI21_X1  g624(.A(G106gat), .B1(new_n793), .B2(new_n552), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n823), .A2(new_n827), .ZN(G1339gat));
  NOR2_X1   g627(.A1(new_n310), .A2(new_n318), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n302), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n310), .A2(new_n318), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n832), .B(KEYINPUT54), .C1(new_n303), .C2(new_n310), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT55), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(new_n316), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n836), .A2(new_n316), .A3(KEYINPUT114), .A4(new_n837), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n263), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n243), .B1(new_n242), .B2(new_n245), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n250), .A2(new_n251), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n258), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n262), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n321), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n719), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n846), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n675), .B2(new_n676), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n840), .A2(new_n841), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n728), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  NOR4_X1   g653(.A1(new_n677), .A2(new_n692), .A3(new_n321), .A4(new_n760), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n413), .A2(new_n700), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n552), .A2(new_n628), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n859), .A2(new_n328), .A3(new_n860), .A4(new_n760), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n862));
  INV_X1    g661(.A(new_n728), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT55), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT55), .B1(new_n831), .B2(new_n833), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT114), .B1(new_n866), .B2(new_n316), .ZN(new_n867));
  INV_X1    g666(.A(new_n841), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n760), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n677), .B1(new_n869), .B2(new_n847), .ZN(new_n870));
  INV_X1    g669(.A(new_n853), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n863), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n855), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n874), .A2(new_n639), .A3(new_n760), .A4(new_n857), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n862), .B1(new_n875), .B2(G113gat), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n639), .B(new_n857), .C1(new_n854), .C2(new_n855), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n862), .B(G113gat), .C1(new_n877), .C2(new_n263), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n861), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT116), .B(new_n861), .C1(new_n876), .C2(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1340gat));
  OAI21_X1  g683(.A(G120gat), .B1(new_n877), .B2(new_n786), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n859), .A2(new_n860), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n321), .A2(new_n326), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(G1341gat));
  NOR3_X1   g687(.A1(new_n877), .A2(new_n331), .A3(new_n863), .ZN(new_n889));
  INV_X1    g688(.A(new_n886), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n691), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n891), .B2(new_n331), .ZN(G1342gat));
  OR4_X1    g691(.A1(KEYINPUT56), .A2(new_n886), .A3(G134gat), .A4(new_n719), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n332), .A3(new_n677), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n877), .B2(new_n719), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(G1343gat));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n898), .B(new_n553), .C1(new_n854), .C2(new_n855), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n847), .B1(new_n263), .B2(new_n838), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n719), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n853), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n855), .B1(new_n902), .B2(new_n692), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT57), .B1(new_n903), .B2(new_n552), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n709), .A2(new_n857), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT117), .Z(new_n906));
  NAND3_X1  g705(.A1(new_n899), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G141gat), .B1(new_n907), .B2(new_n263), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n710), .A2(new_n552), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n874), .A2(new_n857), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n351), .A3(new_n760), .ZN(new_n912));
  XNOR2_X1  g711(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n908), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n908), .B2(new_n912), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(G1344gat));
  NAND3_X1  g715(.A1(new_n911), .A2(new_n353), .A3(new_n321), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n899), .A2(new_n904), .A3(new_n321), .A4(new_n906), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n919), .A3(G148gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT119), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n918), .A2(new_n922), .A3(new_n919), .A4(G148gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT57), .B1(new_n856), .B2(new_n552), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n851), .A2(new_n316), .A3(new_n866), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n691), .B1(new_n926), .B2(new_n901), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n898), .B(new_n553), .C1(new_n927), .C2(new_n855), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n925), .A2(new_n321), .A3(new_n906), .A4(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n919), .B1(new_n929), .B2(G148gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n917), .B1(new_n924), .B2(new_n930), .ZN(G1345gat));
  NOR3_X1   g730(.A1(new_n907), .A2(new_n357), .A3(new_n863), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n910), .A2(new_n692), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n933), .B(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n935), .B2(new_n357), .ZN(G1346gat));
  OAI21_X1  g735(.A(G162gat), .B1(new_n907), .B2(new_n719), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n911), .A2(new_n358), .A3(new_n677), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1347gat));
  INV_X1    g738(.A(new_n413), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n860), .A2(new_n700), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n942), .B2(KEYINPUT121), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n942), .A2(KEYINPUT121), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n943), .B(new_n944), .C1(new_n854), .C2(new_n855), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n257), .A3(new_n760), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n940), .A2(new_n636), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n874), .A2(KEYINPUT123), .A3(new_n639), .A4(new_n949), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n639), .B(new_n949), .C1(new_n854), .C2(new_n855), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n950), .A2(new_n953), .A3(new_n760), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n948), .B1(new_n257), .B2(new_n954), .ZN(G1348gat));
  NAND4_X1  g754(.A1(new_n950), .A2(new_n953), .A3(G176gat), .A4(new_n321), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n956), .A2(KEYINPUT124), .ZN(new_n957));
  AOI21_X1  g756(.A(G176gat), .B1(new_n947), .B2(new_n321), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n956), .A2(KEYINPUT124), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G1349gat));
  NAND3_X1  g759(.A1(new_n950), .A2(new_n953), .A3(new_n728), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G183gat), .ZN(new_n962));
  INV_X1    g761(.A(new_n945), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n963), .B(new_n691), .C1(new_n460), .C2(new_n459), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT60), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n962), .B(new_n964), .C1(new_n966), .C2(new_n967), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1350gat));
  NAND3_X1  g770(.A1(new_n947), .A2(new_n458), .A3(new_n677), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n950), .A2(new_n953), .A3(new_n677), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n973), .A2(new_n974), .A3(G190gat), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n974), .B1(new_n973), .B2(G190gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(G1351gat));
  INV_X1    g776(.A(new_n928), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n874), .A2(new_n553), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(new_n979), .B2(KEYINPUT57), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n709), .A2(new_n949), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n980), .A2(new_n981), .A3(new_n760), .A4(new_n983), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n925), .A2(new_n760), .A3(new_n928), .A4(new_n983), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT127), .ZN(new_n986));
  XOR2_X1   g785(.A(KEYINPUT126), .B(G197gat), .Z(new_n987));
  NAND3_X1  g786(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n856), .A2(new_n552), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(new_n983), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(new_n760), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n988), .B1(new_n987), .B2(new_n992), .ZN(G1352gat));
  NOR3_X1   g792(.A1(new_n990), .A2(G204gat), .A3(new_n786), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT62), .ZN(new_n995));
  OR2_X1    g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n980), .A2(new_n321), .A3(new_n983), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(G204gat), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n994), .A2(new_n995), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(G1353gat));
  OR3_X1    g799(.A1(new_n990), .A2(G211gat), .A3(new_n692), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n925), .A2(new_n691), .A3(new_n928), .A4(new_n983), .ZN(new_n1002));
  AND3_X1   g801(.A1(new_n1002), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1003));
  AOI21_X1  g802(.A(KEYINPUT63), .B1(new_n1002), .B2(G211gat), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(G1354gat));
  AOI21_X1  g804(.A(G218gat), .B1(new_n991), .B2(new_n677), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n980), .A2(new_n983), .ZN(new_n1007));
  AND2_X1   g806(.A1(new_n677), .A2(G218gat), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(G1355gat));
endmodule


