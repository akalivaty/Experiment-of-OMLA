

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n370, n371, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756;

  BUF_X1 U364 ( .A(n718), .Z(n722) );
  XOR2_X1 U365 ( .A(n346), .B(n636), .Z(n360) );
  XNOR2_X1 U366 ( .A(n641), .B(n640), .ZN(n361) );
  BUF_X1 U367 ( .A(n637), .Z(n346) );
  NOR2_X1 U368 ( .A1(n717), .A2(n692), .ZN(n399) );
  OR2_X1 U369 ( .A1(n754), .A2(n703), .ZN(n439) );
  AND2_X1 U370 ( .A1(n436), .A2(n434), .ZN(n401) );
  OR2_X1 U371 ( .A1(n709), .A2(n410), .ZN(n409) );
  NOR2_X1 U372 ( .A1(n658), .A2(n586), .ZN(n566) );
  OR2_X1 U373 ( .A1(n694), .A2(G902), .ZN(n388) );
  OR2_X1 U374 ( .A1(n645), .A2(G902), .ZN(n495) );
  XNOR2_X1 U375 ( .A(n520), .B(n493), .ZN(n645) );
  INV_X1 U376 ( .A(G146), .ZN(n469) );
  NOR2_X1 U377 ( .A1(G953), .A2(G237), .ZN(n544) );
  INV_X2 U378 ( .A(G953), .ZN(n744) );
  NAND2_X1 U379 ( .A1(n390), .A2(n341), .ZN(n344) );
  OR2_X2 U380 ( .A1(n724), .A2(G902), .ZN(n508) );
  NAND2_X1 U381 ( .A1(n389), .A2(n623), .ZN(n341) );
  NOR2_X2 U382 ( .A1(n367), .A2(n605), .ZN(n607) );
  XNOR2_X2 U383 ( .A(n342), .B(n477), .ZN(n367) );
  NOR2_X2 U384 ( .A1(n604), .A2(n603), .ZN(n342) );
  NAND2_X1 U385 ( .A1(n401), .A2(n343), .ZN(n398) );
  NAND2_X1 U386 ( .A1(n348), .A2(n351), .ZN(n343) );
  XNOR2_X2 U387 ( .A(n588), .B(n532), .ZN(n669) );
  XNOR2_X2 U388 ( .A(n433), .B(G134), .ZN(n557) );
  XNOR2_X2 U389 ( .A(n388), .B(n355), .ZN(n658) );
  XNOR2_X2 U390 ( .A(n344), .B(KEYINPUT45), .ZN(n734) );
  AND2_X4 U391 ( .A1(n403), .A2(n345), .ZN(n718) );
  AND2_X2 U392 ( .A1(n386), .A2(n387), .ZN(n345) );
  AND2_X2 U393 ( .A1(n575), .A2(n579), .ZN(n562) );
  XNOR2_X2 U394 ( .A(n448), .B(n572), .ZN(n755) );
  XNOR2_X2 U395 ( .A(n574), .B(n441), .ZN(n604) );
  XNOR2_X2 U396 ( .A(n607), .B(n606), .ZN(n615) );
  XNOR2_X2 U397 ( .A(n368), .B(n565), .ZN(n693) );
  AND2_X2 U398 ( .A1(n611), .A2(n616), .ZN(n628) );
  XOR2_X1 U399 ( .A(G110), .B(KEYINPUT75), .Z(n525) );
  XNOR2_X1 U400 ( .A(n739), .B(n469), .ZN(n547) );
  NOR2_X1 U401 ( .A1(n639), .A2(n634), .ZN(n531) );
  XNOR2_X2 U402 ( .A(n373), .B(KEYINPUT30), .ZN(n442) );
  XOR2_X2 U403 ( .A(G113), .B(G104), .Z(n543) );
  NOR2_X2 U404 ( .A1(n658), .A2(n472), .ZN(n373) );
  NOR2_X1 U405 ( .A1(n707), .A2(n673), .ZN(n578) );
  INV_X1 U406 ( .A(n671), .ZN(n430) );
  XNOR2_X1 U407 ( .A(n393), .B(n392), .ZN(n711) );
  XNOR2_X1 U408 ( .A(n395), .B(n394), .ZN(n724) );
  XNOR2_X1 U409 ( .A(n414), .B(n547), .ZN(n637) );
  XNOR2_X1 U410 ( .A(n470), .B(n547), .ZN(n395) );
  XNOR2_X1 U411 ( .A(n500), .B(n352), .ZN(n394) );
  INV_X1 U412 ( .A(n668), .ZN(n472) );
  XOR2_X2 U413 ( .A(KEYINPUT10), .B(KEYINPUT68), .Z(n349) );
  NAND2_X2 U414 ( .A1(n374), .A2(n380), .ZN(n375) );
  XNOR2_X2 U415 ( .A(n743), .B(n524), .ZN(n520) );
  XNOR2_X2 U416 ( .A(n557), .B(n487), .ZN(n743) );
  XNOR2_X1 U417 ( .A(G125), .B(G140), .ZN(n501) );
  INV_X1 U418 ( .A(KEYINPUT69), .ZN(n486) );
  XNOR2_X1 U419 ( .A(G119), .B(G116), .ZN(n513) );
  XNOR2_X1 U420 ( .A(n439), .B(KEYINPUT44), .ZN(n389) );
  NOR2_X1 U421 ( .A1(n482), .A2(n696), .ZN(n461) );
  XNOR2_X1 U422 ( .A(n454), .B(G122), .ZN(n554) );
  INV_X1 U423 ( .A(G107), .ZN(n454) );
  XNOR2_X1 U424 ( .A(n543), .B(n481), .ZN(n417) );
  XOR2_X1 U425 ( .A(G143), .B(G122), .Z(n481) );
  XNOR2_X1 U426 ( .A(n546), .B(n545), .ZN(n416) );
  XOR2_X1 U427 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n546) );
  XNOR2_X1 U428 ( .A(n740), .B(G101), .ZN(n524) );
  XNOR2_X1 U429 ( .A(G140), .B(G104), .ZN(n489) );
  AND2_X1 U430 ( .A1(n431), .A2(n428), .ZN(n427) );
  INV_X1 U431 ( .A(n709), .ZN(n563) );
  NAND2_X1 U432 ( .A1(n411), .A2(KEYINPUT107), .ZN(n405) );
  NAND2_X1 U433 ( .A1(n408), .A2(n407), .ZN(n406) );
  BUF_X1 U434 ( .A(n611), .Z(n402) );
  NOR2_X1 U435 ( .A1(n719), .A2(G902), .ZN(n451) );
  XNOR2_X1 U436 ( .A(n602), .B(KEYINPUT94), .ZN(n603) );
  XNOR2_X1 U437 ( .A(n535), .B(n534), .ZN(n538) );
  XOR2_X1 U438 ( .A(KEYINPUT90), .B(KEYINPUT14), .Z(n535) );
  XNOR2_X1 U439 ( .A(n533), .B(KEYINPUT73), .ZN(n534) );
  NAND2_X1 U440 ( .A1(G234), .A2(G237), .ZN(n533) );
  AND2_X1 U441 ( .A1(n669), .A2(n580), .ZN(n438) );
  XNOR2_X1 U442 ( .A(KEYINPUT5), .B(KEYINPUT100), .ZN(n514) );
  XOR2_X1 U443 ( .A(G113), .B(KEYINPUT74), .Z(n515) );
  XNOR2_X1 U444 ( .A(n488), .B(KEYINPUT4), .ZN(n740) );
  NAND2_X1 U445 ( .A1(n634), .A2(n464), .ZN(n463) );
  NAND2_X1 U446 ( .A1(KEYINPUT2), .A2(KEYINPUT65), .ZN(n464) );
  NAND2_X1 U447 ( .A1(n528), .A2(KEYINPUT65), .ZN(n465) );
  AND2_X1 U448 ( .A1(n632), .A2(n467), .ZN(n466) );
  NAND2_X1 U449 ( .A1(n634), .A2(KEYINPUT65), .ZN(n462) );
  XOR2_X1 U450 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n522) );
  INV_X1 U451 ( .A(KEYINPUT77), .ZN(n376) );
  NAND2_X1 U452 ( .A1(n429), .A2(n356), .ZN(n428) );
  OR2_X1 U453 ( .A1(n669), .A2(n432), .ZN(n431) );
  INV_X1 U454 ( .A(KEYINPUT39), .ZN(n435) );
  NAND2_X1 U455 ( .A1(n587), .A2(n413), .ZN(n410) );
  NAND2_X1 U456 ( .A1(n624), .A2(n413), .ZN(n407) );
  OR2_X1 U457 ( .A1(n709), .A2(n586), .ZN(n411) );
  NOR2_X1 U458 ( .A1(n681), .A2(G953), .ZN(n537) );
  XNOR2_X1 U459 ( .A(n423), .B(n476), .ZN(n727) );
  INV_X1 U460 ( .A(n527), .ZN(n476) );
  XNOR2_X1 U461 ( .A(n554), .B(n453), .ZN(n555) );
  INV_X1 U462 ( .A(KEYINPUT103), .ZN(n453) );
  XNOR2_X1 U463 ( .A(n452), .B(n503), .ZN(n553) );
  XNOR2_X1 U464 ( .A(n502), .B(KEYINPUT83), .ZN(n452) );
  XNOR2_X1 U465 ( .A(n415), .B(n549), .ZN(n414) );
  XNOR2_X1 U466 ( .A(n417), .B(n416), .ZN(n415) );
  NAND2_X1 U467 ( .A1(n628), .A2(n618), .ZN(n458) );
  INV_X1 U468 ( .A(KEYINPUT19), .ZN(n441) );
  NOR2_X1 U469 ( .A1(n592), .A2(n595), .ZN(n589) );
  INV_X1 U470 ( .A(n621), .ZN(n419) );
  XNOR2_X1 U471 ( .A(n479), .B(n478), .ZN(n754) );
  INV_X1 U472 ( .A(KEYINPUT32), .ZN(n478) );
  INV_X1 U473 ( .A(KEYINPUT31), .ZN(n392) );
  NAND2_X1 U474 ( .A1(n366), .A2(n665), .ZN(n393) );
  INV_X1 U475 ( .A(KEYINPUT56), .ZN(n445) );
  XOR2_X1 U476 ( .A(n350), .B(n496), .Z(n347) );
  AND2_X1 U477 ( .A1(n438), .A2(n627), .ZN(n348) );
  INV_X1 U478 ( .A(KEYINPUT65), .ZN(n467) );
  XOR2_X1 U479 ( .A(KEYINPUT95), .B(KEYINPUT97), .Z(n350) );
  AND2_X1 U480 ( .A1(n610), .A2(n655), .ZN(n616) );
  NAND2_X1 U481 ( .A1(n608), .A2(n480), .ZN(n586) );
  AND2_X1 U482 ( .A1(n442), .A2(n435), .ZN(n351) );
  XOR2_X1 U483 ( .A(G137), .B(G119), .Z(n352) );
  AND2_X1 U484 ( .A1(n628), .A2(n473), .ZN(n665) );
  INV_X1 U485 ( .A(n468), .ZN(n706) );
  AND2_X1 U486 ( .A1(n442), .A2(n627), .ZN(n353) );
  NOR2_X1 U487 ( .A1(n367), .A2(n473), .ZN(n354) );
  XOR2_X1 U488 ( .A(G472), .B(KEYINPUT72), .Z(n355) );
  XOR2_X1 U489 ( .A(KEYINPUT112), .B(KEYINPUT41), .Z(n356) );
  XOR2_X1 U490 ( .A(KEYINPUT71), .B(KEYINPUT34), .Z(n357) );
  INV_X1 U491 ( .A(KEYINPUT107), .ZN(n413) );
  XOR2_X1 U492 ( .A(KEYINPUT87), .B(KEYINPUT35), .Z(n358) );
  XOR2_X1 U493 ( .A(n694), .B(KEYINPUT62), .Z(n359) );
  XOR2_X1 U494 ( .A(n645), .B(n644), .Z(n362) );
  INV_X1 U495 ( .A(n528), .ZN(n634) );
  AND2_X1 U496 ( .A1(n465), .A2(n463), .ZN(n363) );
  NOR2_X1 U497 ( .A1(n744), .A2(G952), .ZN(n726) );
  INV_X1 U498 ( .A(n726), .ZN(n646) );
  XNOR2_X1 U499 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n364) );
  XOR2_X1 U500 ( .A(KEYINPUT113), .B(KEYINPUT63), .Z(n365) );
  BUF_X1 U501 ( .A(n658), .Z(n471) );
  INV_X1 U502 ( .A(n367), .ZN(n366) );
  NOR2_X2 U503 ( .A1(n682), .A2(n367), .ZN(n620) );
  XNOR2_X1 U504 ( .A(n525), .B(KEYINPUT16), .ZN(n475) );
  NAND2_X1 U505 ( .A1(n398), .A2(n563), .ZN(n368) );
  NAND2_X1 U506 ( .A1(n381), .A2(n399), .ZN(n380) );
  INV_X1 U507 ( .A(n714), .ZN(n384) );
  NAND2_X1 U508 ( .A1(n714), .A2(n474), .ZN(n382) );
  AND2_X2 U509 ( .A1(n590), .A2(n402), .ZN(n714) );
  XNOR2_X2 U510 ( .A(n370), .B(KEYINPUT109), .ZN(n571) );
  NAND2_X1 U511 ( .A1(n568), .A2(n567), .ZN(n370) );
  XNOR2_X1 U512 ( .A(n371), .B(n459), .ZN(n390) );
  NAND2_X1 U513 ( .A1(n460), .A2(n461), .ZN(n371) );
  XNOR2_X1 U514 ( .A(n550), .B(n551), .ZN(n569) );
  NAND2_X1 U515 ( .A1(n406), .A2(n405), .ZN(n412) );
  NAND2_X1 U516 ( .A1(n409), .A2(n618), .ZN(n408) );
  NOR2_X1 U517 ( .A1(n633), .A2(n462), .ZN(n404) );
  NAND2_X1 U518 ( .A1(n378), .A2(n399), .ZN(n374) );
  NAND2_X1 U519 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U520 ( .A1(n633), .A2(n466), .ZN(n386) );
  AND2_X1 U521 ( .A1(n375), .A2(KEYINPUT2), .ZN(n635) );
  XNOR2_X2 U522 ( .A(n375), .B(KEYINPUT86), .ZN(n650) );
  INV_X1 U523 ( .A(n387), .ZN(n391) );
  XNOR2_X2 U524 ( .A(n377), .B(n376), .ZN(n387) );
  NAND2_X1 U525 ( .A1(n734), .A2(n635), .ZN(n377) );
  NOR2_X1 U526 ( .A1(n379), .A2(n591), .ZN(n378) );
  NAND2_X1 U527 ( .A1(n384), .A2(KEYINPUT48), .ZN(n379) );
  NAND2_X1 U528 ( .A1(n591), .A2(n474), .ZN(n383) );
  NAND2_X1 U529 ( .A1(n631), .A2(n734), .ZN(n633) );
  NOR2_X1 U530 ( .A1(n649), .A2(n391), .ZN(n653) );
  NAND2_X1 U531 ( .A1(n711), .A2(n699), .ZN(n630) );
  XNOR2_X1 U532 ( .A(n650), .B(KEYINPUT76), .ZN(n631) );
  NAND2_X1 U533 ( .A1(n571), .A2(n396), .ZN(n707) );
  INV_X1 U534 ( .A(n604), .ZN(n396) );
  NAND2_X1 U535 ( .A1(n616), .A2(n397), .ZN(n512) );
  XNOR2_X1 U536 ( .A(n397), .B(KEYINPUT1), .ZN(n611) );
  XNOR2_X1 U537 ( .A(n397), .B(KEYINPUT108), .ZN(n567) );
  XNOR2_X2 U538 ( .A(n495), .B(n494), .ZN(n397) );
  AND2_X1 U539 ( .A1(n398), .A2(n597), .ZN(n692) );
  NAND2_X1 U540 ( .A1(n718), .A2(G472), .ZN(n695) );
  NAND2_X1 U541 ( .A1(n588), .A2(n668), .ZN(n574) );
  XNOR2_X2 U542 ( .A(n531), .B(n530), .ZN(n588) );
  NOR2_X1 U543 ( .A1(n404), .A2(n363), .ZN(n403) );
  NAND2_X1 U544 ( .A1(n412), .A2(n668), .ZN(n592) );
  XNOR2_X2 U545 ( .A(n349), .B(n501), .ZN(n739) );
  NAND2_X1 U546 ( .A1(n753), .A2(KEYINPUT44), .ZN(n460) );
  XNOR2_X2 U547 ( .A(n418), .B(n358), .ZN(n753) );
  NAND2_X1 U548 ( .A1(n420), .A2(n419), .ZN(n418) );
  XNOR2_X1 U549 ( .A(n620), .B(n357), .ZN(n420) );
  XNOR2_X1 U550 ( .A(n421), .B(n727), .ZN(n639) );
  XNOR2_X1 U551 ( .A(n422), .B(n524), .ZN(n421) );
  XNOR2_X1 U552 ( .A(n457), .B(n523), .ZN(n422) );
  XNOR2_X1 U553 ( .A(n475), .B(n526), .ZN(n423) );
  NAND2_X1 U554 ( .A1(n669), .A2(n668), .ZN(n672) );
  NAND2_X1 U555 ( .A1(n427), .A2(n424), .ZN(n683) );
  NAND2_X1 U556 ( .A1(n669), .A2(n425), .ZN(n424) );
  NOR2_X1 U557 ( .A1(n671), .A2(n426), .ZN(n425) );
  NAND2_X1 U558 ( .A1(n432), .A2(n668), .ZN(n426) );
  NAND2_X1 U559 ( .A1(n430), .A2(n668), .ZN(n429) );
  INV_X1 U560 ( .A(n356), .ZN(n432) );
  XNOR2_X1 U561 ( .A(n433), .B(G125), .ZN(n457) );
  XNOR2_X2 U562 ( .A(n485), .B(n484), .ZN(n433) );
  OR2_X1 U563 ( .A1(n438), .A2(n435), .ZN(n434) );
  NAND2_X1 U564 ( .A1(n437), .A2(KEYINPUT39), .ZN(n436) );
  NAND2_X1 U565 ( .A1(n627), .A2(n442), .ZN(n437) );
  INV_X1 U566 ( .A(n439), .ZN(n622) );
  NAND2_X1 U567 ( .A1(n718), .A2(G469), .ZN(n456) );
  XNOR2_X2 U568 ( .A(n512), .B(KEYINPUT99), .ZN(n627) );
  XNOR2_X1 U569 ( .A(n456), .B(n362), .ZN(n483) );
  INV_X1 U570 ( .A(KEYINPUT48), .ZN(n474) );
  XNOR2_X1 U571 ( .A(n443), .B(n364), .ZN(G60) );
  NAND2_X1 U572 ( .A1(n449), .A2(n646), .ZN(n443) );
  XNOR2_X1 U573 ( .A(n444), .B(n365), .ZN(G57) );
  NAND2_X1 U574 ( .A1(n447), .A2(n646), .ZN(n444) );
  XNOR2_X1 U575 ( .A(n446), .B(n445), .ZN(G51) );
  NAND2_X1 U576 ( .A1(n450), .A2(n646), .ZN(n446) );
  XNOR2_X1 U577 ( .A(n695), .B(n359), .ZN(n447) );
  NAND2_X1 U578 ( .A1(n570), .A2(n571), .ZN(n448) );
  XNOR2_X1 U579 ( .A(n638), .B(n360), .ZN(n449) );
  XNOR2_X1 U580 ( .A(n642), .B(n361), .ZN(n450) );
  XNOR2_X2 U581 ( .A(n451), .B(G478), .ZN(n579) );
  XNOR2_X1 U582 ( .A(n455), .B(n556), .ZN(n559) );
  XNOR2_X1 U583 ( .A(n557), .B(n558), .ZN(n455) );
  INV_X1 U584 ( .A(n402), .ZN(n617) );
  XNOR2_X2 U585 ( .A(n458), .B(n619), .ZN(n682) );
  INV_X1 U586 ( .A(KEYINPUT88), .ZN(n459) );
  NAND2_X1 U587 ( .A1(n353), .A2(n582), .ZN(n468) );
  NAND2_X1 U588 ( .A1(n553), .A2(G221), .ZN(n470) );
  XNOR2_X1 U589 ( .A(n658), .B(KEYINPUT6), .ZN(n618) );
  INV_X1 U590 ( .A(n471), .ZN(n473) );
  INV_X1 U591 ( .A(KEYINPUT0), .ZN(n477) );
  NAND2_X1 U592 ( .A1(n615), .A2(n614), .ZN(n479) );
  AND2_X1 U593 ( .A1(n580), .A2(n655), .ZN(n480) );
  AND2_X1 U594 ( .A1(n630), .A2(n629), .ZN(n482) );
  XNOR2_X1 U595 ( .A(n691), .B(n690), .ZN(G75) );
  XNOR2_X2 U596 ( .A(KEYINPUT80), .B(G143), .ZN(n485) );
  INV_X1 U597 ( .A(G128), .ZN(n484) );
  XNOR2_X1 U598 ( .A(n486), .B(G131), .ZN(n548) );
  XNOR2_X1 U599 ( .A(n548), .B(G137), .ZN(n487) );
  XOR2_X1 U600 ( .A(G146), .B(KEYINPUT64), .Z(n488) );
  XOR2_X1 U601 ( .A(G107), .B(n525), .Z(n492) );
  NAND2_X1 U602 ( .A1(G227), .A2(n744), .ZN(n490) );
  XNOR2_X1 U603 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U604 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U605 ( .A(G469), .B(KEYINPUT70), .ZN(n494) );
  XNOR2_X1 U606 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n496) );
  XOR2_X1 U607 ( .A(KEYINPUT96), .B(KEYINPUT82), .Z(n498) );
  XNOR2_X1 U608 ( .A(G128), .B(G110), .ZN(n497) );
  XNOR2_X1 U609 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U610 ( .A(n347), .B(n499), .ZN(n500) );
  XOR2_X1 U611 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n503) );
  NAND2_X1 U612 ( .A1(G234), .A2(n744), .ZN(n502) );
  XOR2_X1 U613 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n506) );
  XNOR2_X1 U614 ( .A(G902), .B(KEYINPUT15), .ZN(n528) );
  NAND2_X1 U615 ( .A1(G234), .A2(n528), .ZN(n504) );
  XNOR2_X1 U616 ( .A(KEYINPUT20), .B(n504), .ZN(n509) );
  NAND2_X1 U617 ( .A1(G217), .A2(n509), .ZN(n505) );
  XNOR2_X1 U618 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X2 U619 ( .A(n508), .B(n507), .ZN(n610) );
  NAND2_X1 U620 ( .A1(n509), .A2(G221), .ZN(n511) );
  XOR2_X1 U621 ( .A(KEYINPUT98), .B(KEYINPUT21), .Z(n510) );
  XNOR2_X1 U622 ( .A(n511), .B(n510), .ZN(n655) );
  XNOR2_X1 U623 ( .A(n513), .B(KEYINPUT3), .ZN(n527) );
  XNOR2_X1 U624 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U625 ( .A(n527), .B(n516), .Z(n518) );
  NAND2_X1 U626 ( .A1(n544), .A2(G210), .ZN(n517) );
  XNOR2_X1 U627 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U628 ( .A(n520), .B(n519), .ZN(n694) );
  OR2_X1 U629 ( .A1(G237), .A2(G902), .ZN(n529) );
  NAND2_X1 U630 ( .A1(G214), .A2(n529), .ZN(n668) );
  NAND2_X1 U631 ( .A1(G224), .A2(n744), .ZN(n521) );
  XNOR2_X1 U632 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U633 ( .A(n543), .B(n554), .ZN(n526) );
  NAND2_X1 U634 ( .A1(G210), .A2(n529), .ZN(n530) );
  INV_X1 U635 ( .A(KEYINPUT38), .ZN(n532) );
  NAND2_X1 U636 ( .A1(n538), .A2(G952), .ZN(n536) );
  XOR2_X1 U637 ( .A(KEYINPUT91), .B(n536), .Z(n681) );
  XNOR2_X1 U638 ( .A(n537), .B(KEYINPUT92), .ZN(n601) );
  NAND2_X1 U639 ( .A1(G902), .A2(n538), .ZN(n599) );
  NOR2_X1 U640 ( .A1(G900), .A2(n599), .ZN(n539) );
  NAND2_X1 U641 ( .A1(G953), .A2(n539), .ZN(n541) );
  INV_X1 U642 ( .A(KEYINPUT106), .ZN(n540) );
  XNOR2_X1 U643 ( .A(n541), .B(n540), .ZN(n542) );
  OR2_X1 U644 ( .A1(n601), .A2(n542), .ZN(n580) );
  XOR2_X1 U645 ( .A(KEYINPUT13), .B(G475), .Z(n551) );
  NAND2_X1 U646 ( .A1(G214), .A2(n544), .ZN(n545) );
  XOR2_X1 U647 ( .A(n548), .B(KEYINPUT12), .Z(n549) );
  NOR2_X1 U648 ( .A1(G902), .A2(n637), .ZN(n550) );
  INV_X1 U649 ( .A(KEYINPUT102), .ZN(n552) );
  XNOR2_X1 U650 ( .A(n569), .B(n552), .ZN(n575) );
  NAND2_X1 U651 ( .A1(n553), .A2(G217), .ZN(n560) );
  XNOR2_X1 U652 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n558) );
  XNOR2_X1 U653 ( .A(n555), .B(G116), .ZN(n556) );
  XNOR2_X1 U654 ( .A(n560), .B(n559), .ZN(n719) );
  INV_X1 U655 ( .A(KEYINPUT104), .ZN(n561) );
  XNOR2_X2 U656 ( .A(n562), .B(n561), .ZN(n709) );
  XNOR2_X1 U657 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n564) );
  XNOR2_X1 U658 ( .A(n564), .B(KEYINPUT110), .ZN(n565) );
  INV_X1 U659 ( .A(n610), .ZN(n608) );
  XNOR2_X1 U660 ( .A(n566), .B(KEYINPUT28), .ZN(n568) );
  NAND2_X1 U661 ( .A1(n579), .A2(n569), .ZN(n671) );
  INV_X1 U662 ( .A(n683), .ZN(n570) );
  INV_X1 U663 ( .A(KEYINPUT42), .ZN(n572) );
  NOR2_X2 U664 ( .A1(n693), .A2(n755), .ZN(n573) );
  XNOR2_X1 U665 ( .A(n573), .B(KEYINPUT46), .ZN(n585) );
  INV_X1 U666 ( .A(n575), .ZN(n577) );
  INV_X1 U667 ( .A(n579), .ZN(n576) );
  NAND2_X1 U668 ( .A1(n577), .A2(n576), .ZN(n712) );
  NAND2_X1 U669 ( .A1(n712), .A2(n709), .ZN(n629) );
  INV_X1 U670 ( .A(n629), .ZN(n673) );
  XNOR2_X1 U671 ( .A(n578), .B(KEYINPUT47), .ZN(n583) );
  OR2_X1 U672 ( .A1(n579), .A2(n569), .ZN(n621) );
  NAND2_X1 U673 ( .A1(n588), .A2(n580), .ZN(n581) );
  NOR2_X1 U674 ( .A1(n621), .A2(n581), .ZN(n582) );
  AND2_X1 U675 ( .A1(n583), .A2(n468), .ZN(n584) );
  NAND2_X1 U676 ( .A1(n585), .A2(n584), .ZN(n591) );
  INV_X1 U677 ( .A(n618), .ZN(n624) );
  INV_X1 U678 ( .A(n586), .ZN(n587) );
  INV_X1 U679 ( .A(n588), .ZN(n595) );
  XNOR2_X1 U680 ( .A(n589), .B(KEYINPUT36), .ZN(n590) );
  NOR2_X1 U681 ( .A1(n592), .A2(n402), .ZN(n594) );
  INV_X1 U682 ( .A(KEYINPUT43), .ZN(n593) );
  XNOR2_X1 U683 ( .A(n594), .B(n593), .ZN(n596) );
  AND2_X1 U684 ( .A1(n596), .A2(n595), .ZN(n717) );
  INV_X1 U685 ( .A(n712), .ZN(n597) );
  NOR2_X1 U686 ( .A1(G898), .A2(n744), .ZN(n598) );
  XNOR2_X1 U687 ( .A(KEYINPUT93), .B(n598), .ZN(n728) );
  NOR2_X1 U688 ( .A1(n599), .A2(n728), .ZN(n600) );
  NOR2_X1 U689 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U690 ( .A1(n430), .A2(n655), .ZN(n605) );
  XNOR2_X1 U691 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n606) );
  NAND2_X1 U692 ( .A1(n615), .A2(n617), .ZN(n626) );
  NAND2_X1 U693 ( .A1(n471), .A2(n608), .ZN(n609) );
  NOR2_X1 U694 ( .A1(n626), .A2(n609), .ZN(n703) );
  XOR2_X1 U695 ( .A(KEYINPUT105), .B(n610), .Z(n654) );
  NOR2_X1 U696 ( .A1(n654), .A2(n618), .ZN(n612) );
  NAND2_X1 U697 ( .A1(n612), .A2(n402), .ZN(n613) );
  XNOR2_X1 U698 ( .A(KEYINPUT79), .B(n613), .ZN(n614) );
  INV_X1 U699 ( .A(n616), .ZN(n659) );
  XNOR2_X1 U700 ( .A(KEYINPUT89), .B(KEYINPUT33), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n622), .A2(n753), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n654), .ZN(n625) );
  NOR2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n696) );
  NAND2_X1 U704 ( .A1(n354), .A2(n627), .ZN(n699) );
  INV_X1 U705 ( .A(KEYINPUT2), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n718), .A2(G475), .ZN(n638) );
  XOR2_X1 U707 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n636) );
  NAND2_X1 U708 ( .A1(n718), .A2(G210), .ZN(n642) );
  XOR2_X1 U709 ( .A(KEYINPUT81), .B(KEYINPUT55), .Z(n641) );
  XNOR2_X1 U710 ( .A(n639), .B(KEYINPUT54), .ZN(n640) );
  XOR2_X1 U711 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n643) );
  XNOR2_X1 U712 ( .A(n643), .B(KEYINPUT118), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n483), .A2(n646), .ZN(n647) );
  XNOR2_X1 U714 ( .A(n647), .B(KEYINPUT119), .ZN(G54) );
  NOR2_X1 U715 ( .A1(n734), .A2(KEYINPUT2), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n648), .B(KEYINPUT84), .ZN(n649) );
  NOR2_X1 U717 ( .A1(n650), .A2(KEYINPUT2), .ZN(n651) );
  XNOR2_X1 U718 ( .A(n651), .B(KEYINPUT85), .ZN(n652) );
  NAND2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n687) );
  NOR2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U721 ( .A(n656), .B(KEYINPUT49), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n471), .A2(n657), .ZN(n662) );
  NAND2_X1 U723 ( .A1(n617), .A2(n659), .ZN(n660) );
  XOR2_X1 U724 ( .A(KEYINPUT50), .B(n660), .Z(n661) );
  NOR2_X1 U725 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U726 ( .A(n663), .B(KEYINPUT116), .ZN(n664) );
  NOR2_X1 U727 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U728 ( .A(KEYINPUT51), .B(n666), .Z(n667) );
  NOR2_X1 U729 ( .A1(n683), .A2(n667), .ZN(n678) );
  NOR2_X1 U730 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U731 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U732 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U733 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U734 ( .A1(n676), .A2(n682), .ZN(n677) );
  NOR2_X1 U735 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U736 ( .A(n679), .B(KEYINPUT52), .ZN(n680) );
  NOR2_X1 U737 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U738 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U739 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U740 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U741 ( .A1(G953), .A2(n688), .ZN(n691) );
  INV_X1 U742 ( .A(KEYINPUT53), .ZN(n689) );
  XNOR2_X1 U743 ( .A(n689), .B(KEYINPUT117), .ZN(n690) );
  XOR2_X1 U744 ( .A(G134), .B(n692), .Z(G36) );
  XOR2_X1 U745 ( .A(n693), .B(G131), .Z(G33) );
  XOR2_X1 U746 ( .A(G101), .B(n696), .Z(G3) );
  NOR2_X1 U747 ( .A1(n709), .A2(n699), .ZN(n697) );
  XOR2_X1 U748 ( .A(KEYINPUT114), .B(n697), .Z(n698) );
  XNOR2_X1 U749 ( .A(G104), .B(n698), .ZN(G6) );
  NOR2_X1 U750 ( .A1(n712), .A2(n699), .ZN(n701) );
  XNOR2_X1 U751 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n700) );
  XNOR2_X1 U752 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U753 ( .A(G107), .B(n702), .ZN(G9) );
  XOR2_X1 U754 ( .A(n703), .B(G110), .Z(G12) );
  NOR2_X1 U755 ( .A1(n712), .A2(n707), .ZN(n705) );
  XNOR2_X1 U756 ( .A(G128), .B(KEYINPUT29), .ZN(n704) );
  XNOR2_X1 U757 ( .A(n705), .B(n704), .ZN(G30) );
  XOR2_X1 U758 ( .A(G143), .B(n706), .Z(G45) );
  NOR2_X1 U759 ( .A1(n709), .A2(n707), .ZN(n708) );
  XOR2_X1 U760 ( .A(G146), .B(n708), .Z(G48) );
  NOR2_X1 U761 ( .A1(n709), .A2(n711), .ZN(n710) );
  XOR2_X1 U762 ( .A(G113), .B(n710), .Z(G15) );
  NOR2_X1 U763 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U764 ( .A(G116), .B(n713), .Z(G18) );
  XOR2_X1 U765 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n716) );
  XNOR2_X1 U766 ( .A(n714), .B(G125), .ZN(n715) );
  XNOR2_X1 U767 ( .A(n716), .B(n715), .ZN(G27) );
  XOR2_X1 U768 ( .A(G140), .B(n717), .Z(G42) );
  NAND2_X1 U769 ( .A1(n722), .A2(G478), .ZN(n720) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U771 ( .A1(n726), .A2(n721), .ZN(G63) );
  NAND2_X1 U772 ( .A1(n722), .A2(G217), .ZN(n723) );
  XNOR2_X1 U773 ( .A(n723), .B(n724), .ZN(n725) );
  NOR2_X1 U774 ( .A1(n726), .A2(n725), .ZN(G66) );
  XNOR2_X1 U775 ( .A(n727), .B(G101), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U777 ( .A(n730), .B(KEYINPUT123), .ZN(n738) );
  NAND2_X1 U778 ( .A1(G224), .A2(G953), .ZN(n731) );
  XNOR2_X1 U779 ( .A(n731), .B(KEYINPUT122), .ZN(n732) );
  XNOR2_X1 U780 ( .A(KEYINPUT61), .B(n732), .ZN(n733) );
  NAND2_X1 U781 ( .A1(G898), .A2(n733), .ZN(n736) );
  NAND2_X1 U782 ( .A1(n734), .A2(n744), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U784 ( .A(n738), .B(n737), .ZN(G69) );
  XOR2_X1 U785 ( .A(n739), .B(KEYINPUT124), .Z(n741) );
  XNOR2_X1 U786 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U787 ( .A(n743), .B(n742), .ZN(n746) );
  XNOR2_X1 U788 ( .A(n650), .B(n746), .ZN(n745) );
  NAND2_X1 U789 ( .A1(n745), .A2(n744), .ZN(n751) );
  XNOR2_X1 U790 ( .A(n746), .B(G227), .ZN(n747) );
  XNOR2_X1 U791 ( .A(n747), .B(KEYINPUT125), .ZN(n748) );
  NAND2_X1 U792 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U793 ( .A1(G953), .A2(n749), .ZN(n750) );
  NAND2_X1 U794 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U795 ( .A(KEYINPUT126), .B(n752), .ZN(G72) );
  XOR2_X1 U796 ( .A(n753), .B(G122), .Z(G24) );
  XOR2_X1 U797 ( .A(n754), .B(G119), .Z(G21) );
  XNOR2_X1 U798 ( .A(G137), .B(KEYINPUT127), .ZN(n756) );
  XNOR2_X1 U799 ( .A(n756), .B(n755), .ZN(G39) );
endmodule

