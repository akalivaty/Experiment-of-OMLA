//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  AND2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G116), .A2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n207), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G68), .A2(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n219), .C1(G97), .C2(G257), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G1), .B2(G20), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n222));
  XNOR2_X1  g0022(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G1), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n224), .A2(new_n225), .A3(G13), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n213), .B(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n230), .A2(KEYINPUT0), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n203), .A2(new_n205), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n217), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(new_n225), .ZN(new_n235));
  AOI22_X1  g0035(.A1(new_n230), .A2(KEYINPUT0), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  AND3_X1   g0036(.A1(new_n223), .A2(new_n231), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(new_n224), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n217), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n256), .A2(new_n234), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n253), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n224), .A2(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G50), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n255), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT66), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n263), .B(new_n255), .C1(new_n258), .C2(new_n260), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G150), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n225), .A2(G33), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .C1(new_n206), .C2(new_n225), .ZN(new_n269));
  INV_X1    g0069(.A(new_n257), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n262), .A2(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G169), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G223), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n277), .B(new_n280), .C1(G77), .C2(new_n273), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n224), .B1(G41), .B2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n279), .A2(new_n282), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n281), .B(new_n285), .C1(new_n218), .C2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n271), .B1(new_n272), .B2(new_n287), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n287), .A2(G179), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT9), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n262), .A2(new_n264), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n269), .A2(new_n270), .ZN(new_n294));
  OAI211_X1 g0094(.A(KEYINPUT71), .B(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT71), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(new_n271), .B2(KEYINPUT9), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n287), .A2(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n271), .A2(KEYINPUT9), .B1(new_n287), .B2(G200), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n298), .A2(new_n304), .A3(new_n300), .A4(new_n301), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n291), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT72), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n285), .B1(new_n286), .B2(new_n211), .ZN(new_n308));
  AND2_X1   g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  NOR2_X1   g0109(.A1(KEYINPUT3), .A2(G33), .ZN(new_n310));
  OAI211_X1 g0110(.A(G232), .B(new_n275), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT67), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT67), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n273), .A2(new_n313), .A3(G232), .A4(new_n275), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n273), .A2(G238), .A3(G1698), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n309), .A2(new_n310), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G107), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n312), .A2(new_n314), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n308), .B1(new_n318), .B2(new_n280), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT68), .ZN(new_n321));
  AOI211_X1 g0121(.A(new_n321), .B(new_n308), .C1(new_n318), .C2(new_n280), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n272), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n320), .B2(new_n322), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n254), .A2(new_n207), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n253), .A2(new_n234), .A3(new_n256), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(G77), .A3(new_n259), .ZN(new_n329));
  INV_X1    g0129(.A(new_n268), .ZN(new_n330));
  XOR2_X1   g0130(.A(KEYINPUT15), .B(G87), .Z(new_n331));
  INV_X1    g0131(.A(new_n267), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n330), .A2(new_n265), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n225), .B2(new_n207), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT69), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n334), .A2(new_n335), .A3(new_n270), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n335), .B1(new_n334), .B2(new_n270), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n327), .B(new_n329), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n324), .A2(new_n326), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n320), .A2(new_n322), .A3(new_n340), .ZN(new_n341));
  OR3_X1    g0141(.A1(new_n341), .A2(new_n338), .A3(KEYINPUT70), .ZN(new_n342));
  OAI21_X1  g0142(.A(G190), .B1(new_n320), .B2(new_n322), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT70), .B1(new_n341), .B2(new_n338), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n306), .A2(new_n307), .A3(new_n339), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(KEYINPUT77), .A2(G169), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G97), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT73), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT73), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(G33), .A3(G97), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(G226), .B(new_n275), .C1(new_n309), .C2(new_n310), .ZN(new_n353));
  OAI211_X1 g0153(.A(G232), .B(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n280), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT74), .ZN(new_n357));
  INV_X1    g0157(.A(new_n286), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G238), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT74), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n355), .A2(new_n360), .A3(new_n280), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n357), .A2(new_n359), .A3(new_n361), .A4(new_n285), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT13), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n284), .B1(new_n356), .B2(KEYINPUT74), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n359), .A4(new_n361), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n347), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(KEYINPUT14), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n363), .A2(G179), .A3(new_n366), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT12), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n254), .B(new_n202), .C1(KEYINPUT76), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(KEYINPUT76), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n328), .A2(G68), .A3(new_n259), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n265), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n207), .B2(new_n267), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT75), .B(KEYINPUT11), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n377), .A2(new_n270), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n378), .B1(new_n377), .B2(new_n270), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n374), .B(new_n375), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n367), .B2(KEYINPUT14), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n370), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT7), .B1(new_n316), .B2(new_n225), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NOR4_X1   g0186(.A1(new_n309), .A2(new_n310), .A3(new_n386), .A4(G20), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n265), .A2(G159), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n201), .A2(new_n202), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n232), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n388), .A2(KEYINPUT16), .A3(new_n389), .A4(new_n391), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n270), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n328), .A2(new_n259), .A3(new_n330), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n253), .B2(new_n330), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT78), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n218), .A2(G1698), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n402), .B1(G223), .B2(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT79), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n404), .B(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n279), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n279), .A2(G232), .A3(new_n282), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n408), .A2(new_n325), .A3(new_n285), .A4(new_n410), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n407), .A2(new_n284), .A3(new_n409), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(G169), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n401), .A2(new_n414), .A3(KEYINPUT18), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT80), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n401), .A2(new_n414), .A3(KEYINPUT80), .A4(KEYINPUT18), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n401), .A2(new_n414), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n417), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n346), .A2(new_n384), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n363), .A2(G190), .A3(new_n366), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n382), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n340), .B1(new_n363), .B2(new_n366), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n408), .A2(new_n299), .A3(new_n285), .A4(new_n410), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n412), .B2(G200), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n396), .A2(new_n400), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n306), .A2(new_n339), .A3(new_n345), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(KEYINPUT72), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n423), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G116), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n256), .A2(new_n234), .B1(G20), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G283), .ZN(new_n438));
  INV_X1    g0238(.A(G97), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n438), .B(new_n225), .C1(G33), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT20), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n437), .A2(KEYINPUT20), .A3(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n254), .A2(new_n436), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n224), .A2(G33), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n253), .A2(new_n447), .A3(new_n234), .A4(new_n256), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT86), .B1(new_n448), .B2(new_n436), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT86), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n328), .A2(new_n450), .A3(G116), .A4(new_n447), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n445), .A2(new_n446), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n275), .A2(G257), .ZN(new_n453));
  OAI221_X1 g0253(.A(new_n453), .B1(new_n229), .B2(new_n275), .C1(new_n309), .C2(new_n310), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT85), .B(G303), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n316), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n456), .A3(new_n280), .ZN(new_n457));
  AND2_X1   g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n224), .A2(G45), .ZN(new_n461));
  OAI211_X1 g0261(.A(G270), .B(new_n279), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n283), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n459), .B2(new_n458), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n457), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G169), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT21), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n465), .A2(new_n325), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n452), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n444), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT20), .B1(new_n437), .B2(new_n440), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n446), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n451), .A2(new_n449), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT87), .B1(new_n475), .B2(new_n466), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT87), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n452), .A2(new_n477), .A3(G169), .A4(new_n465), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n467), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G107), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G20), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G13), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(G1), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT25), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI22_X1  g0288(.A1(KEYINPUT25), .A2(new_n485), .B1(new_n448), .B2(new_n480), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n225), .B(G87), .C1(new_n309), .C2(new_n310), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT22), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT22), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n273), .A2(new_n492), .A3(new_n225), .A4(G87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n332), .A2(G116), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n481), .B(KEYINPUT23), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT24), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n496), .B1(new_n491), .B2(new_n493), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT24), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n501), .A3(new_n495), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(new_n488), .B(new_n489), .C1(new_n503), .C2(new_n270), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n279), .B1(new_n460), .B2(new_n461), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n229), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n228), .A2(G1698), .ZN(new_n507));
  OAI221_X1 g0307(.A(new_n507), .B1(G250), .B2(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G294), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n279), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n464), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n506), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n325), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(G169), .B2(new_n512), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n470), .B(new_n479), .C1(new_n504), .C2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n273), .A2(new_n225), .A3(G68), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n267), .B2(new_n439), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n349), .A2(new_n351), .ZN(new_n519));
  AOI21_X1  g0319(.A(G20), .B1(new_n519), .B2(KEYINPUT19), .ZN(new_n520));
  NOR3_X1   g0320(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n516), .B(new_n518), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n270), .ZN(new_n523));
  INV_X1    g0323(.A(new_n331), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n254), .ZN(new_n525));
  INV_X1    g0325(.A(new_n448), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G87), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n523), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(G33), .A2(G41), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n461), .B(G250), .C1(new_n529), .C2(new_n234), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G238), .B(new_n275), .C1(new_n309), .C2(new_n310), .ZN(new_n532));
  OAI211_X1 g0332(.A(G244), .B(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI211_X1 g0335(.A(new_n463), .B(new_n531), .C1(new_n535), .C2(new_n280), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n340), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT84), .B1(new_n528), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(G190), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(new_n280), .ZN(new_n540));
  INV_X1    g0340(.A(new_n463), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n530), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G200), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n522), .A2(new_n270), .B1(new_n254), .B2(new_n524), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT84), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .A4(new_n527), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n538), .A2(new_n539), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n526), .A2(new_n331), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n523), .A2(new_n525), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n536), .A2(new_n325), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n549), .B(new_n550), .C1(G169), .C2(new_n536), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n498), .A2(KEYINPUT24), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n501), .B1(new_n500), .B2(new_n495), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n270), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n510), .ZN(new_n556));
  INV_X1    g0356(.A(new_n505), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G264), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n556), .A2(new_n558), .A3(new_n299), .A4(new_n464), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n512), .B2(G200), .ZN(new_n560));
  INV_X1    g0360(.A(new_n488), .ZN(new_n561));
  INV_X1    g0361(.A(new_n489), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n555), .A2(new_n560), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n465), .A2(G200), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n475), .B(new_n564), .C1(new_n299), .C2(new_n465), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n515), .A2(new_n552), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(G107), .B1(new_n385), .B2(new_n387), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT6), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n439), .A2(new_n480), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G97), .A2(G107), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n480), .A2(KEYINPUT6), .A3(G97), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n265), .A2(G77), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n568), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n270), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n253), .A2(G97), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n526), .B2(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n273), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n582));
  OAI21_X1  g0382(.A(G244), .B1(new_n309), .B2(new_n310), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT4), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n585), .A3(new_n438), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n273), .A2(G250), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n275), .B1(new_n587), .B2(KEYINPUT4), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n280), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n464), .B1(new_n505), .B2(new_n228), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n272), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(new_n325), .A3(new_n591), .ZN(new_n594));
  AND4_X1   g0394(.A1(KEYINPUT82), .A2(new_n581), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  OR2_X1    g0395(.A1(KEYINPUT3), .A2(G33), .ZN(new_n596));
  NAND2_X1  g0396(.A1(KEYINPUT3), .A2(G33), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n213), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(G1698), .B1(new_n598), .B2(new_n584), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n583), .A2(new_n584), .B1(G33), .B2(G283), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n600), .A3(new_n582), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n590), .B1(new_n601), .B2(new_n280), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n578), .A2(new_n580), .B1(new_n602), .B2(new_n325), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT82), .B1(new_n603), .B2(new_n593), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT83), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT81), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n589), .A2(G190), .A3(new_n591), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n578), .A3(new_n580), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n602), .A2(new_n340), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n592), .A2(G200), .ZN(new_n612));
  INV_X1    g0412(.A(new_n580), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n577), .B2(new_n270), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n612), .A2(KEYINPUT81), .A3(new_n614), .A4(new_n608), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n605), .A2(new_n606), .A3(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n611), .A2(new_n615), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT82), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n386), .B1(new_n273), .B2(G20), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n316), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n622), .A2(G107), .B1(G20), .B2(new_n574), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n257), .B1(new_n623), .B2(new_n576), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n594), .B1(new_n624), .B2(new_n613), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n602), .A2(G169), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n619), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n603), .A2(KEYINPUT82), .A3(new_n593), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT83), .B1(new_n618), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n567), .B1(new_n617), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n435), .A2(new_n631), .ZN(G372));
  AND2_X1   g0432(.A1(new_n423), .A2(new_n434), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT88), .B1(new_n536), .B2(G169), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT88), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n542), .A2(new_n635), .A3(new_n272), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n634), .A2(new_n549), .A3(new_n550), .A4(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n539), .A2(new_n543), .A3(new_n544), .A4(new_n527), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n637), .A2(new_n593), .A3(new_n603), .A4(new_n638), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n640));
  INV_X1    g0440(.A(new_n637), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n547), .A2(new_n551), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n605), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(KEYINPUT26), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT89), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n563), .A2(new_n638), .A3(new_n637), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n489), .B1(new_n503), .B2(new_n270), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n514), .B1(new_n647), .B2(new_n561), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n479), .A2(new_n470), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n646), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n605), .A2(new_n616), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n645), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n637), .A2(new_n638), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n563), .B(new_n655), .C1(new_n648), .C2(new_n650), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n611), .B(new_n615), .C1(new_n595), .C2(new_n604), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT89), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n640), .B(new_n644), .C1(new_n654), .C2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n633), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT90), .ZN(new_n661));
  AOI211_X1 g0461(.A(new_n420), .B(new_n413), .C1(new_n396), .C2(new_n400), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT18), .B1(new_n401), .B2(new_n414), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n339), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n370), .B2(new_n383), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n665), .B1(new_n667), .B2(new_n432), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n303), .A2(new_n305), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n291), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n661), .A2(new_n670), .ZN(G369));
  NOR2_X1   g0471(.A1(new_n483), .A2(G20), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n484), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT92), .Z(new_n675));
  NOR2_X1   g0475(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT91), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n475), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(new_n650), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n683), .A2(new_n565), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n563), .B1(new_n504), .B2(new_n681), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n649), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n648), .A2(new_n681), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n650), .A2(new_n681), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(new_n648), .B2(new_n681), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(G399));
  NOR2_X1   g0495(.A1(new_n227), .A2(G41), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n521), .A2(new_n436), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n696), .A2(new_n697), .A3(new_n224), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n233), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  AND3_X1   g0500(.A1(new_n563), .A2(new_n638), .A3(new_n637), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n515), .A2(new_n701), .A3(new_n618), .A4(new_n629), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT26), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n642), .A2(new_n703), .A3(new_n605), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n641), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n681), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT94), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n706), .A2(KEYINPUT94), .A3(new_n681), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(KEYINPUT29), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n567), .B(new_n681), .C1(new_n617), .C2(new_n630), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT93), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n469), .A2(new_n556), .A3(new_n558), .A4(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n714), .A2(KEYINPUT93), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n602), .A2(new_n536), .ZN(new_n718));
  OR3_X1    g0518(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n465), .A2(new_n325), .ZN(new_n720));
  OR4_X1    g0520(.A1(new_n536), .A2(new_n602), .A3(new_n720), .A4(new_n512), .ZN(new_n721));
  OAI22_X1  g0521(.A1(new_n716), .A2(new_n718), .B1(KEYINPUT93), .B2(new_n714), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n680), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT31), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n726), .A3(new_n680), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n712), .B1(new_n713), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n659), .A2(new_n731), .A3(new_n681), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n711), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n700), .B1(new_n734), .B2(G1), .ZN(G364));
  INV_X1    g0535(.A(new_n696), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n672), .A2(G45), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(G1), .A3(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G311), .ZN(new_n739));
  NAND2_X1  g0539(.A1(G20), .A2(G179), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT96), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G190), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n299), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G322), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n739), .A2(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n299), .A2(new_n340), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n225), .A2(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n273), .B1(new_n751), .B2(G303), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n749), .A2(new_n742), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G329), .ZN(new_n755));
  INV_X1    g0555(.A(G294), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n744), .A2(new_n325), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n752), .B(new_n755), .C1(new_n756), .C2(new_n759), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n741), .A2(KEYINPUT97), .A3(new_n748), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT97), .B1(new_n741), .B2(new_n748), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n747), .B(new_n760), .C1(new_n764), .C2(G326), .ZN(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n340), .A2(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n749), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n741), .A2(KEYINPUT98), .A3(new_n767), .ZN(new_n769));
  AOI21_X1  g0569(.A(KEYINPUT98), .B1(new_n741), .B2(new_n767), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  XOR2_X1   g0572(.A(KEYINPUT33), .B(G317), .Z(new_n773));
  OAI221_X1 g0573(.A(new_n765), .B1(new_n766), .B2(new_n768), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT99), .Z(new_n775));
  OAI21_X1  g0575(.A(new_n273), .B1(new_n745), .B2(new_n201), .ZN(new_n776));
  INV_X1    g0576(.A(new_n743), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n777), .A2(G77), .B1(G87), .B2(new_n751), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n480), .B2(new_n768), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n776), .B(new_n779), .C1(G97), .C2(new_n758), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G50), .A2(new_n764), .B1(new_n771), .B2(G68), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n753), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT32), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n780), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n775), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n234), .B1(G20), .B2(new_n272), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n738), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n227), .A2(new_n273), .ZN(new_n789));
  INV_X1    g0589(.A(G45), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n233), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n789), .B(new_n791), .C1(new_n248), .C2(new_n790), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n273), .A2(new_n226), .A3(G355), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n792), .B(new_n793), .C1(G116), .C2(new_n226), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT95), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n787), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n798), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n788), .B(new_n800), .C1(new_n684), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n684), .A2(G330), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n685), .A2(new_n738), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(G396));
  INV_X1    g0605(.A(KEYINPUT100), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n339), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT100), .A4(new_n338), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n809), .A2(new_n345), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n659), .A2(new_n681), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n659), .A2(new_n681), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n338), .A2(new_n680), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n809), .A2(new_n345), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n666), .A2(new_n680), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n811), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n730), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(KEYINPUT101), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(KEYINPUT101), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n817), .A2(new_n730), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n819), .A2(new_n738), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n745), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n771), .A2(G150), .B1(G143), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n825), .B2(new_n763), .C1(new_n782), .C2(new_n743), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT34), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n273), .B1(new_n753), .B2(new_n828), .C1(new_n217), .C2(new_n750), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G58), .B2(new_n758), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n827), .B(new_n830), .C1(new_n202), .C2(new_n768), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n759), .A2(new_n439), .B1(new_n739), .B2(new_n753), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n316), .B1(new_n768), .B2(new_n212), .C1(new_n480), .C2(new_n750), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n756), .B2(new_n745), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G303), .B2(new_n764), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n836), .B1(new_n436), .B2(new_n743), .C1(new_n766), .C2(new_n772), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n787), .A2(new_n795), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n838), .A2(new_n787), .B1(new_n207), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n738), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n840), .B(new_n841), .C1(new_n797), .C2(new_n816), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n822), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G384));
  XNOR2_X1  g0644(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n678), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n401), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n419), .A2(new_n848), .A3(new_n430), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT104), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n419), .A2(new_n848), .A3(new_n852), .A4(new_n430), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT105), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n396), .A2(new_n400), .A3(new_n429), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n678), .B1(new_n396), .B2(new_n400), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT105), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(new_n852), .A4(new_n419), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT104), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n849), .A2(new_n860), .A3(KEYINPUT37), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n851), .A2(new_n854), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT17), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n430), .B(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n856), .B1(new_n664), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n846), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n848), .B1(new_n422), .B2(new_n431), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n852), .B1(new_n857), .B2(new_n419), .ZN(new_n868));
  INV_X1    g0668(.A(new_n853), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n867), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n425), .A2(new_n426), .B1(new_n382), .B2(new_n681), .ZN(new_n874));
  INV_X1    g0674(.A(new_n369), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n875), .A2(new_n367), .A3(KEYINPUT14), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n367), .A2(KEYINPUT14), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n381), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n874), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n370), .A2(new_n383), .A3(new_n681), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n815), .B2(new_n814), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n713), .A2(new_n728), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT106), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT40), .B1(new_n873), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n871), .B1(new_n867), .B2(new_n870), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n850), .A2(new_n853), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n663), .B1(new_n662), .B2(KEYINPUT80), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n864), .B1(new_n888), .B2(new_n417), .ZN(new_n889));
  OAI211_X1 g0689(.A(KEYINPUT38), .B(new_n887), .C1(new_n889), .C2(new_n848), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(KEYINPUT106), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n892), .A2(new_n883), .A3(new_n894), .A4(new_n882), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n885), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n633), .A2(new_n883), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(G330), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n809), .A2(new_n680), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n811), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n886), .A2(new_n890), .ZN(new_n903));
  INV_X1    g0703(.A(new_n881), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n664), .A2(new_n678), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n866), .B2(new_n872), .ZN(new_n908));
  INV_X1    g0708(.A(new_n880), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n886), .A2(new_n890), .A3(KEYINPUT39), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n905), .A2(new_n906), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n435), .B1(new_n711), .B2(new_n732), .ZN(new_n913));
  INV_X1    g0713(.A(new_n670), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n912), .B(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n899), .B(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n224), .B2(new_n672), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n436), .B1(new_n574), .B2(KEYINPUT35), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(new_n235), .C1(KEYINPUT35), .C2(new_n574), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT36), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n233), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(G50), .B2(new_n202), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(G1), .A3(new_n483), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT102), .Z(new_n925));
  NAND3_X1  g0725(.A1(new_n918), .A2(new_n921), .A3(new_n925), .ZN(G367));
  NAND2_X1  g0726(.A1(new_n737), .A2(G1), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n653), .B1(new_n614), .B2(new_n681), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n680), .A2(new_n603), .A3(new_n593), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n694), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT45), .ZN(new_n932));
  OR3_X1    g0732(.A1(new_n694), .A2(KEYINPUT44), .A3(new_n930), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT44), .B1(new_n694), .B2(new_n930), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n690), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT45), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n931), .B(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n938), .A2(new_n691), .A3(new_n934), .A4(new_n933), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n693), .A2(KEYINPUT108), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n689), .A2(new_n692), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n693), .A2(KEYINPUT108), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT109), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n685), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n734), .B1(new_n940), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n696), .B(KEYINPUT41), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n927), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n693), .A2(new_n653), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT42), .ZN(new_n954));
  INV_X1    g0754(.A(new_n528), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n655), .B1(new_n955), .B2(new_n681), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n641), .A2(new_n528), .A3(new_n680), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n930), .A2(new_n648), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n680), .B1(new_n959), .B2(new_n629), .ZN(new_n960));
  OR4_X1    g0760(.A1(KEYINPUT43), .A2(new_n954), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n958), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT43), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(new_n954), .C2(new_n960), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n690), .A2(new_n930), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n961), .A2(new_n968), .A3(new_n966), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT107), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n952), .A2(new_n970), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n764), .A2(G143), .ZN(new_n976));
  INV_X1    g0776(.A(G150), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n217), .A2(new_n743), .B1(new_n745), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n768), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(G77), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n771), .A2(G159), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n273), .B1(new_n753), .B2(new_n825), .C1(new_n201), .C2(new_n750), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G68), .B2(new_n758), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n976), .A2(new_n980), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G311), .A2(new_n764), .B1(new_n771), .B2(G294), .ZN(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n316), .B1(new_n753), .B2(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n745), .A2(new_n455), .B1(new_n439), .B2(new_n768), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(G283), .C2(new_n777), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n985), .B(new_n989), .C1(new_n480), .C2(new_n759), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n750), .A2(new_n436), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT46), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n984), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n787), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n962), .A2(new_n798), .ZN(new_n996));
  INV_X1    g0796(.A(new_n789), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n799), .B1(new_n226), .B2(new_n524), .C1(new_n244), .C2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT110), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n995), .A2(new_n996), .A3(new_n841), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n975), .A2(new_n1000), .ZN(G387));
  NAND2_X1  g0801(.A1(new_n948), .A2(new_n733), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n947), .A2(new_n734), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(new_n696), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n768), .A2(new_n436), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n273), .B1(new_n754), .B2(G326), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n771), .A2(G311), .B1(G317), .B2(new_n823), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n746), .B2(new_n763), .C1(new_n455), .C2(new_n743), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT48), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n766), .B2(new_n759), .C1(new_n756), .C2(new_n750), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1006), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1005), .B(new_n1012), .C1(new_n1011), .C2(new_n1010), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n751), .A2(G77), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n743), .B2(new_n202), .C1(new_n217), .C2(new_n745), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n273), .B1(new_n753), .B2(new_n977), .C1(new_n439), .C2(new_n768), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n331), .B2(new_n758), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n763), .B2(new_n782), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1015), .B(new_n1018), .C1(new_n330), .C2(new_n771), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n787), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n997), .B1(new_n241), .B2(G45), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n268), .A2(G50), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT111), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1023), .A2(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n697), .B1(new_n1023), .B2(KEYINPUT50), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(G68), .A2(G77), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n790), .A4(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1021), .A2(new_n1027), .B1(new_n480), .B2(new_n227), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n697), .A2(new_n226), .A3(new_n273), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n689), .A2(new_n798), .B1(new_n799), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1020), .A2(new_n841), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n927), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1004), .B(new_n1032), .C1(new_n1033), .C2(new_n948), .ZN(G393));
  AOI21_X1  g0834(.A(new_n736), .B1(new_n940), .B2(new_n1003), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n940), .B2(new_n1003), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n936), .A2(new_n939), .A3(new_n927), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n772), .A2(new_n217), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n273), .B1(new_n768), .B2(new_n212), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G143), .B2(new_n754), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n207), .B2(new_n759), .C1(new_n268), .C2(new_n743), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n763), .A2(new_n977), .B1(new_n782), .B2(new_n745), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT113), .Z(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1038), .B(new_n1041), .C1(new_n1044), .C2(KEYINPUT51), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(KEYINPUT51), .B2(new_n1044), .C1(new_n202), .C2(new_n750), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n763), .A2(new_n986), .B1(new_n739), .B2(new_n745), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT52), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n316), .B1(new_n768), .B2(new_n480), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G283), .B2(new_n751), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n436), .B2(new_n759), .C1(new_n756), .C2(new_n743), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n455), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(new_n1052), .B2(new_n771), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1048), .B(new_n1053), .C1(new_n746), .C2(new_n753), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1046), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n738), .B1(new_n1055), .B2(new_n787), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n799), .B1(new_n439), .B2(new_n226), .C1(new_n251), .C2(new_n997), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n801), .C2(new_n930), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1036), .A2(new_n1037), .A3(new_n1058), .ZN(G390));
  INV_X1    g0859(.A(KEYINPUT116), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n904), .B1(new_n729), .B2(new_n816), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1061), .A2(KEYINPUT114), .B1(new_n811), .B2(new_n901), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT114), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n729), .A2(new_n882), .ZN(new_n1064));
  AOI221_X4 g0864(.A(new_n712), .B1(new_n814), .B2(new_n815), .C1(new_n713), .C2(new_n728), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1063), .B(new_n1064), .C1(new_n1065), .C2(new_n904), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n709), .A2(new_n710), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n900), .B1(new_n1067), .B2(new_n816), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n883), .A2(G330), .A3(new_n816), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1069), .A2(new_n881), .B1(new_n729), .B2(new_n882), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1062), .A2(new_n1066), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n710), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT94), .B1(new_n706), .B2(new_n681), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1072), .A2(new_n1073), .A3(new_n731), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n659), .A2(new_n731), .A3(new_n681), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n633), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n633), .A2(G330), .A3(new_n883), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n1077), .A3(new_n670), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT115), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1080));
  AOI221_X4 g0880(.A(KEYINPUT114), .B1(new_n729), .B2(new_n882), .C1(new_n1069), .C2(new_n881), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1069), .A2(KEYINPUT114), .A3(new_n881), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n902), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1080), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT115), .ZN(new_n1085));
  AND4_X1   g0885(.A1(G330), .A2(new_n423), .A3(new_n434), .A4(new_n883), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n913), .A2(new_n914), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1079), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n873), .A2(new_n909), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1068), .B2(new_n881), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n908), .A2(new_n910), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n881), .B1(new_n811), .B2(new_n901), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n909), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1091), .A2(new_n1094), .A3(new_n1064), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1064), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1060), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1064), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1091), .A2(new_n1094), .A3(new_n1064), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1103), .A2(KEYINPUT116), .A3(new_n1088), .A4(new_n1079), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1089), .A2(new_n1097), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1098), .A2(new_n696), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1092), .A2(new_n796), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n316), .B1(new_n754), .B2(G125), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1108), .B1(new_n217), .B2(new_n768), .C1(new_n782), .C2(new_n759), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n751), .A2(G150), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT53), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(G132), .C2(new_n823), .ZN(new_n1112));
  XOR2_X1   g0912(.A(KEYINPUT54), .B(G143), .Z(new_n1113));
  NAND2_X1  g0913(.A1(new_n777), .A2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G128), .A2(new_n764), .B1(new_n771), .B2(G137), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n764), .A2(G283), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n439), .A2(new_n743), .B1(new_n745), .B2(new_n436), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G77), .B2(new_n758), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n771), .A2(G107), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n316), .B1(new_n753), .B2(new_n756), .C1(new_n212), .C2(new_n750), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G68), .B2(new_n979), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1116), .A2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1124), .A2(new_n787), .B1(new_n268), .B2(new_n839), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1107), .A2(new_n841), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1097), .B2(new_n927), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1106), .A2(new_n1127), .ZN(G378));
  NAND2_X1  g0928(.A1(new_n823), .A2(G128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n825), .B2(new_n743), .C1(new_n977), .C2(new_n759), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n764), .B2(G125), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n751), .A2(new_n1113), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT118), .Z(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(new_n828), .C2(new_n772), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1136));
  AOI21_X1  g0936(.A(G33), .B1(new_n979), .B2(G159), .ZN(new_n1137));
  AOI21_X1  g0937(.A(G41), .B1(new_n754), .B2(G124), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n217), .B1(new_n309), .B2(G41), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1014), .B1(new_n201), .B2(new_n768), .C1(new_n766), .C2(new_n753), .ZN(new_n1141));
  AOI211_X1 g0941(.A(G41), .B(new_n1141), .C1(G68), .C2(new_n758), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n316), .B1(new_n743), .B2(new_n524), .C1(new_n480), .C2(new_n745), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n771), .B2(G97), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(new_n436), .C2(new_n763), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1146));
  XNOR2_X1  g0946(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1139), .A2(new_n1140), .A3(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1148), .A2(new_n787), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT119), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n306), .B(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n678), .A2(new_n271), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n738), .B(new_n1149), .C1(new_n1159), .C2(new_n796), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n839), .A2(new_n217), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT106), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n713), .A2(new_n728), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n816), .A2(new_n904), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n848), .B1(new_n665), .B2(new_n431), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n849), .A2(new_n860), .A3(KEYINPUT37), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n860), .B1(new_n849), .B2(KEYINPUT37), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n854), .A2(new_n859), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1167), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n890), .B1(new_n1172), .B2(new_n846), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n891), .B1(new_n1166), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n895), .ZN(new_n1175));
  OAI21_X1  g0975(.A(G330), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT120), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1159), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1176), .A2(new_n912), .A3(new_n1177), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n912), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n886), .A2(new_n890), .A3(KEYINPUT39), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n907), .B2(new_n1173), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1183), .A2(new_n909), .B1(new_n1093), .B2(new_n903), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n712), .B1(new_n885), .B2(new_n895), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1184), .B(new_n906), .C1(new_n1185), .C2(KEYINPUT120), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1158), .B1(new_n1185), .B2(KEYINPUT120), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1176), .A2(new_n912), .A3(new_n1177), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1181), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1162), .B1(new_n1190), .B2(new_n1033), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1078), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n736), .B1(new_n1193), .B2(KEYINPUT57), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT57), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1191), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(G375));
  NAND2_X1  g0998(.A1(new_n1084), .A2(new_n927), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT121), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n881), .A2(new_n795), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n763), .A2(new_n756), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n759), .A2(new_n524), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n480), .A2(new_n743), .B1(new_n745), .B2(new_n766), .ZN(new_n1204));
  INV_X1    g1004(.A(G303), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n316), .B1(new_n753), .B2(new_n1205), .C1(new_n207), .C2(new_n768), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n439), .B2(new_n750), .C1(new_n436), .C2(new_n772), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n745), .A2(new_n825), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G159), .A2(new_n751), .B1(new_n754), .B2(G128), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT122), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n1210), .A2(new_n1211), .B1(new_n201), .B2(new_n768), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n316), .B(new_n1212), .C1(G50), .C2(new_n758), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n771), .A2(new_n1113), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n764), .A2(G132), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1210), .A2(new_n1211), .B1(new_n777), .B2(G150), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1208), .B1(new_n1209), .B2(new_n1217), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1218), .A2(new_n787), .B1(new_n202), .B2(new_n839), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1201), .A2(new_n841), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1200), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n950), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1071), .A2(new_n1078), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1079), .A2(new_n1088), .A3(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1222), .B1(new_n1223), .B2(new_n1225), .ZN(G381));
  NOR2_X1   g1026(.A1(G375), .A2(G378), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n951), .A2(new_n973), .A3(new_n969), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1000), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1229), .A2(new_n1230), .A3(G390), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1227), .A2(new_n1228), .A3(new_n1231), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT123), .Z(G407));
  NAND2_X1  g1033(.A1(new_n1227), .A2(new_n679), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(G407), .A2(G213), .A3(new_n1234), .ZN(G409));
  INV_X1    g1035(.A(G390), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n975), .A2(new_n1236), .A3(new_n1000), .ZN(new_n1237));
  OAI21_X1  g1037(.A(G390), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  XOR2_X1   g1039(.A(G393), .B(G396), .Z(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1240), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1237), .A2(new_n1242), .A3(new_n1238), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n679), .A2(G213), .ZN(new_n1245));
  INV_X1    g1045(.A(G378), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1190), .A2(new_n1192), .A3(new_n1223), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(new_n1191), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1245), .B(new_n1249), .C1(new_n1197), .C2(new_n1246), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1225), .A2(KEYINPUT60), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1224), .A2(new_n1252), .ZN(new_n1253));
  AND4_X1   g1053(.A1(KEYINPUT125), .A2(new_n1251), .A3(new_n696), .A4(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n736), .B1(new_n1225), .B2(KEYINPUT60), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT125), .B1(new_n1255), .B2(new_n1253), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1222), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n843), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1251), .A2(new_n696), .A3(new_n1253), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT125), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1255), .A2(KEYINPUT125), .A3(new_n1253), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(G384), .A3(new_n1222), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1258), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT62), .B1(new_n1250), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1105), .A2(new_n1087), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1187), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1267), .A2(new_n1270), .A3(KEYINPUT57), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(new_n1196), .A3(new_n696), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1191), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1272), .A2(new_n1273), .B1(new_n1127), .B2(new_n1106), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(G378), .A2(new_n1191), .A3(new_n1247), .ZN(new_n1275));
  OAI21_X1  g1075(.A(KEYINPUT124), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1265), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT124), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1278), .B(new_n1249), .C1(new_n1197), .C2(new_n1246), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1276), .A2(new_n1277), .A3(new_n1279), .A4(new_n1245), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1244), .B(new_n1266), .C1(new_n1280), .C2(KEYINPUT62), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n679), .A2(G213), .A3(G2897), .ZN(new_n1284));
  AOI21_X1  g1084(.A(G384), .B1(new_n1263), .B2(new_n1222), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n843), .B(new_n1221), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1284), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1284), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1258), .A2(new_n1264), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1283), .B(KEYINPUT61), .C1(new_n1290), .C2(new_n1250), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1258), .A2(new_n1264), .A3(new_n1288), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1288), .B1(new_n1258), .B2(new_n1264), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1250), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT126), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1291), .A2(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1250), .A2(new_n1265), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1298), .B2(KEYINPUT63), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1276), .A2(new_n1279), .A3(new_n1245), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1300), .B1(new_n1301), .B2(new_n1290), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1280), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1299), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1244), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n1282), .A2(new_n1297), .B1(new_n1304), .B2(new_n1305), .ZN(G405));
  INV_X1    g1106(.A(KEYINPUT127), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1237), .A2(new_n1242), .A3(new_n1238), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1242), .B1(new_n1238), .B2(new_n1237), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1307), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1241), .A2(KEYINPUT127), .A3(new_n1243), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1277), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1310), .A2(new_n1311), .A3(new_n1265), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1227), .A2(new_n1274), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1315), .B(new_n1316), .ZN(G402));
endmodule


