//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1122, new_n1123;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n458), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT3), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n460), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n463), .A2(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NOR3_X1   g046(.A1(new_n461), .A2(new_n469), .A3(new_n471), .ZN(G160));
  INV_X1    g047(.A(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n460), .A2(G112), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  OAI22_X1  g050(.A1(new_n467), .A2(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n464), .A2(G2105), .A3(new_n466), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n476), .B1(new_n478), .B2(G124), .ZN(G162));
  NAND4_X1  g054(.A1(new_n464), .A2(G126), .A3(G2105), .A4(new_n466), .ZN(new_n480));
  OR2_X1    g055(.A1(G102), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G114), .C2(new_n460), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT4), .B1(new_n467), .B2(new_n484), .ZN(new_n485));
  XOR2_X1   g060(.A(KEYINPUT70), .B(KEYINPUT4), .Z(new_n486));
  NAND4_X1  g061(.A1(new_n486), .A2(G138), .A3(new_n460), .A4(new_n458), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n483), .B1(new_n485), .B2(new_n487), .ZN(G164));
  INV_X1    g063(.A(G543), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(KEYINPUT5), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT5), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G543), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n489), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT6), .B(G651), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  XOR2_X1   g073(.A(KEYINPUT72), .B(G88), .Z(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n498), .A2(new_n499), .B1(G50), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n495), .A2(G62), .ZN(new_n505));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  XOR2_X1   g081(.A(new_n506), .B(KEYINPUT73), .Z(new_n507));
  AOI21_X1  g082(.A(new_n504), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n503), .A2(new_n508), .ZN(G166));
  NAND2_X1  g084(.A1(new_n498), .A2(G89), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT7), .ZN(new_n511));
  NAND2_X1  g086(.A1(G76), .A2(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(new_n504), .ZN(new_n513));
  XOR2_X1   g088(.A(KEYINPUT75), .B(G51), .Z(new_n514));
  NAND2_X1  g089(.A1(new_n501), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n510), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n517));
  AOI211_X1 g092(.A(new_n517), .B(new_n490), .C1(new_n493), .C2(new_n494), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n493), .A2(new_n494), .ZN(new_n519));
  INV_X1    g094(.A(new_n490), .ZN(new_n520));
  AOI21_X1  g095(.A(KEYINPUT74), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G63), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n522), .A2(new_n523), .B1(new_n511), .B2(new_n512), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n516), .B1(new_n524), .B2(G651), .ZN(G168));
  XNOR2_X1  g100(.A(KEYINPUT78), .B(G52), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n501), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n497), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n530));
  OAI21_X1  g105(.A(G64), .B1(new_n518), .B2(new_n521), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G651), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n532), .B1(new_n531), .B2(new_n533), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n489), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n539));
  AOI21_X1  g114(.A(KEYINPUT71), .B1(new_n489), .B2(KEYINPUT5), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n520), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(new_n517), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n495), .A2(KEYINPUT74), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n538), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n533), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT76), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n546), .A2(KEYINPUT77), .A3(new_n534), .A4(G651), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n529), .B1(new_n537), .B2(new_n547), .ZN(G171));
  XOR2_X1   g123(.A(KEYINPUT79), .B(G43), .Z(new_n549));
  NAND2_X1  g124(.A1(new_n501), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n495), .A2(G81), .A3(new_n496), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g127(.A(G56), .B1(new_n518), .B2(new_n521), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n552), .B1(new_n555), .B2(G651), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n501), .A2(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n563), .B2(KEYINPUT80), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(KEYINPUT80), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n541), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(new_n498), .B2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(new_n529), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n542), .A2(new_n543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n545), .B1(new_n573), .B2(G64), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n504), .B1(new_n574), .B2(new_n532), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT77), .B1(new_n575), .B2(new_n546), .ZN(new_n576));
  INV_X1    g151(.A(new_n547), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n572), .B1(new_n576), .B2(new_n577), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  NOR3_X1   g154(.A1(new_n503), .A2(KEYINPUT81), .A3(new_n508), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n581));
  INV_X1    g156(.A(new_n508), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n581), .B1(new_n502), .B2(new_n582), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n580), .A2(new_n583), .ZN(G303));
  AOI22_X1  g159(.A1(new_n498), .A2(G87), .B1(G49), .B2(new_n501), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n573), .A2(G74), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n504), .ZN(G288));
  AOI22_X1  g162(.A1(new_n498), .A2(G86), .B1(G48), .B2(new_n501), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n495), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n504), .B2(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n573), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(new_n504), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n498), .A2(G85), .B1(G47), .B2(new_n501), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G290));
  AND3_X1   g169(.A1(new_n495), .A2(G92), .A3(new_n496), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n501), .A2(G54), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n495), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n504), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT83), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n597), .A2(new_n598), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n599), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G284));
  OAI21_X1  g183(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G860), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n605), .B1(G559), .B2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT84), .Z(G148));
  INV_X1    g191(.A(G56), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n542), .B2(new_n543), .ZN(new_n618));
  INV_X1    g193(.A(new_n554), .ZN(new_n619));
  OAI21_X1  g194(.A(G651), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n552), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n606), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n605), .A2(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g201(.A(new_n467), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n460), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n478), .A2(G123), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n628), .B1(new_n629), .B2(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n458), .A2(new_n470), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2435), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT86), .B(KEYINPUT16), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  AND3_X1   g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(G401));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT87), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2084), .B(G2090), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n659), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n662), .B1(new_n663), .B2(KEYINPUT17), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n665));
  AOI211_X1 g240(.A(new_n660), .B(new_n664), .C1(new_n663), .C2(new_n665), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n658), .A2(new_n661), .A3(new_n659), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT18), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT88), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n676), .A2(KEYINPUT89), .ZN(new_n677));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(KEYINPUT89), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n674), .A2(new_n675), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n676), .B2(new_n679), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(KEYINPUT90), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT91), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n687), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G21), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G168), .B2(new_n696), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT102), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G1966), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT103), .Z(new_n701));
  NAND2_X1  g276(.A1(G171), .A2(G16), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G5), .B2(G16), .ZN(new_n703));
  INV_X1    g278(.A(G1961), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n701), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT23), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G299), .B2(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n696), .A2(G20), .ZN(new_n710));
  MUX2_X1   g285(.A(new_n708), .B(new_n709), .S(new_n710), .Z(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G2090), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT29), .Z(new_n717));
  OAI22_X1  g292(.A1(new_n712), .A2(G1956), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G1956), .B2(new_n712), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT105), .Z(new_n720));
  AND2_X1   g295(.A1(new_n714), .A2(G26), .ZN(new_n721));
  OR2_X1    g296(.A1(G104), .A2(G2105), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n722), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT100), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n627), .A2(G140), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(KEYINPUT99), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(KEYINPUT99), .B2(new_n725), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n478), .A2(G128), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(G29), .ZN(new_n731));
  MUX2_X1   g306(.A(new_n721), .B(new_n731), .S(KEYINPUT28), .Z(new_n732));
  INV_X1    g307(.A(G2067), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G19), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n556), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT98), .B(G1341), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n734), .A2(new_n735), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n634), .A2(G29), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT104), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n627), .A2(G139), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n458), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n744));
  AOI21_X1  g319(.A(KEYINPUT25), .B1(new_n470), .B2(G103), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n470), .A2(KEYINPUT25), .A3(G103), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n743), .B1(new_n460), .B2(new_n744), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  MUX2_X1   g322(.A(G33), .B(new_n747), .S(G29), .Z(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G2072), .Z(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT31), .B(G11), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT30), .B(G28), .Z(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G29), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n714), .B1(KEYINPUT24), .B2(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(KEYINPUT24), .B2(G34), .ZN(new_n754));
  INV_X1    g329(.A(G160), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2084), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n752), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n749), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G32), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT26), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n470), .A2(G105), .ZN(new_n763));
  INV_X1    g338(.A(G141), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n762), .B(new_n763), .C1(new_n467), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n478), .B2(G129), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n760), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n756), .A2(new_n757), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT101), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n714), .A2(G27), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G164), .B2(new_n714), .ZN(new_n773));
  INV_X1    g348(.A(G2078), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n759), .A2(new_n769), .A3(new_n771), .A4(new_n775), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n742), .B(new_n776), .C1(new_n713), .C2(new_n717), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n696), .A2(G4), .ZN(new_n778));
  INV_X1    g353(.A(new_n605), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n696), .ZN(new_n780));
  INV_X1    g355(.A(G1348), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n777), .B(new_n782), .C1(G1966), .C2(new_n699), .ZN(new_n783));
  OR4_X1    g358(.A1(new_n707), .A2(new_n720), .A3(new_n740), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n714), .A2(G25), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(G95), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n788));
  INV_X1    g363(.A(G131), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n467), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n478), .B2(G119), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT93), .Z(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT94), .Z(new_n793));
  AOI21_X1  g368(.A(new_n786), .B1(new_n793), .B2(G29), .ZN(new_n794));
  MUX2_X1   g369(.A(new_n786), .B(new_n794), .S(KEYINPUT92), .Z(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT35), .B(G1991), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n696), .A2(G23), .ZN(new_n798));
  INV_X1    g373(.A(G288), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n696), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT33), .B(G1976), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT95), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n800), .B(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G6), .B(G305), .S(G16), .Z(new_n804));
  XOR2_X1   g379(.A(KEYINPUT32), .B(G1981), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n696), .A2(G22), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n696), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G1971), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(G1971), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n803), .A2(new_n806), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT34), .Z(new_n812));
  AND2_X1   g387(.A1(new_n696), .A2(G24), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G290), .B2(G16), .ZN(new_n814));
  INV_X1    g389(.A(G1986), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n814), .A2(new_n815), .B1(new_n817), .B2(KEYINPUT36), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n797), .A2(new_n812), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n817), .B1(KEYINPUT96), .B2(KEYINPUT36), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n784), .A2(new_n821), .ZN(G311));
  INV_X1    g397(.A(G311), .ZN(G150));
  NAND3_X1  g398(.A1(new_n620), .A2(KEYINPUT107), .A3(new_n621), .ZN(new_n824));
  OAI21_X1  g399(.A(G67), .B1(new_n518), .B2(new_n521), .ZN(new_n825));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n519), .A2(G93), .A3(new_n520), .A4(new_n496), .ZN(new_n828));
  INV_X1    g403(.A(G55), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n500), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT106), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n828), .B(KEYINPUT106), .C1(new_n829), .C2(new_n500), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n827), .A2(G651), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n824), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT108), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT107), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n622), .B2(new_n837), .ZN(new_n838));
  AOI211_X1 g413(.A(KEYINPUT107), .B(KEYINPUT108), .C1(new_n620), .C2(new_n621), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT108), .B1(new_n556), .B2(KEYINPUT107), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n622), .A2(new_n837), .A3(new_n836), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n841), .A2(new_n842), .A3(new_n834), .A4(new_n824), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n779), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n848));
  AOI21_X1  g423(.A(G860), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n834), .A2(new_n614), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT110), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT109), .B(KEYINPUT37), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n854), .ZN(G145));
  XNOR2_X1  g430(.A(new_n755), .B(G162), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n634), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n485), .A2(new_n487), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n480), .A2(KEYINPUT111), .A3(new_n482), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT111), .B1(new_n480), .B2(new_n482), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n857), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n729), .B(new_n792), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n766), .B(new_n637), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n863), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n627), .A2(G142), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n460), .A2(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(G130), .B2(new_n478), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n747), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G37), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n867), .B2(new_n873), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g453(.A(G290), .B(G288), .ZN(new_n879));
  XNOR2_X1  g454(.A(G166), .B(G305), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G290), .B(new_n799), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n880), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT114), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT113), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT113), .B1(new_n884), .B2(new_n882), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n886), .B1(new_n892), .B2(new_n885), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n888), .B1(new_n893), .B2(KEYINPUT114), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n611), .A2(new_n605), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n597), .B(KEYINPUT10), .ZN(new_n897));
  AOI21_X1  g472(.A(G299), .B1(new_n897), .B2(new_n603), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n895), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n896), .A2(new_n898), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(KEYINPUT112), .B(KEYINPUT41), .Z(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n899), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n844), .B(new_n624), .ZN(new_n905));
  MUX2_X1   g480(.A(new_n904), .B(new_n901), .S(new_n905), .Z(new_n906));
  XNOR2_X1  g481(.A(new_n894), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(G868), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(G868), .B2(new_n834), .ZN(G295));
  OAI21_X1  g484(.A(new_n908), .B1(G868), .B2(new_n834), .ZN(G331));
  INV_X1    g485(.A(KEYINPUT115), .ZN(new_n911));
  NAND2_X1  g486(.A1(G301), .A2(G168), .ZN(new_n912));
  NAND2_X1  g487(.A1(G171), .A2(G286), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n912), .A2(new_n843), .A3(new_n913), .A4(new_n840), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n537), .A2(new_n547), .ZN(new_n915));
  AOI21_X1  g490(.A(G286), .B1(new_n915), .B2(new_n572), .ZN(new_n916));
  AOI211_X1 g491(.A(G168), .B(new_n529), .C1(new_n537), .C2(new_n547), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n838), .A2(new_n839), .A3(new_n835), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n841), .A2(new_n842), .B1(new_n834), .B2(new_n824), .ZN(new_n919));
  OAI22_X1  g494(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n911), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n916), .A2(new_n917), .ZN(new_n922));
  INV_X1    g497(.A(new_n844), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT115), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n904), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT116), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n901), .A2(new_n914), .A3(new_n920), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT116), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n928), .B(new_n904), .C1(new_n921), .C2(new_n924), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n926), .A2(new_n891), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n844), .A2(new_n916), .A3(new_n917), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n912), .A2(new_n913), .B1(new_n843), .B2(new_n840), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT115), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n914), .A2(new_n911), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n928), .B1(new_n936), .B2(new_n904), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n929), .A2(new_n927), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n892), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n875), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n931), .B1(new_n940), .B2(KEYINPUT117), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT117), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(new_n942), .A3(new_n875), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT43), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n930), .A2(new_n875), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n900), .A2(new_n895), .ZN(new_n946));
  OAI221_X1 g521(.A(new_n946), .B1(new_n900), .B2(new_n903), .C1(new_n932), .C2(new_n933), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n921), .A2(new_n900), .A3(new_n924), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n948), .B2(KEYINPUT118), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT118), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n936), .A2(new_n950), .A3(new_n900), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n892), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n945), .A2(KEYINPUT43), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT44), .B1(new_n944), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n941), .B2(new_n943), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n952), .A2(new_n956), .A3(new_n875), .A4(new_n930), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT119), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n945), .A2(KEYINPUT119), .A3(new_n956), .A4(new_n952), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n955), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n954), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n861), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n968));
  INV_X1    g543(.A(G40), .ZN(new_n969));
  NOR4_X1   g544(.A1(new_n461), .A2(new_n469), .A3(new_n969), .A4(new_n471), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n729), .B(G2067), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1996), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n766), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n972), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n792), .B(new_n796), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n972), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n592), .A2(new_n815), .A3(new_n593), .ZN(new_n981));
  NAND2_X1  g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n971), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(KEYINPUT123), .B(G8), .Z(new_n985));
  INV_X1    g560(.A(new_n970), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  NOR2_X1   g562(.A1(G164), .A2(G1384), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n967), .B2(new_n987), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(G2090), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n970), .B1(new_n988), .B2(KEYINPUT45), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT120), .B1(new_n966), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT120), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n861), .A2(new_n995), .A3(KEYINPUT45), .A4(new_n965), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n992), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(G1971), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n985), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(G8), .B1(new_n580), .B2(new_n583), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT55), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n966), .A2(new_n986), .ZN(new_n1003));
  INV_X1    g578(.A(new_n985), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(new_n1006), .B2(G288), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n799), .A2(G1976), .ZN(new_n1008));
  OR3_X1    g583(.A1(new_n1007), .A2(KEYINPUT52), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(G305), .B(G1981), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT49), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n1005), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(KEYINPUT52), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1009), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n861), .A2(new_n987), .A3(new_n965), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1016), .A2(new_n713), .A3(new_n970), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n997), .B2(G1971), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1015), .B1(new_n1019), .B2(KEYINPUT121), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1001), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT121), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1022), .B(new_n1018), .C1(new_n997), .C2(G1971), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT122), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT122), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1020), .A2(new_n1021), .A3(new_n1026), .A4(new_n1023), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1014), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1016), .A2(new_n970), .A3(new_n1017), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G2084), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n988), .A2(KEYINPUT45), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n970), .B(new_n1031), .C1(new_n967), .C2(KEYINPUT45), .ZN(new_n1032));
  INV_X1    g607(.A(G1966), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1030), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(G168), .A2(new_n1004), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1034), .A2(new_n1004), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1036), .B1(new_n1034), .B2(new_n1015), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT51), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1037), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(G171), .B(KEYINPUT54), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT53), .B1(new_n997), .B2(new_n774), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n704), .B2(new_n1029), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n774), .A2(KEYINPUT53), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n968), .A2(new_n986), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1031), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1044), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n994), .A2(new_n996), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1046), .A2(new_n1044), .A3(new_n1052), .ZN(new_n1053));
  OR3_X1    g628(.A1(new_n1043), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  XOR2_X1   g629(.A(G299), .B(KEYINPUT57), .Z(new_n1055));
  INV_X1    g630(.A(G1956), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT56), .B(G2072), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1056), .A2(new_n990), .B1(new_n997), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1059), .A2(KEYINPUT126), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1060), .A2(KEYINPUT61), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1029), .A2(new_n781), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1003), .A2(new_n733), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n779), .B1(new_n1065), .B2(KEYINPUT60), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(KEYINPUT60), .ZN(new_n1067));
  MUX2_X1   g642(.A(new_n779), .B(new_n1066), .S(new_n1067), .Z(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT58), .B(G1341), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1003), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n997), .B2(new_n975), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(new_n622), .ZN(new_n1072));
  XOR2_X1   g647(.A(new_n1072), .B(KEYINPUT59), .Z(new_n1073));
  NAND2_X1  g648(.A1(new_n1059), .A2(KEYINPUT61), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1061), .A2(new_n1068), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1065), .A2(new_n605), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n1059), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1054), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n1081));
  OAI211_X1 g656(.A(G171), .B(new_n1080), .C1(new_n1043), .C2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n1081), .B2(new_n1043), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1002), .B(new_n1028), .C1(new_n1079), .C2(new_n1083), .ZN(new_n1084));
  AOI211_X1 g659(.A(G1976), .B(G288), .C1(new_n1011), .C2(new_n1005), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G305), .A2(G1981), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1005), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n1014), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1014), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1038), .A2(G286), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1088), .A2(new_n1002), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT63), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1028), .A2(KEYINPUT124), .A3(new_n1002), .A4(new_n1091), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1001), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1028), .A2(KEYINPUT63), .A3(new_n1091), .A4(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1089), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1084), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g678(.A(KEYINPUT125), .B(new_n1089), .C1(new_n1097), .C2(new_n1100), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n984), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n971), .B1(new_n973), .B2(new_n766), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT46), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n972), .A2(new_n975), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT47), .Z(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n971), .B2(new_n981), .ZN(new_n1113));
  OR3_X1    g688(.A1(new_n971), .A2(new_n981), .A3(new_n1112), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n977), .A2(new_n979), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n793), .A2(new_n796), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n977), .A2(new_n1116), .B1(new_n733), .B2(new_n729), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1117), .B2(new_n971), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1111), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1105), .A2(new_n1119), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g695(.A1(new_n694), .A2(G319), .A3(new_n671), .ZN(new_n1122));
  NOR3_X1   g696(.A1(new_n877), .A2(G401), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g697(.A(new_n1123), .B1(new_n957), .B2(new_n962), .ZN(G225));
  INV_X1    g698(.A(G225), .ZN(G308));
endmodule


