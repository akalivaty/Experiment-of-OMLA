//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  XNOR2_X1  g0004(.A(KEYINPUT64), .B(G20), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G1), .A2(G13), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n202), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT65), .Z(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n211), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n210), .B(new_n214), .C1(new_n221), .C2(KEYINPUT1), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0023(.A(G226), .B(G232), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT67), .ZN(new_n225));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  INV_X1    g0040(.A(G33), .ZN(new_n241));
  INV_X1    g0041(.A(G41), .ZN(new_n242));
  OAI211_X1 g0042(.A(G1), .B(G13), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G45), .ZN(new_n244));
  AOI21_X1  g0044(.A(G1), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n243), .A2(G274), .A3(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n247), .B1(G238), .B2(new_n251), .ZN(new_n252));
  OR2_X1    g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G226), .ZN(new_n258));
  INV_X1    g0058(.A(G97), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n257), .A2(new_n258), .B1(new_n241), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT75), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n255), .A2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G232), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n256), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(KEYINPUT75), .A3(G232), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n260), .B1(new_n264), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n252), .B1(new_n270), .B2(new_n243), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT13), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT13), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n273), .B(new_n252), .C1(new_n270), .C2(new_n243), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(KEYINPUT76), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT76), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n271), .A2(new_n276), .A3(KEYINPUT13), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G169), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT14), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT14), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n275), .A2(new_n280), .A3(G169), .A4(new_n277), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n272), .A2(G179), .A3(new_n274), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT77), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OR2_X1    g0084(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n279), .A2(new_n281), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G68), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT64), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT64), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n241), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G77), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n206), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT69), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT69), .B1(new_n299), .B2(new_n206), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(KEYINPUT11), .ZN(new_n307));
  INV_X1    g0107(.A(G13), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(G1), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G20), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n288), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT12), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n306), .A2(KEYINPUT11), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n310), .B1(new_n302), .B2(new_n303), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n248), .A2(G20), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G68), .A3(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n307), .A2(new_n313), .A3(new_n314), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n286), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n274), .A2(G190), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n319), .B1(new_n321), .B2(new_n272), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n275), .A2(G200), .A3(new_n277), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n326));
  INV_X1    g0126(.A(G150), .ZN(new_n327));
  INV_X1    g0127(.A(new_n287), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT70), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G58), .ZN(new_n330));
  XOR2_X1   g0130(.A(new_n330), .B(KEYINPUT8), .Z(new_n331));
  OAI221_X1 g0131(.A(new_n326), .B1(new_n327), .B2(new_n328), .C1(new_n331), .C2(new_n296), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n304), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n317), .A2(G50), .ZN(new_n334));
  XOR2_X1   g0134(.A(new_n334), .B(KEYINPUT71), .Z(new_n335));
  OAI221_X1 g0135(.A(new_n333), .B1(G50), .B2(new_n310), .C1(new_n315), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT9), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n246), .B1(new_n250), .B2(new_n258), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n267), .A2(G1698), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(G222), .B1(G77), .B2(new_n267), .ZN(new_n340));
  XOR2_X1   g0140(.A(KEYINPUT68), .B(G223), .Z(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n262), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n206), .B1(G33), .B2(G41), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n338), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n336), .A2(new_n337), .B1(new_n344), .B2(G190), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  OAI221_X1 g0146(.A(new_n345), .B1(new_n337), .B2(new_n336), .C1(new_n346), .C2(new_n344), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT10), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n336), .B1(new_n344), .B2(G169), .ZN(new_n349));
  INV_X1    g0149(.A(G179), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n344), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n331), .A2(new_n311), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n330), .B(KEYINPUT8), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n317), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n354), .B1(new_n356), .B2(new_n315), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT79), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n354), .B(KEYINPUT79), .C1(new_n315), .C2(new_n356), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n302), .A2(new_n303), .ZN(new_n362));
  INV_X1    g0162(.A(G58), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n288), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n364), .A2(new_n201), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(G20), .B1(G159), .B2(new_n287), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n253), .A2(new_n291), .A3(new_n293), .A4(new_n254), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT78), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT78), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n372), .A3(new_n369), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n290), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n367), .B1(new_n375), .B2(G68), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n362), .B1(new_n376), .B2(KEYINPUT16), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n368), .A2(KEYINPUT7), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n267), .A2(new_n369), .A3(new_n290), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n366), .B1(new_n380), .B2(new_n288), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n361), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n246), .B1(new_n250), .B2(new_n263), .ZN(new_n385));
  INV_X1    g0185(.A(G223), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n256), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n258), .A2(G1698), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n387), .B(new_n388), .C1(new_n265), .C2(new_n266), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n243), .B1(new_n391), .B2(KEYINPUT80), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT80), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n393), .A3(new_n390), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n385), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n395), .A2(G190), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n346), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n384), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n359), .A2(new_n360), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n267), .B2(new_n205), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n374), .B1(new_n403), .B2(new_n372), .ZN(new_n404));
  INV_X1    g0204(.A(new_n373), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(KEYINPUT16), .A3(new_n366), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n304), .A3(new_n383), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n398), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT17), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n401), .A2(new_n410), .ZN(new_n411));
  AOI211_X1 g0211(.A(G179), .B(new_n385), .C1(new_n392), .C2(new_n394), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n391), .A2(KEYINPUT80), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(new_n343), .A3(new_n394), .ZN(new_n414));
  INV_X1    g0214(.A(new_n385), .ZN(new_n415));
  AOI21_X1  g0215(.A(G169), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT81), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n350), .A3(new_n415), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT81), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n418), .B(new_n419), .C1(G169), .C2(new_n395), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n384), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT18), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n384), .B2(new_n421), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n411), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT15), .B(G87), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT73), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n295), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n430), .A2(KEYINPUT74), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT8), .B(G58), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n297), .A2(new_n205), .B1(new_n432), .B2(new_n328), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n430), .B2(KEYINPUT74), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n362), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n316), .A2(G77), .A3(new_n317), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(G77), .B2(new_n310), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n247), .B1(G244), .B2(new_n251), .ZN(new_n440));
  INV_X1    g0240(.A(G238), .ZN(new_n441));
  INV_X1    g0241(.A(G107), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n262), .A2(new_n441), .B1(new_n442), .B2(new_n255), .ZN(new_n443));
  OR3_X1    g0243(.A1(new_n257), .A2(KEYINPUT72), .A3(new_n263), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT72), .B1(new_n257), .B2(new_n263), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n440), .B1(new_n446), .B2(new_n243), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n447), .A2(G179), .ZN(new_n448));
  INV_X1    g0248(.A(G169), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n439), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(G200), .ZN(new_n452));
  INV_X1    g0252(.A(G190), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n438), .B(new_n452), .C1(new_n453), .C2(new_n447), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n325), .A2(new_n353), .A3(new_n427), .A4(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n339), .A2(KEYINPUT4), .A3(G244), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n255), .A2(G244), .A3(new_n256), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT4), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n268), .A2(G250), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n457), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n343), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n248), .B(G45), .C1(new_n242), .C2(KEYINPUT5), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G274), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n343), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n465), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n343), .B1(new_n472), .B2(new_n470), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G257), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n464), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n449), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n442), .A2(KEYINPUT6), .A3(G97), .ZN(new_n477));
  XOR2_X1   g0277(.A(G97), .B(G107), .Z(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(KEYINPUT6), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n479), .A2(new_n294), .B1(G77), .B2(new_n287), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n442), .B2(new_n380), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n304), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n248), .A2(G33), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n362), .A2(new_n310), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G97), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n310), .A2(G97), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n482), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n463), .A2(new_n343), .B1(G257), .B2(new_n473), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n350), .A3(new_n471), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n476), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT83), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n482), .A2(new_n486), .A3(new_n488), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n475), .A2(G200), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n496), .C1(new_n453), .C2(new_n475), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n476), .A2(new_n489), .A3(KEYINPUT83), .A4(new_n491), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G250), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n244), .B2(G1), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n248), .A2(new_n468), .A3(G45), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n243), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT84), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n257), .B2(new_n441), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n339), .A2(KEYINPUT84), .A3(G238), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G244), .ZN(new_n509));
  INV_X1    g0309(.A(G116), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n262), .A2(new_n509), .B1(new_n241), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n504), .B1(new_n513), .B2(new_n343), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n350), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n506), .B2(new_n507), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n503), .B1(new_n516), .B2(new_n243), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n449), .ZN(new_n518));
  NOR3_X1   g0318(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n519), .B(KEYINPUT85), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n241), .A2(new_n259), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n294), .B1(KEYINPUT19), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n255), .A2(new_n205), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n520), .A2(new_n522), .B1(new_n288), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT19), .B1(new_n295), .B2(G97), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n304), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n429), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n311), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n528), .C1(new_n527), .C2(new_n484), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n515), .A2(new_n518), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n514), .A2(G190), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n517), .A2(G200), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n526), .A2(new_n528), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n485), .A2(G87), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  XNOR2_X1  g0335(.A(KEYINPUT88), .B(KEYINPUT22), .ZN(new_n536));
  INV_X1    g0336(.A(G87), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n523), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT22), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(KEYINPUT88), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n255), .A2(new_n205), .A3(G87), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT89), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n294), .A2(new_n543), .A3(new_n544), .A4(new_n442), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n442), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT89), .B1(new_n205), .B2(new_n546), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n241), .A2(new_n510), .A3(G20), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(G20), .B2(new_n442), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  OR3_X1    g0351(.A1(new_n542), .A2(KEYINPUT24), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT24), .B1(new_n542), .B2(new_n551), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n304), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n484), .A2(new_n442), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n309), .A2(G20), .A3(new_n442), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n557), .B(KEYINPUT25), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n473), .A2(G264), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n471), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n268), .A2(G257), .B1(G33), .B2(G294), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n339), .A2(G250), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n243), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(G200), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n564), .ZN(new_n567));
  INV_X1    g0367(.A(G257), .ZN(new_n568));
  INV_X1    g0368(.A(G294), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n262), .A2(new_n568), .B1(new_n241), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n343), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n471), .A3(new_n561), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n566), .B1(new_n572), .B2(new_n453), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n530), .B(new_n535), .C1(new_n560), .C2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n499), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT87), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(KEYINPUT21), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT86), .B1(new_n257), .B2(new_n568), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT86), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n339), .A2(new_n579), .A3(G257), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(G264), .ZN(new_n582));
  INV_X1    g0382(.A(G303), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n262), .A2(new_n582), .B1(new_n583), .B2(new_n255), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n243), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n473), .A2(G270), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n471), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(G169), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n484), .A2(new_n510), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n311), .A2(new_n510), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n205), .B(new_n462), .C1(G33), .C2(new_n259), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n299), .A2(new_n206), .B1(G20), .B2(new_n510), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT20), .B1(new_n592), .B2(new_n593), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n577), .B1(new_n589), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n471), .A2(new_n587), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n584), .B1(new_n580), .B2(new_n578), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n243), .B2(new_n600), .ZN(new_n601));
  OAI221_X1 g0401(.A(new_n591), .B1(new_n594), .B2(new_n595), .C1(new_n484), .C2(new_n510), .ZN(new_n602));
  INV_X1    g0402(.A(new_n577), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(G169), .A4(new_n603), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n586), .A2(new_n588), .A3(new_n350), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n602), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n598), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n449), .B1(new_n562), .B2(new_n565), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n572), .B2(G179), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n555), .B2(new_n559), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n586), .A2(new_n588), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n597), .B1(new_n611), .B2(new_n346), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n601), .A2(new_n453), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n607), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n456), .A2(new_n575), .A3(new_n615), .ZN(G372));
  AND2_X1   g0416(.A1(new_n494), .A2(new_n498), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n535), .A2(new_n530), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT26), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n618), .A2(new_n492), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n530), .C1(KEYINPUT26), .C2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n575), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n607), .A2(new_n610), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n456), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT90), .B1(new_n384), .B2(new_n421), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n408), .A2(new_n402), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(new_n417), .A4(new_n420), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n424), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n627), .A2(new_n630), .A3(KEYINPUT18), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n451), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n286), .A2(new_n319), .B1(new_n324), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n401), .A2(new_n410), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n351), .B1(new_n638), .B2(new_n348), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n626), .A2(new_n639), .ZN(G369));
  AOI21_X1  g0440(.A(new_n362), .B1(new_n552), .B2(new_n553), .ZN(new_n641));
  INV_X1    g0441(.A(new_n559), .ZN(new_n642));
  OAI221_X1 g0442(.A(new_n608), .B1(G179), .B2(new_n572), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n573), .A2(new_n641), .A3(new_n642), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n205), .A2(new_n309), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n646), .A2(G213), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G343), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n555), .B2(new_n559), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n643), .B1(new_n644), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n610), .A2(new_n649), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT91), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n649), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n602), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n607), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n614), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n607), .A2(new_n649), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n655), .A2(new_n656), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(new_n652), .A3(new_n665), .ZN(G399));
  INV_X1    g0466(.A(new_n212), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G41), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n248), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n520), .A2(new_n510), .ZN(new_n671));
  INV_X1    g0471(.A(new_n668), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n670), .A2(new_n671), .B1(new_n208), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  INV_X1    g0474(.A(G330), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT30), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n562), .A2(new_n565), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n514), .A2(new_n490), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n611), .A2(G179), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n517), .A2(new_n572), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(KEYINPUT30), .A3(new_n605), .A4(new_n490), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n677), .A2(G179), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n475), .A3(new_n517), .A4(new_n601), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT31), .B1(new_n685), .B2(new_n658), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(KEYINPUT92), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n685), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n687), .B(new_n688), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n618), .A2(new_n644), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n690), .A2(new_n615), .A3(new_n691), .A4(new_n649), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT93), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT93), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n575), .A2(new_n694), .A3(new_n615), .A4(new_n649), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n675), .B1(new_n689), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n649), .B1(new_n622), .B2(new_n625), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n624), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n701), .A2(KEYINPUT94), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(KEYINPUT94), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n702), .A2(new_n623), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n530), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n621), .B2(KEYINPUT26), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n619), .B2(KEYINPUT26), .ZN(new_n707));
  OAI211_X1 g0507(.A(KEYINPUT29), .B(new_n649), .C1(new_n704), .C2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n697), .B1(new_n700), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n674), .B1(new_n709), .B2(G1), .ZN(G364));
  NOR3_X1   g0510(.A1(new_n294), .A2(new_n308), .A3(new_n244), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT95), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n670), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n662), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n661), .A2(G330), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G13), .A2(G33), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G20), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n660), .B2(new_n614), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n667), .A2(new_n267), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G355), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G116), .B2(new_n212), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n236), .A2(new_n244), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n667), .A2(new_n255), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n244), .B2(new_n209), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n724), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n206), .B1(G20), .B2(new_n449), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n720), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n713), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G190), .A2(G200), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n294), .A2(new_n350), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT97), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(KEYINPUT97), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G329), .ZN(new_n741));
  INV_X1    g0541(.A(G326), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n205), .A2(new_n350), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n744), .A2(new_n453), .A3(new_n346), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n744), .A2(G190), .A3(new_n346), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT33), .B(G317), .Z(new_n749));
  OAI221_X1 g0549(.A(new_n741), .B1(new_n742), .B2(new_n746), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  NOR4_X1   g0550(.A1(new_n290), .A2(new_n453), .A3(new_n346), .A4(G179), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n255), .B1(new_n751), .B2(G303), .ZN(new_n752));
  INV_X1    g0552(.A(G283), .ZN(new_n753));
  NOR4_X1   g0553(.A1(new_n205), .A2(G179), .A3(G190), .A4(new_n346), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n453), .A2(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n744), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G322), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n752), .B1(new_n753), .B2(new_n755), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n743), .A2(new_n734), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n294), .B1(new_n757), .B2(G179), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n762), .A2(new_n763), .B1(new_n765), .B2(new_n569), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n750), .A2(new_n761), .A3(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT98), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n754), .A2(G107), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n267), .B1(new_n751), .B2(G87), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n770), .B(new_n771), .C1(new_n759), .C2(new_n363), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(G50), .B2(new_n745), .ZN(new_n773));
  INV_X1    g0573(.A(new_n762), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n774), .A2(G77), .B1(G97), .B2(new_n764), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT96), .B(G159), .Z(new_n776));
  NAND2_X1  g0576(.A1(new_n736), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT32), .Z(new_n778));
  NAND2_X1  g0578(.A1(new_n747), .A2(G68), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n773), .A2(new_n775), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n768), .A2(KEYINPUT98), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n769), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n733), .B1(new_n782), .B2(new_n730), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n717), .B1(new_n721), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(G396));
  OAI21_X1  g0585(.A(KEYINPUT101), .B1(new_n451), .B2(new_n649), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n438), .B1(new_n449), .B2(new_n447), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT101), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n787), .A2(new_n788), .A3(new_n448), .A4(new_n658), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n451), .A2(KEYINPUT100), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT100), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n439), .A2(new_n792), .A3(new_n448), .A4(new_n450), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n439), .A2(new_n658), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n791), .A2(new_n454), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n698), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT102), .ZN(new_n798));
  INV_X1    g0598(.A(new_n796), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n649), .B(new_n799), .C1(new_n622), .C2(new_n625), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n697), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n698), .A2(KEYINPUT102), .A3(new_n796), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n804), .A2(KEYINPUT103), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n802), .B1(new_n801), .B2(new_n803), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n805), .A2(new_n713), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(KEYINPUT103), .B2(new_n804), .ZN(new_n808));
  INV_X1    g0608(.A(new_n730), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n719), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n713), .B1(G77), .B2(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G143), .A2(new_n758), .B1(new_n774), .B2(new_n776), .ZN(new_n812));
  INV_X1    g0612(.A(G137), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n748), .B2(new_n327), .C1(new_n813), .C2(new_n746), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT34), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n765), .A2(new_n363), .ZN(new_n818));
  INV_X1    g0618(.A(G50), .ZN(new_n819));
  INV_X1    g0619(.A(new_n751), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n255), .B1(new_n819), .B2(new_n820), .C1(new_n755), .C2(new_n288), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n818), .B(new_n821), .C1(new_n740), .C2(G132), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n816), .A2(new_n817), .A3(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n758), .A2(G294), .B1(G97), .B2(new_n764), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT99), .Z(new_n825));
  AOI21_X1  g0625(.A(new_n255), .B1(new_n751), .B2(G107), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n826), .B1(new_n762), .B2(new_n510), .C1(new_n755), .C2(new_n537), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n740), .B2(G311), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G283), .A2(new_n747), .B1(new_n745), .B2(G303), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n825), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n823), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n811), .B1(new_n831), .B2(new_n730), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n799), .B2(new_n719), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n808), .A2(new_n833), .ZN(G384));
  OR2_X1    g0634(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n835), .A2(G116), .A3(new_n207), .A4(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT36), .Z(new_n838));
  OR3_X1    g0638(.A1(new_n208), .A2(new_n297), .A3(new_n364), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n819), .A2(G68), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n248), .B(G13), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  INV_X1    g0643(.A(new_n648), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n384), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(new_n422), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n409), .A2(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n631), .A2(new_n399), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT105), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n409), .B1(new_n627), .B2(new_n630), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT105), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n845), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n849), .B1(new_n855), .B2(KEYINPUT37), .ZN(new_n856));
  INV_X1    g0656(.A(new_n845), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n634), .B2(new_n411), .ZN(new_n858));
  OAI211_X1 g0658(.A(KEYINPUT106), .B(new_n843), .C1(new_n856), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n406), .A2(new_n366), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n382), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n361), .B1(new_n377), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n399), .B1(new_n421), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n844), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n848), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n637), .B1(new_n425), .B2(new_n423), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n377), .A2(new_n861), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n648), .B1(new_n868), .B2(new_n361), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n866), .B(KEYINPUT38), .C1(new_n867), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n859), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n858), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n851), .B2(new_n854), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n874), .B2(new_n849), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT106), .B1(new_n875), .B2(new_n843), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT110), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT106), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n858), .B1(new_n879), .B2(new_n848), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n878), .B1(new_n880), .B2(KEYINPUT38), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT110), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n881), .A2(new_n882), .A3(new_n870), .A4(new_n859), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT108), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n686), .B1(new_n884), .B2(new_n688), .ZN(new_n885));
  AOI211_X1 g0685(.A(KEYINPUT108), .B(KEYINPUT31), .C1(new_n685), .C2(new_n658), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n696), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n319), .A2(new_n658), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n320), .A2(new_n324), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n324), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n319), .B(new_n658), .C1(new_n891), .C2(new_n286), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n796), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n888), .A2(KEYINPUT40), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n877), .A2(new_n883), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n869), .B1(new_n411), .B2(new_n426), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n869), .B(new_n399), .C1(new_n421), .C2(new_n862), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n898), .A2(KEYINPUT37), .B1(new_n846), .B2(new_n847), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n843), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n870), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n888), .A3(new_n893), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT109), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n904), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT109), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n896), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n456), .A2(new_n888), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n675), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n700), .A2(new_n456), .A3(new_n708), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n639), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT107), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n901), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n881), .A2(new_n870), .A3(new_n859), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n917), .B2(new_n915), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n320), .A2(new_n658), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT104), .Z(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n634), .A2(new_n648), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n791), .A2(new_n793), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n649), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n800), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n890), .A2(new_n892), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n922), .B1(new_n927), .B2(new_n901), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n914), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n911), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(G1), .B1(new_n294), .B2(new_n308), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n911), .A2(new_n930), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n842), .B1(new_n933), .B2(new_n934), .ZN(G367));
  NAND2_X1  g0735(.A1(new_n489), .A2(new_n658), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n690), .A2(KEYINPUT111), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n492), .B2(new_n649), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT111), .B1(new_n690), .B2(new_n936), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n665), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT112), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n610), .B1(new_n938), .B2(new_n939), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n658), .B1(new_n945), .B2(new_n617), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n942), .B2(KEYINPUT42), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n533), .A2(new_n534), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n705), .A2(new_n948), .A3(new_n658), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n658), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(new_n535), .A3(new_n530), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n944), .A2(new_n947), .B1(KEYINPUT43), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n952), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n663), .A2(new_n940), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n944), .A2(new_n955), .A3(new_n954), .A4(new_n947), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n958), .B1(new_n957), .B2(new_n959), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n668), .B(KEYINPUT41), .Z(new_n963));
  NAND2_X1  g0763(.A1(new_n665), .A2(new_n652), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(new_n940), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT113), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(KEYINPUT113), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n966), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n964), .A2(new_n940), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT44), .Z(new_n973));
  NAND3_X1  g0773(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n663), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n657), .B(new_n662), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(new_n664), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n970), .A2(new_n973), .A3(new_n971), .A4(new_n663), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n976), .A2(new_n709), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n963), .B1(new_n980), .B2(new_n709), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n712), .A2(new_n248), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n962), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT46), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n820), .B2(new_n510), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n751), .A2(KEYINPUT46), .A3(G116), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(new_n755), .C2(new_n259), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G311), .B2(new_n745), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n569), .B2(new_n748), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n255), .B1(new_n736), .B2(G317), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n759), .B2(new_n583), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n762), .A2(new_n753), .B1(new_n765), .B2(new_n442), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n745), .A2(G143), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n736), .A2(G137), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n754), .A2(G77), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n267), .B1(new_n751), .B2(G58), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n764), .A2(G68), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n819), .B2(new_n762), .C1(new_n759), .C2(new_n327), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n999), .B(new_n1001), .C1(new_n747), .C2(new_n776), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n994), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT47), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n730), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n954), .A2(new_n720), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n732), .B1(new_n232), .B2(new_n726), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n212), .B2(new_n527), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1005), .A2(new_n713), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n984), .A2(new_n1009), .ZN(G387));
  NOR2_X1   g0810(.A1(new_n978), .A2(new_n709), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT115), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n978), .A2(new_n709), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(KEYINPUT115), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1012), .A2(new_n668), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n727), .B1(new_n229), .B2(G45), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n671), .B2(new_n722), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n432), .A2(G50), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT50), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n244), .B1(new_n288), .B2(new_n297), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n671), .B(new_n1020), .C1(new_n1019), .C2(new_n1018), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1017), .A2(new_n1021), .B1(G107), .B2(new_n212), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n714), .B1(new_n1022), .B2(new_n731), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n429), .A2(new_n764), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n288), .B2(new_n762), .C1(new_n759), .C2(new_n819), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n820), .A2(new_n297), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n267), .B(new_n1026), .C1(new_n754), .C2(G97), .ZN(new_n1027));
  INV_X1    g0827(.A(G159), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1027), .B1(new_n327), .B2(new_n735), .C1(new_n1028), .C2(new_n746), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1025), .B(new_n1029), .C1(new_n355), .C2(new_n747), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n764), .A2(G283), .B1(new_n751), .B2(G294), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G317), .A2(new_n758), .B1(new_n774), .B2(G303), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n748), .B2(new_n763), .C1(new_n760), .C2(new_n746), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT114), .Z(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1031), .B1(new_n1035), .B2(KEYINPUT48), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(KEYINPUT48), .B2(new_n1035), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT49), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n267), .B1(new_n742), .B2(new_n735), .C1(new_n755), .C2(new_n510), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n1037), .B2(KEYINPUT49), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1030), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1023), .B1(new_n1041), .B2(new_n809), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n657), .B2(new_n720), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n978), .B2(new_n983), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1015), .A2(new_n1044), .ZN(G393));
  NAND2_X1  g0845(.A1(new_n976), .A2(new_n979), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n1013), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1047), .A2(new_n668), .A3(new_n980), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n762), .A2(new_n432), .B1(new_n765), .B2(new_n297), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n255), .B1(new_n288), .B2(new_n820), .C1(new_n755), .C2(new_n537), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G143), .C2(new_n736), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n746), .A2(new_n327), .B1(new_n759), .B2(new_n1028), .ZN(new_n1052));
  XOR2_X1   g0852(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1051), .B(new_n1054), .C1(new_n819), .C2(new_n748), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n745), .A2(G317), .B1(new_n758), .B2(G311), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n770), .B(new_n267), .C1(new_n753), .C2(new_n820), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G322), .B2(new_n736), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n774), .A2(G294), .B1(G116), .B2(new_n764), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n583), .C2(new_n748), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1055), .A2(new_n1056), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n730), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n239), .A2(new_n726), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1065), .B(new_n731), .C1(new_n259), .C2(new_n212), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n713), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n940), .B2(new_n720), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1046), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n983), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1048), .A2(new_n1070), .ZN(G390));
  OAI211_X1 g0871(.A(new_n649), .B(new_n799), .C1(new_n704), .C2(new_n707), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n924), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n920), .B1(new_n1073), .B2(new_n926), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n877), .A2(new_n883), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1075), .B1(new_n918), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n675), .B1(new_n696), .B2(new_n887), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1078), .A2(new_n893), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n697), .A2(new_n799), .A3(new_n926), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1075), .B(new_n1081), .C1(new_n918), .C2(new_n1076), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n456), .A2(new_n1078), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n912), .A2(new_n639), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n926), .B1(new_n697), .B2(new_n799), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n925), .B1(new_n1087), .B2(new_n1079), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1073), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1078), .A2(new_n799), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1081), .B(new_n1089), .C1(new_n926), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n672), .B1(new_n1083), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1093), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1080), .A2(new_n1082), .A3(new_n1095), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n713), .B1(new_n355), .B2(new_n810), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n740), .A2(G125), .B1(G137), .B2(new_n747), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n745), .A2(G128), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n267), .B1(new_n754), .B2(G50), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n751), .A2(G150), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT53), .Z(new_n1103));
  NAND4_X1  g0903(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT54), .B(G143), .Z(new_n1105));
  NAND2_X1  g0905(.A1(new_n774), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(G132), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1106), .B1(new_n1028), .B2(new_n765), .C1(new_n759), .C2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G116), .A2(new_n758), .B1(new_n774), .B2(G97), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n267), .B1(new_n820), .B2(new_n537), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G68), .B2(new_n754), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(new_n297), .C2(new_n765), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G107), .A2(new_n747), .B1(new_n745), .B2(G283), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n569), .B2(new_n739), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1104), .A2(new_n1108), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1098), .B1(new_n1115), .B2(new_n730), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n918), .B2(new_n719), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n1083), .B2(new_n982), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1097), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(G378));
  INV_X1    g0920(.A(new_n929), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n675), .B1(new_n907), .B2(new_n905), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n895), .A2(new_n1122), .A3(KEYINPUT117), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT117), .B1(new_n895), .B2(new_n1122), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n336), .A2(new_n648), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n353), .B(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1123), .A2(new_n1124), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1129), .A2(new_n895), .A3(new_n1122), .A4(KEYINPUT117), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1121), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n895), .A2(new_n1122), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT117), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n895), .A2(new_n1122), .A3(KEYINPUT117), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n1137), .A3(new_n1128), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n929), .A3(new_n1131), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1133), .A2(KEYINPUT118), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1096), .A2(new_n1086), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT118), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1138), .A2(new_n1142), .A3(new_n929), .A4(new_n1131), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT57), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1096), .B2(new_n1086), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1138), .A2(new_n929), .A3(new_n1131), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n929), .B1(new_n1138), .B2(new_n1131), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n668), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1140), .A2(new_n983), .A3(new_n1143), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1129), .A2(new_n718), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n713), .B1(G50), .B2(new_n810), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G97), .A2(new_n747), .B1(new_n745), .B2(G116), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n753), .B2(new_n739), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1026), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n754), .A2(G58), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n255), .A2(G41), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1159), .A2(new_n1000), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n759), .A2(new_n442), .B1(new_n527), .B2(new_n762), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1158), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT58), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G125), .A2(new_n745), .B1(new_n747), .B2(G132), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n764), .A2(G150), .B1(new_n751), .B2(new_n1105), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G128), .A2(new_n758), .B1(new_n774), .B2(G137), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n736), .A2(G124), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G33), .B(G41), .C1(new_n754), .C2(new_n776), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1164), .A2(KEYINPUT58), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1161), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1176), .B(new_n819), .C1(G33), .C2(G41), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1165), .A2(new_n1174), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1156), .B1(new_n1178), .B2(new_n730), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1155), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1154), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1153), .A2(new_n1182), .ZN(G375));
  INV_X1    g0983(.A(new_n963), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1085), .A2(new_n1088), .A3(new_n1091), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1093), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n890), .A2(new_n718), .A3(new_n892), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n713), .B1(G68), .B2(new_n810), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT119), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n745), .A2(G294), .B1(G107), .B2(new_n774), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n510), .B2(new_n748), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT120), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n255), .B1(new_n751), .B2(G97), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1024), .A2(new_n997), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G283), .B2(new_n758), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1192), .B(new_n1195), .C1(new_n583), .C2(new_n739), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n774), .A2(G150), .B1(G159), .B2(new_n751), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n819), .B2(new_n765), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1160), .A2(new_n255), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT121), .Z(new_n1200));
  AOI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(G128), .C2(new_n740), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT122), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n747), .A2(new_n1105), .B1(new_n758), .B2(G137), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1107), .B2(new_n746), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1196), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1189), .B1(new_n1205), .B2(new_n730), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1092), .A2(new_n983), .B1(new_n1187), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1186), .A2(new_n1207), .ZN(G381));
  NOR2_X1   g1008(.A1(G393), .A2(G396), .ZN(new_n1209));
  INV_X1    g1009(.A(G384), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OR3_X1    g1011(.A1(G390), .A2(G381), .A3(new_n1211), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(G375), .A2(new_n1212), .A3(G387), .A4(G378), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT123), .ZN(G407));
  INV_X1    g1014(.A(G343), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(G213), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT124), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1153), .A2(new_n1182), .A3(new_n1119), .A4(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT125), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(G407), .A2(G213), .A3(new_n1219), .ZN(G409));
  NAND3_X1  g1020(.A1(new_n984), .A2(G390), .A3(new_n1009), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(KEYINPUT127), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(G393), .B(new_n784), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(G390), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G387), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1221), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1222), .A2(new_n1226), .A3(new_n1221), .A4(new_n1223), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1093), .A2(KEYINPUT60), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(new_n1185), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(new_n672), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1185), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1207), .ZN(new_n1236));
  OR3_X1    g1036(.A1(new_n1235), .A2(new_n1210), .A3(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1210), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(KEYINPUT62), .A3(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1153), .A2(G378), .A3(new_n1182), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n982), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1155), .B2(new_n1179), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1140), .A2(new_n1184), .A3(new_n1141), .A4(new_n1143), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1119), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1217), .B(new_n1239), .C1(new_n1240), .C2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1151), .B1(new_n1145), .B2(new_n1144), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1247), .A2(new_n1119), .A3(new_n1181), .ZN(new_n1248));
  AOI21_X1  g1048(.A(G378), .B1(new_n1243), .B2(new_n1242), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT126), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT126), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1240), .A2(new_n1245), .A3(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1216), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT62), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1246), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1217), .B1(new_n1240), .B2(new_n1245), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1237), .A2(new_n1238), .B1(G2897), .B2(new_n1217), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1215), .A2(G213), .A3(G2897), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1260), .B1(new_n1252), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1258), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1230), .B1(new_n1257), .B2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1228), .A2(new_n1258), .A3(new_n1229), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1251), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1265), .B1(new_n1259), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1255), .A2(new_n1266), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1250), .A2(new_n1216), .A3(new_n1254), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1268), .B(new_n1269), .C1(new_n1270), .C2(new_n1262), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1264), .A2(new_n1271), .ZN(G405));
  XNOR2_X1  g1072(.A(G375), .B(G378), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1273), .A2(new_n1251), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1251), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1230), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1274), .A2(new_n1229), .A3(new_n1228), .A4(new_n1275), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(G402));
endmodule


