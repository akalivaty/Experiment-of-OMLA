

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745;

  NOR2_X1 U370 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U371 ( .A(n346), .B(KEYINPUT78), .ZN(n701) );
  OR2_X2 U372 ( .A1(n733), .A2(KEYINPUT2), .ZN(n346) );
  XNOR2_X1 U373 ( .A(n569), .B(KEYINPUT39), .ZN(n602) );
  NOR2_X1 U374 ( .A1(n538), .A2(n539), .ZN(n540) );
  BUF_X1 U375 ( .A(n530), .Z(n351) );
  XNOR2_X1 U376 ( .A(n350), .B(G469), .ZN(n572) );
  NOR2_X2 U377 ( .A1(n636), .A2(G902), .ZN(n350) );
  BUF_X1 U378 ( .A(G128), .Z(n349) );
  BUF_X1 U379 ( .A(G104), .Z(n347) );
  XNOR2_X1 U380 ( .A(n480), .B(KEYINPUT4), .ZN(n449) );
  XNOR2_X1 U381 ( .A(G122), .B(G104), .ZN(n461) );
  INV_X1 U382 ( .A(G953), .ZN(n734) );
  NAND2_X1 U383 ( .A1(n593), .A2(n594), .ZN(n595) );
  XNOR2_X1 U384 ( .A(n686), .B(KEYINPUT76), .ZN(n593) );
  XNOR2_X2 U385 ( .A(n474), .B(n475), .ZN(n538) );
  NAND2_X1 U386 ( .A1(n348), .A2(n598), .ZN(n599) );
  NAND2_X1 U387 ( .A1(n596), .A2(n652), .ZN(n348) );
  INV_X1 U388 ( .A(n648), .ZN(n658) );
  NAND2_X1 U389 ( .A1(n678), .A2(n544), .ZN(n524) );
  XNOR2_X1 U390 ( .A(n523), .B(n522), .ZN(n678) );
  NOR2_X2 U391 ( .A1(n621), .A2(n717), .ZN(n623) );
  NOR2_X2 U392 ( .A1(n630), .A2(n717), .ZN(n631) );
  XOR2_X1 U393 ( .A(n540), .B(KEYINPUT99), .Z(n648) );
  XNOR2_X1 U394 ( .A(n385), .B(n384), .ZN(n745) );
  NOR2_X2 U395 ( .A1(n613), .A2(n717), .ZN(n615) );
  NAND2_X2 U396 ( .A1(n527), .A2(n526), .ZN(n529) );
  NOR2_X1 U397 ( .A1(n699), .A2(n608), .ZN(n702) );
  NOR2_X1 U398 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X2 U399 ( .A1(n742), .A2(n745), .ZN(n577) );
  XNOR2_X1 U400 ( .A(n387), .B(n355), .ZN(n742) );
  OR2_X1 U401 ( .A1(n418), .A2(n533), .ZN(n419) );
  XNOR2_X1 U402 ( .A(n389), .B(n388), .ZN(n533) );
  BUF_X1 U403 ( .A(n634), .Z(n713) );
  XNOR2_X2 U404 ( .A(n529), .B(n528), .ZN(n536) );
  XNOR2_X1 U405 ( .A(n436), .B(G472), .ZN(n530) );
  XNOR2_X2 U406 ( .A(n564), .B(n563), .ZN(n718) );
  OR2_X1 U407 ( .A1(n627), .A2(n379), .ZN(n378) );
  NOR2_X1 U408 ( .A1(n380), .A2(n375), .ZN(n374) );
  INV_X1 U409 ( .A(KEYINPUT19), .ZN(n375) );
  INV_X1 U410 ( .A(G137), .ZN(n429) );
  XOR2_X1 U411 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n477) );
  XOR2_X1 U412 ( .A(G137), .B(G140), .Z(n411) );
  XNOR2_X1 U413 ( .A(n358), .B(G101), .ZN(n444) );
  XNOR2_X1 U414 ( .A(KEYINPUT3), .B(G113), .ZN(n358) );
  NAND2_X1 U415 ( .A1(n364), .A2(n362), .ZN(n361) );
  NAND2_X1 U416 ( .A1(n456), .A2(n365), .ZN(n364) );
  NAND2_X1 U417 ( .A1(n607), .A2(n363), .ZN(n362) );
  NAND2_X1 U418 ( .A1(KEYINPUT2), .A2(n365), .ZN(n363) );
  NOR2_X1 U419 ( .A1(n573), .A2(KEYINPUT19), .ZN(n372) );
  AND2_X1 U420 ( .A1(n377), .A2(KEYINPUT19), .ZN(n376) );
  AND2_X1 U421 ( .A1(n382), .A2(n381), .ZN(n380) );
  NAND2_X1 U422 ( .A1(n459), .A2(n607), .ZN(n381) );
  NAND2_X1 U423 ( .A1(G234), .A2(n734), .ZN(n412) );
  XNOR2_X1 U424 ( .A(n509), .B(KEYINPUT0), .ZN(n547) );
  XNOR2_X1 U425 ( .A(n571), .B(KEYINPUT28), .ZN(n588) );
  AND2_X1 U426 ( .A1(n570), .A2(n351), .ZN(n571) );
  XNOR2_X1 U427 ( .A(n417), .B(n354), .ZN(n388) );
  OR2_X1 U428 ( .A1(n714), .A2(G902), .ZN(n389) );
  INV_X1 U429 ( .A(KEYINPUT65), .ZN(n365) );
  XNOR2_X1 U430 ( .A(G113), .B(G143), .ZN(n468) );
  XOR2_X1 U431 ( .A(KEYINPUT93), .B(G131), .Z(n469) );
  XOR2_X1 U432 ( .A(G107), .B(G110), .Z(n397) );
  XNOR2_X1 U433 ( .A(G101), .B(KEYINPUT83), .ZN(n396) );
  XNOR2_X1 U434 ( .A(KEYINPUT83), .B(KEYINPUT16), .ZN(n441) );
  NOR2_X1 U435 ( .A1(n493), .A2(n492), .ZN(n570) );
  XNOR2_X1 U436 ( .A(n488), .B(n487), .ZN(n501) );
  INV_X1 U437 ( .A(G478), .ZN(n487) );
  XNOR2_X1 U438 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U439 ( .A(n479), .B(n478), .ZN(n483) );
  XNOR2_X1 U440 ( .A(G134), .B(G122), .ZN(n476) );
  XNOR2_X1 U441 ( .A(G125), .B(G146), .ZN(n452) );
  INV_X1 U442 ( .A(n702), .ZN(n368) );
  BUF_X1 U443 ( .A(n678), .Z(n695) );
  NAND2_X1 U444 ( .A1(n380), .A2(n378), .ZN(n504) );
  NOR2_X1 U445 ( .A1(n376), .A2(n374), .ZN(n373) );
  XNOR2_X1 U446 ( .A(n512), .B(n511), .ZN(n554) );
  XNOR2_X1 U447 ( .A(n416), .B(n390), .ZN(n714) );
  INV_X1 U448 ( .A(n731), .ZN(n390) );
  AND2_X1 U449 ( .A1(n612), .A2(G953), .ZN(n717) );
  INV_X1 U450 ( .A(KEYINPUT42), .ZN(n384) );
  AND2_X1 U451 ( .A1(n696), .A2(n587), .ZN(n386) );
  AND2_X1 U452 ( .A1(n682), .A2(n669), .ZN(n352) );
  AND2_X1 U453 ( .A1(n366), .A2(n361), .ZN(n353) );
  XOR2_X1 U454 ( .A(KEYINPUT89), .B(KEYINPUT25), .Z(n354) );
  XOR2_X1 U455 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n355) );
  XOR2_X1 U456 ( .A(KEYINPUT70), .B(KEYINPUT34), .Z(n356) );
  AND2_X1 U457 ( .A1(n607), .A2(n365), .ZN(n357) );
  AND2_X2 U458 ( .A1(n369), .A2(n368), .ZN(n634) );
  XNOR2_X1 U459 ( .A(n732), .B(G146), .ZN(n435) );
  NAND2_X1 U460 ( .A1(n353), .A2(n359), .ZN(n369) );
  NAND2_X1 U461 ( .A1(n360), .A2(n357), .ZN(n359) );
  INV_X1 U462 ( .A(n606), .ZN(n360) );
  NAND2_X1 U463 ( .A1(n606), .A2(n367), .ZN(n366) );
  AND2_X1 U464 ( .A1(n698), .A2(KEYINPUT65), .ZN(n367) );
  NAND2_X1 U465 ( .A1(n373), .A2(n370), .ZN(n589) );
  NAND2_X1 U466 ( .A1(n380), .A2(n371), .ZN(n370) );
  AND2_X1 U467 ( .A1(n378), .A2(n372), .ZN(n371) );
  NAND2_X1 U468 ( .A1(n378), .A2(n679), .ZN(n377) );
  OR2_X1 U469 ( .A1(n459), .A2(n607), .ZN(n379) );
  NAND2_X1 U470 ( .A1(n627), .A2(n459), .ZN(n382) );
  XNOR2_X1 U471 ( .A(n383), .B(n442), .ZN(n414) );
  XNOR2_X2 U472 ( .A(G119), .B(G110), .ZN(n442) );
  XNOR2_X1 U473 ( .A(n413), .B(n349), .ZN(n383) );
  NAND2_X1 U474 ( .A1(n386), .A2(n588), .ZN(n385) );
  NAND2_X1 U475 ( .A1(n602), .A2(n651), .ZN(n387) );
  AND2_X1 U476 ( .A1(n666), .A2(n542), .ZN(n391) );
  AND2_X1 U477 ( .A1(G214), .A2(n470), .ZN(n392) );
  AND2_X1 U478 ( .A1(n514), .A2(n519), .ZN(n393) );
  NOR2_X1 U479 ( .A1(G953), .A2(G237), .ZN(n470) );
  XNOR2_X1 U480 ( .A(n411), .B(n398), .ZN(n399) );
  XNOR2_X1 U481 ( .A(n432), .B(n431), .ZN(n433) );
  NOR2_X1 U482 ( .A1(n501), .A2(n538), .ZN(n503) );
  XNOR2_X1 U483 ( .A(n471), .B(n392), .ZN(n472) );
  XNOR2_X1 U484 ( .A(n473), .B(n472), .ZN(n618) );
  XNOR2_X1 U485 ( .A(n579), .B(KEYINPUT36), .ZN(n580) );
  XNOR2_X1 U486 ( .A(n483), .B(n482), .ZN(n486) );
  XNOR2_X1 U487 ( .A(n581), .B(n580), .ZN(n582) );
  NAND2_X1 U488 ( .A1(n554), .A2(n393), .ZN(n517) );
  XOR2_X1 U489 ( .A(G131), .B(G134), .Z(n394) );
  XNOR2_X1 U490 ( .A(KEYINPUT68), .B(n394), .ZN(n395) );
  XNOR2_X2 U491 ( .A(G143), .B(G128), .ZN(n480) );
  XNOR2_X1 U492 ( .A(n395), .B(n449), .ZN(n732) );
  XOR2_X1 U493 ( .A(n397), .B(n396), .Z(n400) );
  NAND2_X1 U494 ( .A1(G227), .A2(n734), .ZN(n398) );
  XNOR2_X1 U495 ( .A(n400), .B(n399), .ZN(n402) );
  XNOR2_X1 U496 ( .A(n347), .B(KEYINPUT73), .ZN(n401) );
  XNOR2_X1 U497 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U498 ( .A(n435), .B(n403), .ZN(n404) );
  INV_X1 U499 ( .A(n404), .ZN(n636) );
  XNOR2_X1 U500 ( .A(G902), .B(KEYINPUT15), .ZN(n456) );
  NAND2_X1 U501 ( .A1(n456), .A2(G234), .ZN(n407) );
  XNOR2_X1 U502 ( .A(KEYINPUT88), .B(KEYINPUT20), .ZN(n406) );
  XNOR2_X1 U503 ( .A(n407), .B(n406), .ZN(n410) );
  NAND2_X1 U504 ( .A1(n410), .A2(G221), .ZN(n409) );
  XNOR2_X1 U505 ( .A(KEYINPUT90), .B(KEYINPUT21), .ZN(n408) );
  XNOR2_X1 U506 ( .A(n409), .B(n408), .ZN(n518) );
  OR2_X1 U507 ( .A1(n572), .A2(n518), .ZN(n418) );
  NAND2_X1 U508 ( .A1(G217), .A2(n410), .ZN(n417) );
  XNOR2_X1 U509 ( .A(n452), .B(KEYINPUT10), .ZN(n466) );
  XNOR2_X1 U510 ( .A(n411), .B(n466), .ZN(n731) );
  XOR2_X1 U511 ( .A(KEYINPUT8), .B(n412), .Z(n484) );
  NAND2_X1 U512 ( .A1(n484), .A2(G221), .ZN(n415) );
  XNOR2_X1 U513 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n413) );
  XNOR2_X1 U514 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X2 U515 ( .A(KEYINPUT91), .B(n419), .ZN(n567) );
  NAND2_X1 U516 ( .A1(G234), .A2(G237), .ZN(n420) );
  XNOR2_X1 U517 ( .A(KEYINPUT14), .B(n420), .ZN(n423) );
  INV_X1 U518 ( .A(G902), .ZN(n438) );
  NOR2_X1 U519 ( .A1(n734), .A2(n438), .ZN(n421) );
  NAND2_X1 U520 ( .A1(n423), .A2(n421), .ZN(n505) );
  XOR2_X1 U521 ( .A(KEYINPUT105), .B(n505), .Z(n422) );
  NOR2_X1 U522 ( .A1(G900), .A2(n422), .ZN(n426) );
  NAND2_X1 U523 ( .A1(n423), .A2(G952), .ZN(n424) );
  XOR2_X1 U524 ( .A(KEYINPUT85), .B(n424), .Z(n694) );
  NOR2_X1 U525 ( .A1(n694), .A2(G953), .ZN(n425) );
  XNOR2_X1 U526 ( .A(n425), .B(KEYINPUT86), .ZN(n507) );
  NOR2_X1 U527 ( .A1(n426), .A2(n507), .ZN(n493) );
  XOR2_X1 U528 ( .A(KEYINPUT5), .B(KEYINPUT72), .Z(n428) );
  NAND2_X1 U529 ( .A1(n470), .A2(G210), .ZN(n427) );
  XNOR2_X1 U530 ( .A(n428), .B(n427), .ZN(n432) );
  XNOR2_X1 U531 ( .A(G119), .B(G116), .ZN(n430) );
  XNOR2_X1 U532 ( .A(n433), .B(n444), .ZN(n434) );
  XNOR2_X1 U533 ( .A(n435), .B(n434), .ZN(n609) );
  NAND2_X1 U534 ( .A1(n609), .A2(n438), .ZN(n436) );
  INV_X1 U535 ( .A(G237), .ZN(n437) );
  NAND2_X1 U536 ( .A1(n438), .A2(n437), .ZN(n457) );
  NAND2_X1 U537 ( .A1(n457), .A2(G214), .ZN(n679) );
  NAND2_X1 U538 ( .A1(n530), .A2(n679), .ZN(n439) );
  XNOR2_X1 U539 ( .A(KEYINPUT30), .B(n439), .ZN(n440) );
  NOR2_X1 U540 ( .A1(n493), .A2(n440), .ZN(n566) );
  NAND2_X1 U541 ( .A1(n567), .A2(n566), .ZN(n460) );
  XNOR2_X1 U542 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U543 ( .A(n444), .B(n443), .ZN(n447) );
  INV_X1 U544 ( .A(G116), .ZN(n445) );
  XNOR2_X1 U545 ( .A(n445), .B(G107), .ZN(n481) );
  XNOR2_X1 U546 ( .A(n481), .B(n461), .ZN(n446) );
  XNOR2_X1 U547 ( .A(n447), .B(n446), .ZN(n724) );
  NAND2_X1 U548 ( .A1(n734), .A2(G224), .ZN(n448) );
  XNOR2_X1 U549 ( .A(n448), .B(KEYINPUT74), .ZN(n450) );
  XNOR2_X1 U550 ( .A(n450), .B(n449), .ZN(n454) );
  XNOR2_X1 U551 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n451) );
  XNOR2_X1 U552 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U553 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U554 ( .A(n724), .B(n455), .ZN(n627) );
  INV_X1 U555 ( .A(n456), .ZN(n607) );
  NAND2_X1 U556 ( .A1(n457), .A2(G210), .ZN(n458) );
  XNOR2_X1 U557 ( .A(n458), .B(KEYINPUT84), .ZN(n459) );
  OR2_X1 U558 ( .A1(n460), .A2(n504), .ZN(n491) );
  XNOR2_X1 U559 ( .A(KEYINPUT13), .B(G475), .ZN(n475) );
  XOR2_X1 U560 ( .A(n461), .B(KEYINPUT11), .Z(n465) );
  XOR2_X1 U561 ( .A(KEYINPUT95), .B(KEYINPUT12), .Z(n463) );
  XNOR2_X1 U562 ( .A(G140), .B(KEYINPUT94), .ZN(n462) );
  XNOR2_X1 U563 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U564 ( .A(n465), .B(n464), .ZN(n467) );
  XOR2_X1 U565 ( .A(n467), .B(n466), .Z(n473) );
  XNOR2_X1 U566 ( .A(n469), .B(n468), .ZN(n471) );
  NOR2_X1 U567 ( .A1(G902), .A2(n618), .ZN(n474) );
  XNOR2_X1 U568 ( .A(n477), .B(n476), .ZN(n479) );
  XOR2_X1 U569 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n478) );
  XNOR2_X1 U570 ( .A(n480), .B(n481), .ZN(n482) );
  NAND2_X1 U571 ( .A1(G217), .A2(n484), .ZN(n485) );
  XNOR2_X1 U572 ( .A(n486), .B(n485), .ZN(n710) );
  NOR2_X1 U573 ( .A1(G902), .A2(n710), .ZN(n488) );
  AND2_X1 U574 ( .A1(n538), .A2(n501), .ZN(n490) );
  INV_X1 U575 ( .A(KEYINPUT104), .ZN(n489) );
  XNOR2_X1 U576 ( .A(n490), .B(n489), .ZN(n525) );
  NOR2_X1 U577 ( .A1(n491), .A2(n525), .ZN(n583) );
  XOR2_X1 U578 ( .A(n583), .B(G143), .Z(G45) );
  XNOR2_X2 U579 ( .A(n572), .B(KEYINPUT1), .ZN(n666) );
  INV_X1 U580 ( .A(n666), .ZN(n497) );
  INV_X1 U581 ( .A(n518), .ZN(n669) );
  NAND2_X1 U582 ( .A1(n669), .A2(n533), .ZN(n492) );
  XNOR2_X1 U583 ( .A(n351), .B(KEYINPUT6), .ZN(n519) );
  INV_X1 U584 ( .A(n501), .ZN(n539) );
  NAND2_X1 U585 ( .A1(n539), .A2(n538), .ZN(n494) );
  XNOR2_X1 U586 ( .A(KEYINPUT98), .B(n494), .ZN(n655) );
  INV_X1 U587 ( .A(n655), .ZN(n651) );
  NAND2_X1 U588 ( .A1(n679), .A2(n651), .ZN(n495) );
  NOR2_X1 U589 ( .A1(n519), .A2(n495), .ZN(n496) );
  NAND2_X1 U590 ( .A1(n570), .A2(n496), .ZN(n578) );
  NOR2_X1 U591 ( .A1(n497), .A2(n578), .ZN(n499) );
  XNOR2_X1 U592 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n498) );
  XOR2_X1 U593 ( .A(n499), .B(n498), .Z(n500) );
  NAND2_X1 U594 ( .A1(n500), .A2(n504), .ZN(n603) );
  XNOR2_X1 U595 ( .A(n603), .B(G140), .ZN(G42) );
  INV_X1 U596 ( .A(KEYINPUT101), .ZN(n502) );
  XNOR2_X1 U597 ( .A(n503), .B(n502), .ZN(n682) );
  INV_X1 U598 ( .A(n679), .ZN(n573) );
  NOR2_X1 U599 ( .A1(n505), .A2(G898), .ZN(n506) );
  OR2_X1 U600 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U601 ( .A1(n589), .A2(n508), .ZN(n509) );
  INV_X1 U602 ( .A(n547), .ZN(n510) );
  NAND2_X1 U603 ( .A1(n352), .A2(n510), .ZN(n512) );
  INV_X1 U604 ( .A(KEYINPUT22), .ZN(n511) );
  INV_X1 U605 ( .A(KEYINPUT102), .ZN(n513) );
  XNOR2_X1 U606 ( .A(n533), .B(n513), .ZN(n668) );
  NOR2_X1 U607 ( .A1(n666), .A2(n668), .ZN(n514) );
  INV_X1 U608 ( .A(KEYINPUT75), .ZN(n515) );
  XNOR2_X1 U609 ( .A(n515), .B(KEYINPUT32), .ZN(n516) );
  XNOR2_X1 U610 ( .A(n517), .B(n516), .ZN(n535) );
  XNOR2_X1 U611 ( .A(n535), .B(G119), .ZN(G21) );
  XNOR2_X1 U612 ( .A(n547), .B(KEYINPUT87), .ZN(n544) );
  OR2_X1 U613 ( .A1(n533), .A2(n518), .ZN(n665) );
  NOR2_X1 U614 ( .A1(n666), .A2(n665), .ZN(n546) );
  INV_X1 U615 ( .A(n519), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n546), .A2(n551), .ZN(n523) );
  XOR2_X1 U617 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n521) );
  INV_X1 U618 ( .A(KEYINPUT103), .ZN(n520) );
  XNOR2_X1 U619 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U620 ( .A(n524), .B(n356), .ZN(n527) );
  INV_X1 U621 ( .A(n525), .ZN(n526) );
  INV_X1 U622 ( .A(KEYINPUT35), .ZN(n528) );
  XNOR2_X1 U623 ( .A(n536), .B(G122), .ZN(G24) );
  INV_X1 U624 ( .A(n351), .ZN(n542) );
  NAND2_X1 U625 ( .A1(n554), .A2(n391), .ZN(n532) );
  INV_X1 U626 ( .A(KEYINPUT66), .ZN(n531) );
  XNOR2_X1 U627 ( .A(n532), .B(n531), .ZN(n534) );
  NAND2_X1 U628 ( .A1(n534), .A2(n533), .ZN(n632) );
  AND2_X1 U629 ( .A1(n632), .A2(n535), .ZN(n537) );
  NAND2_X1 U630 ( .A1(n537), .A2(n536), .ZN(n560) );
  NAND2_X1 U631 ( .A1(n560), .A2(KEYINPUT44), .ZN(n557) );
  NAND2_X1 U632 ( .A1(n658), .A2(n655), .ZN(n541) );
  XNOR2_X1 U633 ( .A(n541), .B(KEYINPUT100), .ZN(n686) );
  INV_X1 U634 ( .A(n567), .ZN(n543) );
  NOR2_X1 U635 ( .A1(n543), .A2(n351), .ZN(n545) );
  NAND2_X1 U636 ( .A1(n545), .A2(n544), .ZN(n642) );
  NAND2_X1 U637 ( .A1(n546), .A2(n351), .ZN(n674) );
  NOR2_X1 U638 ( .A1(n674), .A2(n547), .ZN(n549) );
  XNOR2_X1 U639 ( .A(KEYINPUT92), .B(KEYINPUT31), .ZN(n548) );
  XNOR2_X1 U640 ( .A(n549), .B(n548), .ZN(n659) );
  NAND2_X1 U641 ( .A1(n642), .A2(n659), .ZN(n550) );
  AND2_X1 U642 ( .A1(n593), .A2(n550), .ZN(n555) );
  NAND2_X1 U643 ( .A1(n666), .A2(n668), .ZN(n552) );
  NOR2_X1 U644 ( .A1(n552), .A2(n551), .ZN(n553) );
  AND2_X1 U645 ( .A1(n554), .A2(n553), .ZN(n640) );
  NOR2_X1 U646 ( .A1(n555), .A2(n640), .ZN(n556) );
  NAND2_X1 U647 ( .A1(n557), .A2(n556), .ZN(n559) );
  INV_X1 U648 ( .A(KEYINPUT79), .ZN(n558) );
  XNOR2_X1 U649 ( .A(n559), .B(n558), .ZN(n562) );
  NOR2_X1 U650 ( .A1(n560), .A2(KEYINPUT44), .ZN(n561) );
  NOR2_X2 U651 ( .A1(n562), .A2(n561), .ZN(n564) );
  XOR2_X1 U652 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n563) );
  INV_X1 U653 ( .A(KEYINPUT38), .ZN(n565) );
  XNOR2_X1 U654 ( .A(n504), .B(n565), .ZN(n574) );
  INV_X1 U655 ( .A(n574), .ZN(n680) );
  AND2_X1 U656 ( .A1(n566), .A2(n680), .ZN(n568) );
  NAND2_X1 U657 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U658 ( .A(n572), .B(KEYINPUT107), .ZN(n587) );
  NOR2_X1 U659 ( .A1(n574), .A2(n573), .ZN(n685) );
  AND2_X1 U660 ( .A1(n682), .A2(n685), .ZN(n576) );
  XNOR2_X1 U661 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n575) );
  XNOR2_X1 U662 ( .A(n576), .B(n575), .ZN(n696) );
  XNOR2_X1 U663 ( .A(n577), .B(KEYINPUT46), .ZN(n586) );
  NOR2_X1 U664 ( .A1(n578), .A2(n504), .ZN(n581) );
  INV_X1 U665 ( .A(KEYINPUT110), .ZN(n579) );
  NOR2_X1 U666 ( .A1(n666), .A2(n582), .ZN(n662) );
  XOR2_X1 U667 ( .A(KEYINPUT77), .B(n583), .Z(n584) );
  NOR2_X1 U668 ( .A1(n662), .A2(n584), .ZN(n585) );
  NAND2_X1 U669 ( .A1(n586), .A2(n585), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n588), .A2(n587), .ZN(n591) );
  INV_X1 U671 ( .A(n589), .ZN(n590) );
  NOR2_X1 U672 ( .A1(n591), .A2(n590), .ZN(n652) );
  NAND2_X1 U673 ( .A1(n686), .A2(n652), .ZN(n592) );
  NAND2_X1 U674 ( .A1(n592), .A2(KEYINPUT47), .ZN(n598) );
  XNOR2_X1 U675 ( .A(KEYINPUT67), .B(KEYINPUT47), .ZN(n594) );
  XNOR2_X1 U676 ( .A(KEYINPUT71), .B(n595), .ZN(n596) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT48), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n602), .A2(n648), .ZN(n664) );
  AND2_X1 U679 ( .A1(n603), .A2(n664), .ZN(n604) );
  AND2_X2 U680 ( .A1(n605), .A2(n604), .ZN(n733) );
  NAND2_X1 U681 ( .A1(n718), .A2(n733), .ZN(n606) );
  INV_X1 U682 ( .A(KEYINPUT2), .ZN(n698) );
  INV_X1 U683 ( .A(n718), .ZN(n699) );
  NAND2_X1 U684 ( .A1(n733), .A2(KEYINPUT2), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n634), .A2(G472), .ZN(n611) );
  XOR2_X1 U686 ( .A(KEYINPUT62), .B(n609), .Z(n610) );
  XNOR2_X1 U687 ( .A(n611), .B(n610), .ZN(n613) );
  INV_X1 U688 ( .A(G952), .ZN(n612) );
  XOR2_X1 U689 ( .A(KEYINPUT80), .B(KEYINPUT63), .Z(n614) );
  XNOR2_X1 U690 ( .A(n615), .B(n614), .ZN(G57) );
  NAND2_X1 U691 ( .A1(n634), .A2(G475), .ZN(n620) );
  XNOR2_X1 U692 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n616), .B(KEYINPUT59), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n620), .B(n619), .ZN(n621) );
  XOR2_X1 U696 ( .A(KEYINPUT121), .B(KEYINPUT60), .Z(n622) );
  XNOR2_X1 U697 ( .A(n623), .B(n622), .ZN(G60) );
  NAND2_X1 U698 ( .A1(n634), .A2(G210), .ZN(n629) );
  XNOR2_X1 U699 ( .A(KEYINPUT82), .B(KEYINPUT54), .ZN(n625) );
  XNOR2_X1 U700 ( .A(KEYINPUT55), .B(KEYINPUT81), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U702 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n631), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U705 ( .A(G110), .B(KEYINPUT113), .Z(n633) );
  XNOR2_X1 U706 ( .A(n632), .B(n633), .ZN(G12) );
  NAND2_X1 U707 ( .A1(n713), .A2(G469), .ZN(n638) );
  XOR2_X1 U708 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n635) );
  XNOR2_X1 U709 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(n639) );
  NOR2_X1 U711 ( .A1(n639), .A2(n717), .ZN(G54) );
  XOR2_X1 U712 ( .A(G101), .B(n640), .Z(G3) );
  NOR2_X1 U713 ( .A1(n655), .A2(n642), .ZN(n641) );
  XOR2_X1 U714 ( .A(n347), .B(n641), .Z(G6) );
  NOR2_X1 U715 ( .A1(n658), .A2(n642), .ZN(n647) );
  XOR2_X1 U716 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n644) );
  XNOR2_X1 U717 ( .A(G107), .B(KEYINPUT26), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U719 ( .A(KEYINPUT27), .B(n645), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(G9) );
  XOR2_X1 U721 ( .A(n349), .B(KEYINPUT29), .Z(n650) );
  NAND2_X1 U722 ( .A1(n652), .A2(n648), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(G30) );
  NAND2_X1 U724 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n653), .B(KEYINPUT114), .ZN(n654) );
  XNOR2_X1 U726 ( .A(G146), .B(n654), .ZN(G48) );
  XNOR2_X1 U727 ( .A(G113), .B(KEYINPUT115), .ZN(n657) );
  NOR2_X1 U728 ( .A1(n655), .A2(n659), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n657), .B(n656), .ZN(G15) );
  NOR2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U731 ( .A(KEYINPUT116), .B(n660), .Z(n661) );
  XNOR2_X1 U732 ( .A(G116), .B(n661), .ZN(G18) );
  XNOR2_X1 U733 ( .A(G125), .B(n662), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n663), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U735 ( .A(G134), .B(n664), .ZN(G36) );
  NAND2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U737 ( .A(n667), .B(KEYINPUT50), .ZN(n673) );
  NOR2_X1 U738 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U739 ( .A(KEYINPUT49), .B(n670), .Z(n671) );
  NOR2_X1 U740 ( .A1(n351), .A2(n671), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U743 ( .A(KEYINPUT51), .B(n676), .Z(n677) );
  NAND2_X1 U744 ( .A1(n696), .A2(n677), .ZN(n691) );
  NOR2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U746 ( .A(KEYINPUT117), .B(n681), .ZN(n683) );
  NAND2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U748 ( .A(n684), .B(KEYINPUT118), .ZN(n688) );
  NAND2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U751 ( .A1(n695), .A2(n689), .ZN(n690) );
  NAND2_X1 U752 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U753 ( .A(KEYINPUT52), .B(n692), .Z(n693) );
  NOR2_X1 U754 ( .A1(n694), .A2(n693), .ZN(n707) );
  NAND2_X1 U755 ( .A1(n696), .A2(n695), .ZN(n705) );
  NAND2_X1 U756 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U757 ( .A1(n701), .A2(n700), .ZN(n703) );
  OR2_X1 U758 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U759 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U760 ( .A1(n734), .A2(n708), .ZN(n709) );
  XOR2_X1 U761 ( .A(KEYINPUT53), .B(n709), .Z(G75) );
  NAND2_X1 U762 ( .A1(n713), .A2(G478), .ZN(n711) );
  XNOR2_X1 U763 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U764 ( .A1(n717), .A2(n712), .ZN(G63) );
  NAND2_X1 U765 ( .A1(n713), .A2(G217), .ZN(n715) );
  XNOR2_X1 U766 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U767 ( .A1(n717), .A2(n716), .ZN(G66) );
  NAND2_X1 U768 ( .A1(n718), .A2(n734), .ZN(n723) );
  NAND2_X1 U769 ( .A1(G224), .A2(G953), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n719), .B(KEYINPUT122), .ZN(n720) );
  XNOR2_X1 U771 ( .A(KEYINPUT61), .B(n720), .ZN(n721) );
  NAND2_X1 U772 ( .A1(n721), .A2(G898), .ZN(n722) );
  NAND2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n729) );
  XOR2_X1 U774 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n725) );
  XNOR2_X1 U775 ( .A(n724), .B(n725), .ZN(n727) );
  NOR2_X1 U776 ( .A1(G898), .A2(n734), .ZN(n726) );
  NOR2_X1 U777 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(n730) );
  XOR2_X1 U779 ( .A(KEYINPUT125), .B(n730), .Z(G69) );
  XOR2_X1 U780 ( .A(n732), .B(n731), .Z(n736) );
  XOR2_X1 U781 ( .A(n736), .B(n733), .Z(n735) );
  NAND2_X1 U782 ( .A1(n735), .A2(n734), .ZN(n741) );
  INV_X1 U783 ( .A(n736), .ZN(n737) );
  XOR2_X1 U784 ( .A(G227), .B(n737), .Z(n738) );
  NAND2_X1 U785 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U786 ( .A1(n739), .A2(G953), .ZN(n740) );
  NAND2_X1 U787 ( .A1(n741), .A2(n740), .ZN(G72) );
  XNOR2_X1 U788 ( .A(n742), .B(G131), .ZN(n743) );
  XNOR2_X1 U789 ( .A(n743), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U790 ( .A(G137), .B(KEYINPUT126), .Z(n744) );
  XNOR2_X1 U791 ( .A(n745), .B(n744), .ZN(G39) );
endmodule

