//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n461), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  AND3_X1   g042(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT3), .B1(KEYINPUT67), .B2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n461), .B1(new_n476), .B2(new_n477), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n480), .B2(G126), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(new_n461), .A3(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n490), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n494), .A2(new_n461), .A3(G138), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n462), .A2(new_n497), .A3(KEYINPUT68), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n478), .B2(G138), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n489), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT69), .A3(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(G543), .A3(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n509), .A2(new_n514), .A3(new_n510), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n503), .A2(new_n511), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n517), .A2(KEYINPUT70), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(KEYINPUT70), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n518), .A2(new_n519), .B1(new_n505), .B2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  INV_X1    g097(.A(new_n511), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G51), .ZN(new_n524));
  INV_X1    g099(.A(new_n515), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n528), .A2(new_n529), .B1(new_n514), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n524), .A2(new_n526), .A3(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  AOI22_X1  g108(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n505), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n523), .A2(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n525), .A2(G90), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  AND2_X1   g114(.A1(G68), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n540), .B1(new_n514), .B2(G56), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n505), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT71), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n525), .A2(G81), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n545), .B1(new_n541), .B2(new_n505), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT72), .B(G43), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n523), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n543), .A2(new_n544), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  AND2_X1   g130(.A1(G53), .A2(G543), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n509), .A2(new_n510), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT73), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n509), .A2(new_n559), .A3(new_n510), .A4(new_n556), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(KEYINPUT9), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n515), .A2(KEYINPUT74), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n509), .A2(new_n563), .A3(new_n514), .A4(new_n510), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(G91), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n557), .A2(KEYINPUT73), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n505), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n561), .A2(new_n565), .A3(new_n567), .A4(new_n569), .ZN(G299));
  OR2_X1    g145(.A1(new_n514), .A2(G74), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n523), .A2(G49), .B1(new_n571), .B2(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n562), .A2(new_n564), .ZN(new_n573));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n512), .A2(new_n513), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n523), .A2(G48), .B1(new_n579), .B2(G651), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n573), .B2(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(G72), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G60), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n577), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n505), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n587), .B1(new_n586), .B2(new_n585), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n523), .A2(G47), .B1(new_n525), .B2(G85), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  XOR2_X1   g167(.A(KEYINPUT76), .B(G66), .Z(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n577), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n523), .A2(G54), .B1(new_n594), .B2(G651), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n562), .A2(new_n596), .A3(G92), .A4(new_n564), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT10), .B1(new_n573), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G284));
  XOR2_X1   g177(.A(G284), .B(KEYINPUT77), .Z(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT78), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G299), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(G280));
  XOR2_X1   g183(.A(G280), .B(KEYINPUT79), .Z(G297));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n601), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n598), .A2(new_n600), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n612), .A2(KEYINPUT80), .A3(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT80), .B1(new_n612), .B2(G559), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  MUX2_X1   g190(.A(new_n549), .B(new_n615), .S(G868), .Z(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n462), .A2(new_n466), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(G123), .A2(new_n480), .B1(new_n478), .B2(G135), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(G111), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n624), .A2(KEYINPUT81), .B1(new_n625), .B2(G2105), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(KEYINPUT81), .B2(new_n624), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G2096), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n639), .A2(new_n642), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT83), .ZN(new_n648));
  INV_X1    g223(.A(G14), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n643), .A2(new_n646), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n649), .B1(new_n650), .B2(new_n644), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  INV_X1    g228(.A(KEYINPUT18), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n621), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n629), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n669), .B2(new_n675), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT84), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT85), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n684), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n667), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n681), .A2(new_n684), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n681), .A2(new_n684), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n666), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(G229));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G33), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT25), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  AOI22_X1  g271(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n478), .A2(KEYINPUT89), .A3(G139), .ZN(new_n698));
  AOI21_X1  g273(.A(KEYINPUT89), .B1(new_n478), .B2(G139), .ZN(new_n699));
  OAI221_X1 g274(.A(new_n696), .B1(new_n461), .B2(new_n697), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT90), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n693), .B1(new_n702), .B2(new_n692), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT91), .B(G2072), .Z(new_n704));
  XOR2_X1   g279(.A(new_n703), .B(new_n704), .Z(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT30), .B(G28), .ZN(new_n706));
  OR2_X1    g281(.A1(KEYINPUT31), .A2(G11), .ZN(new_n707));
  NAND2_X1  g282(.A1(KEYINPUT31), .A2(G11), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n706), .A2(new_n692), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n628), .B2(new_n692), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT26), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n713), .A2(new_n714), .B1(G105), .B2(new_n466), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n478), .A2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n480), .A2(G129), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(new_n692), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n692), .B2(G32), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT27), .B(G1996), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n710), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G2084), .ZN(new_n724));
  NAND2_X1  g299(.A1(G160), .A2(G29), .ZN(new_n725));
  AND2_X1   g300(.A1(KEYINPUT24), .A2(G34), .ZN(new_n726));
  NOR2_X1   g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n692), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT92), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G5), .A2(G16), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT93), .Z(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(G301), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n723), .B1(new_n724), .B2(new_n730), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n692), .A2(G26), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT88), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n478), .A2(G140), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n480), .A2(G128), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n461), .A2(G116), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n740), .B(new_n741), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n739), .B1(G29), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2067), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n550), .A2(G16), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G16), .B2(G19), .ZN(new_n748));
  INV_X1    g323(.A(G1341), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n721), .A2(new_n722), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n735), .B2(new_n734), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n730), .A2(new_n724), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT94), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n733), .A2(G21), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G168), .B2(new_n733), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n752), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  OR4_X1    g334(.A1(new_n705), .A2(new_n736), .A3(new_n750), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n692), .A2(G27), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G164), .B2(new_n692), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2078), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n748), .B2(new_n749), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n692), .A2(G35), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G162), .B2(new_n692), .ZN(new_n766));
  INV_X1    g341(.A(G2090), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G4), .A2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n601), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT87), .B(G1348), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(G299), .A2(G16), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n733), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n760), .A2(new_n771), .A3(new_n775), .A4(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n733), .A2(G23), .ZN(new_n784));
  INV_X1    g359(.A(G288), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n733), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT33), .ZN(new_n787));
  INV_X1    g362(.A(G1976), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(G166), .A2(G16), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G16), .B2(G22), .ZN(new_n791));
  INV_X1    g366(.A(G1971), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G6), .B(G305), .S(G16), .Z(new_n794));
  XOR2_X1   g369(.A(KEYINPUT32), .B(G1981), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n791), .B2(new_n792), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n789), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT34), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n692), .A2(G25), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n478), .A2(G131), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n480), .A2(G119), .ZN(new_n803));
  OR2_X1    g378(.A1(G95), .A2(G2105), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n804), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n801), .B1(new_n807), .B2(new_n692), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT35), .B(G1991), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G24), .B(G290), .S(G16), .Z(new_n811));
  XOR2_X1   g386(.A(KEYINPUT86), .B(G1986), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n800), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n798), .A2(new_n799), .ZN(new_n815));
  OR3_X1    g390(.A1(new_n814), .A2(KEYINPUT36), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT36), .B1(new_n814), .B2(new_n815), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n783), .B1(new_n816), .B2(new_n817), .ZN(G311));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(new_n782), .ZN(G150));
  NAND2_X1  g395(.A1(new_n601), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n523), .A2(G55), .B1(new_n525), .B2(G93), .ZN(new_n823));
  INV_X1    g398(.A(G67), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n512), .B2(new_n513), .ZN(new_n825));
  AND2_X1   g400(.A1(G80), .A2(G543), .ZN(new_n826));
  OR3_X1    g401(.A1(new_n825), .A2(KEYINPUT97), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(KEYINPUT97), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n827), .A2(G651), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n830), .A2(new_n549), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n549), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n822), .B(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n835), .A2(new_n836), .A3(G860), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n830), .A2(G860), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n837), .A2(new_n839), .ZN(G145));
  NAND2_X1  g415(.A1(new_n478), .A2(G142), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n480), .A2(G130), .ZN(new_n842));
  OR2_X1    g417(.A1(G106), .A2(G2105), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n501), .B(new_n744), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n718), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n501), .B(new_n744), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(new_n719), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n848), .A2(new_n700), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n701), .B1(new_n848), .B2(new_n850), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n846), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n619), .ZN(new_n854));
  INV_X1    g429(.A(new_n850), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n849), .A2(new_n719), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n702), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n848), .A2(new_n700), .A3(new_n850), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n845), .A3(new_n858), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n853), .A2(new_n854), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n854), .B1(new_n853), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n806), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n859), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n845), .B1(new_n857), .B2(new_n858), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n619), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n853), .A2(new_n854), .A3(new_n859), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n807), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n862), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(G160), .B(KEYINPUT98), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G162), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n628), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G37), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n862), .A2(new_n867), .A3(new_n868), .A4(new_n872), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g453(.A(new_n615), .B1(new_n831), .B2(new_n832), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n613), .A2(new_n614), .A3(new_n833), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n882));
  OR2_X1    g457(.A1(G299), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(G299), .A2(new_n882), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n601), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n612), .A2(new_n882), .A3(G299), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n886), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n879), .A2(new_n880), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(G303), .B(G290), .ZN(new_n895));
  XNOR2_X1  g470(.A(G305), .B(G288), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n895), .B(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n895), .B(new_n896), .ZN(new_n901));
  INV_X1    g476(.A(new_n899), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n894), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n900), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(new_n889), .A3(new_n893), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(G868), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT102), .B1(new_n830), .B2(new_n606), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT102), .A4(G868), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(G295));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n909), .A2(new_n912), .A3(new_n910), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n909), .B2(new_n910), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(G331));
  OAI21_X1  g490(.A(G171), .B1(new_n831), .B2(new_n832), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n548), .A2(new_n546), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n542), .A2(KEYINPUT71), .B1(new_n525), .B2(G81), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n829), .A4(new_n823), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n830), .A2(new_n549), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(G301), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(G168), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n919), .A2(new_n920), .A3(G301), .ZN(new_n923));
  AOI21_X1  g498(.A(G301), .B1(new_n919), .B2(new_n920), .ZN(new_n924));
  OAI21_X1  g499(.A(G286), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n892), .A2(new_n890), .A3(new_n922), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n888), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n875), .B1(new_n929), .B2(new_n898), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n926), .A2(new_n932), .A3(new_n928), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n898), .B1(new_n926), .B2(new_n932), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT105), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n886), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT41), .B1(new_n885), .B2(new_n886), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n927), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n901), .B1(new_n939), .B2(KEYINPUT104), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n926), .A2(new_n932), .A3(new_n928), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n931), .B1(new_n935), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT105), .B1(new_n933), .B2(new_n934), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n940), .A2(new_n936), .A3(new_n941), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n930), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n930), .B1(new_n929), .B2(new_n898), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n949), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n944), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  AOI211_X1 g529(.A(KEYINPUT43), .B(new_n930), .C1(new_n946), .C2(new_n947), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n952), .A2(new_n949), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(G397));
  XNOR2_X1  g533(.A(KEYINPUT119), .B(G1961), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G40), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n465), .A2(new_n472), .A3(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(G138), .B(new_n461), .C1(new_n468), .C2(new_n469), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT4), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n496), .A3(new_n498), .ZN(new_n965));
  AOI21_X1  g540(.A(G1384), .B1(new_n965), .B2(new_n489), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n962), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI211_X1 g544(.A(KEYINPUT50), .B(G1384), .C1(new_n965), .C2(new_n489), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n960), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(G160), .A2(G40), .ZN(new_n973));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n501), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT111), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n966), .A2(new_n980), .A3(KEYINPUT45), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(G2078), .ZN(new_n983));
  AND4_X1   g558(.A1(new_n977), .A2(new_n979), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G2078), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n978), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n966), .A2(KEYINPUT45), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n966), .A2(new_n986), .A3(KEYINPUT45), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n985), .B(new_n962), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n972), .B(new_n984), .C1(new_n991), .C2(new_n982), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT120), .B1(new_n992), .B2(G301), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n982), .ZN(new_n994));
  INV_X1    g569(.A(new_n972), .ZN(new_n995));
  INV_X1    g570(.A(new_n984), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n998), .A3(G171), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n977), .A2(new_n981), .A3(new_n979), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n968), .A2(new_n970), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n1003), .A2(new_n757), .B1(new_n1004), .B2(new_n724), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n1005), .B2(G168), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n757), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n724), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G286), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1001), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1007), .A2(G168), .A3(new_n1008), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(G8), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(KEYINPUT51), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT62), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(G166), .B2(new_n1002), .ZN(new_n1017));
  NAND3_X1  g592(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n962), .B1(new_n989), .B2(new_n990), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1021), .A2(new_n792), .B1(new_n767), .B2(new_n1004), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1020), .B1(new_n1022), .B2(new_n1002), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1004), .A2(new_n767), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n975), .A2(new_n976), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(new_n986), .A3(new_n978), .ZN(new_n1026));
  INV_X1    g601(.A(new_n990), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n973), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1024), .B1(new_n1028), .B2(G1971), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(G8), .A3(new_n1019), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n966), .A2(new_n962), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1031), .B(G8), .C1(G288), .C2(new_n788), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT52), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n785), .B2(G1976), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1031), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(new_n1002), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n579), .A2(G651), .ZN(new_n1039));
  INV_X1    g614(.A(G48), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(new_n511), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n515), .A2(new_n581), .ZN(new_n1042));
  OAI21_X1  g617(.A(G1981), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1981), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n580), .B(new_n1044), .C1(new_n581), .C2(new_n573), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1045), .A3(KEYINPUT49), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT49), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT110), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1048), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(new_n1038), .A4(new_n1046), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1036), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1023), .A2(new_n1030), .A3(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1005), .A2(G168), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT51), .B1(new_n1013), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT62), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1006), .A2(new_n1001), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1000), .A2(new_n1015), .A3(new_n1054), .A4(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G168), .A2(G8), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1005), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1023), .A2(new_n1030), .A3(new_n1053), .A4(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1005), .A2(new_n1064), .A3(new_n1061), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1053), .A2(new_n1030), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1022), .B2(new_n1002), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1029), .A2(KEYINPUT112), .A3(G8), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1020), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1065), .A2(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1074), .A2(new_n1030), .A3(new_n1036), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n785), .A2(new_n788), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1045), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1075), .B1(new_n1038), .B2(new_n1077), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1060), .A2(new_n1073), .A3(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n962), .B(new_n1080), .C1(new_n989), .C2(new_n990), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1004), .A2(G1956), .ZN(new_n1082));
  XOR2_X1   g657(.A(G299), .B(KEYINPUT57), .Z(new_n1083));
  AND3_X1   g658(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G2067), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1037), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT113), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1004), .A2(G1348), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n601), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1083), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1084), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n601), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1087), .A2(KEYINPUT60), .A3(new_n612), .A4(new_n1088), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1096), .A2(new_n1097), .B1(new_n1095), .B2(new_n1089), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT114), .B(G1996), .Z(new_n1101));
  NOR2_X1   g676(.A1(new_n973), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n989), .B2(new_n990), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT115), .B(KEYINPUT58), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(new_n749), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1031), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1100), .B1(new_n1107), .B2(new_n550), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1102), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1106), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1100), .B(new_n550), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1099), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1083), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1084), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1093), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n550), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT116), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(KEYINPUT59), .A3(new_n1112), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1114), .A2(new_n1117), .A3(new_n1119), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1098), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1126), .A2(KEYINPUT117), .A3(new_n1122), .A4(new_n1114), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1094), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n985), .B1(new_n982), .B2(KEYINPUT122), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(KEYINPUT122), .B2(new_n985), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n966), .B2(KEYINPUT45), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n977), .A2(KEYINPUT121), .ZN(new_n1132));
  OAI211_X1 g707(.A(KEYINPUT121), .B(new_n962), .C1(new_n966), .C2(KEYINPUT45), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1131), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n994), .A2(G301), .A3(new_n995), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT123), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n972), .B1(new_n991), .B2(new_n982), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1138), .A2(new_n1139), .A3(G301), .A4(new_n1135), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n993), .A2(new_n999), .A3(new_n1137), .A4(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1054), .A2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g720(.A(G2078), .B(new_n973), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n995), .B(new_n1135), .C1(new_n1146), .C2(KEYINPUT53), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT124), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1138), .A2(new_n1149), .A3(new_n1135), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(G171), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n992), .B2(G301), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1151), .A2(KEYINPUT125), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT125), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1143), .B(new_n1145), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1079), .B1(new_n1128), .B2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n744), .B(G2067), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT107), .ZN(new_n1159));
  INV_X1    g734(.A(G1996), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n718), .B(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n806), .B(new_n809), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT108), .Z(new_n1164));
  NOR2_X1   g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(G290), .B(G1986), .Z(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1025), .A2(new_n973), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1157), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1168), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1171), .A2(G1986), .A3(G290), .ZN(new_n1172));
  XOR2_X1   g747(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1173));
  XNOR2_X1  g748(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1165), .A2(new_n1171), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1171), .B1(new_n1159), .B2(new_n719), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1168), .A2(KEYINPUT46), .A3(new_n1160), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT46), .B1(new_n1168), .B2(new_n1160), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT47), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n807), .A2(new_n809), .ZN(new_n1182));
  OAI22_X1  g757(.A1(new_n1162), .A2(new_n1182), .B1(G2067), .B2(new_n744), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1176), .B(new_n1181), .C1(new_n1168), .C2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1170), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g760(.A(G229), .ZN(new_n1187));
  NOR2_X1   g761(.A1(G227), .A2(new_n459), .ZN(new_n1188));
  INV_X1    g762(.A(new_n1188), .ZN(new_n1189));
  OAI21_X1  g763(.A(KEYINPUT127), .B1(G401), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n1191));
  NAND3_X1  g765(.A1(new_n652), .A2(new_n1191), .A3(new_n1188), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n877), .A2(new_n1187), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g768(.A1(new_n955), .A2(new_n956), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1194), .A2(new_n1195), .ZN(G308));
  AOI21_X1  g770(.A(G229), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1197));
  OAI211_X1 g771(.A(new_n1197), .B(new_n877), .C1(new_n956), .C2(new_n955), .ZN(G225));
endmodule


