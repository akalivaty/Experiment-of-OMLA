//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT75), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT22), .B(G137), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G140), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n198), .A3(KEYINPUT74), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT74), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n197), .A3(G140), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(KEYINPUT16), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT16), .B1(new_n195), .B2(G125), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G119), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G128), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT24), .B(G110), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n209), .B2(G128), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n216));
  INV_X1    g030(.A(G110), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n210), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  XNOR2_X1  g033(.A(G125), .B(G140), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n213), .A2(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n206), .A2(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n202), .A2(new_n219), .A3(new_n204), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n219), .B1(new_n202), .B2(new_n204), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n211), .A2(new_n212), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n215), .A2(new_n210), .A3(new_n216), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT73), .A3(G110), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT73), .B1(new_n227), .B2(G110), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n222), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n194), .B1(new_n232), .B2(KEYINPUT76), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(KEYINPUT76), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT76), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n235), .B(new_n222), .C1(new_n225), .C2(new_n231), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n233), .B1(new_n237), .B2(new_n194), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT25), .B1(new_n238), .B2(new_n188), .ZN(new_n239));
  INV_X1    g053(.A(new_n236), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n227), .A2(G110), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT73), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n228), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n244), .B(new_n226), .C1(new_n223), .C2(new_n224), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n235), .B1(new_n245), .B2(new_n222), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n194), .B1(new_n240), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n233), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n189), .B1(new_n239), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n238), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n189), .A2(G902), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n256));
  XOR2_X1   g070(.A(G116), .B(G119), .Z(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT2), .B(G113), .ZN(new_n258));
  OR2_X1    g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n258), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n219), .A2(G143), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT66), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n266), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n268), .A2(new_n262), .A3(new_n264), .A4(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT0), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n207), .A3(KEYINPUT64), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT64), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(KEYINPUT0), .B2(G128), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n268), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT65), .B1(new_n263), .B2(G146), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n219), .A3(G143), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(new_n278), .A3(new_n264), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n267), .A2(new_n270), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(G137), .ZN(new_n283));
  INV_X1    g097(.A(G137), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT11), .A3(G134), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(G137), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT67), .A2(G131), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n283), .A2(new_n285), .A3(new_n288), .A4(new_n286), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n280), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT1), .B1(new_n263), .B2(G146), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n262), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(G128), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n265), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n298), .A2(new_n279), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n286), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n282), .A2(G137), .ZN(new_n303));
  OAI21_X1  g117(.A(G131), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n287), .B2(G131), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n261), .B1(new_n293), .B2(new_n306), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n290), .A2(KEYINPUT69), .A3(new_n291), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT69), .B1(new_n290), .B2(new_n291), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n280), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n261), .ZN(new_n311));
  OAI21_X1  g125(.A(G128), .B1(new_n294), .B2(new_n295), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT68), .B1(new_n262), .B2(KEYINPUT1), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n279), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n300), .A2(new_n262), .A3(new_n264), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n287), .A2(G131), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n304), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n310), .A2(new_n311), .A3(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n307), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n321));
  OAI21_X1  g135(.A(new_n256), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n319), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n323), .B1(new_n319), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n321), .B1(new_n307), .B2(new_n319), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT71), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n322), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(G237), .A2(G953), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G210), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT27), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT26), .B(G101), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT30), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n293), .B2(new_n306), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n310), .A2(KEYINPUT30), .A3(new_n318), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n261), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n335), .A3(new_n319), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT31), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n340), .A2(KEYINPUT31), .A3(new_n335), .A4(new_n319), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n330), .A2(new_n336), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(G472), .A2(G902), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT32), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n319), .A2(new_n324), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT72), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n319), .A2(new_n323), .A3(new_n324), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n350), .B(new_n351), .C1(new_n328), .C2(KEYINPUT71), .ZN(new_n352));
  INV_X1    g166(.A(new_n329), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n336), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n343), .A2(new_n344), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT32), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n346), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n348), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n340), .A2(new_n319), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n360), .B2(new_n336), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n330), .B2(new_n336), .ZN(new_n362));
  INV_X1    g176(.A(new_n319), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n311), .B1(new_n310), .B2(new_n318), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT28), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n335), .A2(KEYINPUT29), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n327), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n367), .A2(new_n188), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G472), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n255), .B1(new_n359), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G469), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT79), .B1(new_n308), .B2(new_n309), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT69), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n292), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n290), .A2(KEYINPUT69), .A3(new_n291), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G107), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(G104), .ZN(new_n381));
  NOR2_X1   g195(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(G104), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(G107), .ZN(new_n387));
  NAND2_X1  g201(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n387), .B1(new_n389), .B2(new_n382), .ZN(new_n390));
  INV_X1    g204(.A(G101), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(G107), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n384), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT10), .B1(new_n301), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n384), .B1(new_n383), .B2(new_n388), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n393), .B1(new_n387), .B2(new_n382), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n394), .B1(new_n400), .B2(new_n391), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT10), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n207), .B1(new_n262), .B2(KEYINPUT1), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n315), .B1(new_n299), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n407), .B(G101), .C1(new_n398), .C2(new_n399), .ZN(new_n408));
  OAI211_X1 g222(.A(KEYINPUT78), .B(G101), .C1(new_n398), .C2(new_n399), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n392), .A3(KEYINPUT4), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n391), .B1(new_n385), .B2(new_n390), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT78), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n280), .B(new_n408), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n379), .A2(new_n406), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G110), .B(G140), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n190), .A2(G227), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n301), .A2(new_n396), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n404), .A2(new_n392), .A3(new_n395), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n420), .A2(new_n421), .B1(new_n377), .B2(new_n375), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT80), .B1(new_n422), .B2(KEYINPUT12), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n421), .B1(new_n401), .B2(new_n316), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n375), .A2(new_n377), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT80), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT12), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n424), .A2(KEYINPUT12), .A3(new_n292), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n419), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n406), .A2(new_n413), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n425), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n418), .B1(new_n434), .B2(new_n414), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n372), .B(new_n188), .C1(new_n432), .C2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n419), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n434), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n379), .A2(new_n406), .A3(new_n413), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n430), .B2(new_n431), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n438), .B(G469), .C1(new_n440), .C2(new_n418), .ZN(new_n441));
  NAND2_X1  g255(.A1(G469), .A2(G902), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT9), .B(G234), .ZN(new_n444));
  OAI21_X1  g258(.A(G221), .B1(new_n444), .B2(G902), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n190), .A2(G952), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(G234), .B2(G237), .ZN(new_n449));
  NAND2_X1  g263(.A1(G234), .A2(G237), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(G902), .A3(G953), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(G898), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G122), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n261), .A2(new_n408), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n409), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n459));
  INV_X1    g273(.A(new_n412), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n209), .A3(G116), .ZN(new_n463));
  OAI211_X1 g277(.A(G113), .B(new_n463), .C1(new_n257), .C2(new_n462), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n259), .A2(new_n464), .A3(new_n392), .A4(new_n395), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n457), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n410), .A2(new_n412), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n465), .B(new_n456), .C1(new_n468), .C2(new_n458), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n470));
  OR3_X1    g284(.A1(new_n280), .A2(KEYINPUT81), .A3(new_n197), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT81), .B1(new_n280), .B2(new_n197), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n314), .A2(new_n197), .A3(new_n315), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G224), .ZN(new_n475));
  OR3_X1    g289(.A1(new_n475), .A2(KEYINPUT82), .A3(G953), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT82), .B1(new_n475), .B2(G953), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n478), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n471), .A2(new_n472), .A3(new_n480), .A4(new_n473), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n483), .B(new_n457), .C1(new_n461), .C2(new_n466), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n470), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n464), .A2(new_n259), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n396), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n465), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n456), .B(KEYINPUT8), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n473), .B1(new_n197), .B2(new_n280), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n480), .A2(KEYINPUT7), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n488), .A2(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(new_n478), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(new_n493), .B2(new_n478), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n471), .A2(new_n472), .A3(new_n473), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n469), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n497), .A2(new_n188), .ZN(new_n498));
  OAI21_X1  g312(.A(G210), .B1(G237), .B2(G902), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT84), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n485), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(new_n485), .B2(new_n498), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n447), .B(new_n455), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n444), .A2(new_n187), .A3(G953), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n263), .A2(G128), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT13), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n207), .A2(G143), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT88), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT88), .B1(new_n207), .B2(G143), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(G134), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n282), .B(new_n507), .C1(new_n512), .C2(new_n513), .ZN(new_n516));
  INV_X1    g330(.A(G122), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G116), .ZN(new_n518));
  INV_X1    g332(.A(G116), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G122), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(G107), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n515), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n380), .B1(new_n518), .B2(KEYINPUT14), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n525), .A2(new_n521), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n521), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G134), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n516), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n506), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n516), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n526), .A3(new_n527), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n523), .A3(new_n505), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G478), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT89), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  AOI211_X1 g358(.A(G902), .B(new_n542), .C1(new_n532), .C2(new_n535), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n202), .A2(new_n219), .A3(new_n204), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n331), .A2(G143), .A3(G214), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(G143), .B1(new_n331), .B2(G214), .ZN(new_n550));
  OAI21_X1  g364(.A(G131), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n551), .A2(KEYINPUT17), .ZN(new_n552));
  INV_X1    g366(.A(G237), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n190), .A3(G214), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n263), .ZN(new_n555));
  INV_X1    g369(.A(G131), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n548), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT17), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n547), .B(new_n206), .C1(new_n552), .C2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(G113), .B(G122), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(new_n386), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n548), .ZN(new_n562));
  NAND2_X1  g376(.A1(KEYINPUT18), .A2(G131), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n195), .A2(KEYINPUT74), .A3(G125), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(new_n220), .B2(KEYINPUT74), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT85), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(G146), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(G146), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n220), .B2(new_n219), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n564), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n559), .A2(new_n561), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n561), .B1(new_n559), .B2(new_n572), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n188), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G475), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT20), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n551), .A2(new_n557), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n199), .A2(KEYINPUT19), .A3(new_n201), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT86), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT19), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n220), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n220), .B2(new_n581), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n206), .B(new_n578), .C1(new_n584), .C2(G146), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n572), .ZN(new_n586));
  INV_X1    g400(.A(new_n561), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n559), .A2(new_n561), .A3(new_n572), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(G475), .A2(G902), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT87), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n577), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  AOI211_X1 g408(.A(KEYINPUT20), .B(new_n592), .C1(new_n588), .C2(new_n589), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n546), .B(new_n576), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n446), .A2(new_n504), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n371), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  NAND2_X1  g413(.A1(new_n356), .A2(new_n346), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n345), .A2(G902), .ZN(new_n601));
  INV_X1    g415(.A(G472), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n603), .A2(new_n255), .A3(new_n446), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n576), .B1(new_n594), .B2(new_n595), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n535), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n505), .B1(new_n534), .B2(new_n523), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT33), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n532), .A2(new_n610), .A3(new_n535), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(G478), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n537), .A2(new_n188), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n536), .B2(new_n537), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n504), .A2(new_n606), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n604), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(new_n386), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  INV_X1    g434(.A(new_n594), .ZN(new_n621));
  INV_X1    g435(.A(new_n595), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT91), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT91), .B1(new_n594), .B2(new_n595), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n544), .A2(new_n545), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n624), .A2(new_n625), .A3(new_n576), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n447), .ZN(new_n629));
  INV_X1    g443(.A(new_n503), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n485), .A2(new_n498), .A3(new_n501), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n628), .A2(new_n632), .A3(KEYINPUT92), .A4(new_n455), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT92), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(new_n504), .B2(new_n627), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n604), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  NAND2_X1  g453(.A1(new_n356), .A2(new_n188), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n640), .A2(G472), .B1(new_n356), .B2(new_n346), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n194), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n232), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n253), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT93), .B1(new_n251), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n189), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n247), .A2(new_n188), .A3(new_n248), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT25), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n646), .B1(new_n649), .B2(new_n249), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT93), .ZN(new_n651));
  INV_X1    g465(.A(new_n644), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n597), .A2(new_n641), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  AOI21_X1  g471(.A(new_n357), .B1(new_n356), .B2(new_n346), .ZN(new_n658));
  AOI211_X1 g472(.A(KEYINPUT32), .B(new_n347), .C1(new_n354), .C2(new_n355), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n370), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n446), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n447), .B1(new_n502), .B2(new_n503), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n190), .A2(G900), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(G902), .A3(new_n450), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT94), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n666), .A2(new_n667), .A3(new_n449), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n669), .A2(KEYINPUT95), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(KEYINPUT95), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n662), .A2(new_n627), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n660), .A2(new_n654), .A3(new_n661), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  OAI21_X1  g490(.A(new_n336), .B1(new_n363), .B2(new_n364), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n677), .A2(KEYINPUT97), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT97), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n341), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n602), .B1(new_n680), .B2(new_n188), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n658), .B2(new_n659), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT98), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n681), .B1(new_n348), .B2(new_n358), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT98), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n502), .A2(new_n503), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n251), .A2(new_n644), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n605), .A2(new_n626), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n692), .A2(new_n629), .A3(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT40), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n672), .B(KEYINPUT39), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n661), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n661), .A2(new_n697), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n688), .A2(new_n695), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  AND2_X1   g516(.A1(new_n612), .A2(new_n614), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n605), .A2(new_n703), .A3(new_n672), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n662), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n660), .A2(new_n654), .A3(new_n661), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT99), .B(G146), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G48));
  NOR2_X1   g522(.A1(new_n432), .A2(new_n435), .ZN(new_n709));
  OAI21_X1  g523(.A(G469), .B1(new_n709), .B2(G902), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n445), .A3(new_n436), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n371), .A2(new_n616), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND2_X1  g529(.A1(new_n371), .A2(new_n712), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n633), .A2(new_n635), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n519), .ZN(G18));
  OAI21_X1  g533(.A(new_n651), .B1(new_n650), .B2(new_n652), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n251), .A2(KEYINPUT93), .A3(new_n644), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n596), .A2(new_n454), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n723), .A2(new_n662), .A3(new_n711), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n660), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT100), .B(G119), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G21));
  INV_X1    g541(.A(KEYINPUT101), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n693), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n605), .A2(KEYINPUT101), .A3(new_n626), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n504), .ZN(new_n732));
  INV_X1    g546(.A(new_n255), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n327), .A2(new_n365), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n336), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n347), .B1(new_n735), .B2(new_n355), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n640), .B2(G472), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n732), .A2(new_n733), .A3(new_n712), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  NOR2_X1   g553(.A1(new_n711), .A2(new_n662), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT102), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n704), .B(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n740), .A2(new_n742), .A3(new_n737), .A4(new_n692), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  NOR3_X1   g558(.A1(new_n502), .A2(new_n503), .A3(new_n629), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n442), .B(KEYINPUT103), .Z(new_n746));
  NAND3_X1  g560(.A1(new_n436), .A2(new_n441), .A3(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n745), .A2(new_n445), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n660), .A2(new_n748), .A3(new_n742), .A4(new_n733), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n371), .A2(KEYINPUT42), .A3(new_n742), .A4(new_n748), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NOR2_X1   g568(.A1(new_n627), .A2(new_n673), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n660), .A2(new_n748), .A3(new_n733), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  INV_X1    g571(.A(new_n445), .ZN(new_n758));
  INV_X1    g572(.A(new_n436), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n438), .B1(new_n440), .B2(new_n418), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n372), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n746), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n759), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n764), .A2(KEYINPUT46), .A3(new_n746), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n758), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(new_n697), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n745), .B(KEYINPUT105), .Z(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n605), .A2(KEYINPUT43), .A3(new_n615), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n615), .B1(new_n605), .B2(KEYINPUT104), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(KEYINPUT104), .B2(new_n605), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n773), .B1(new_n775), .B2(KEYINPUT43), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n603), .A3(new_n692), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT44), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n776), .A2(new_n779), .A3(new_n603), .A4(new_n692), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n772), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n770), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  INV_X1    g597(.A(new_n745), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n660), .A2(new_n733), .A3(new_n704), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n769), .A2(KEYINPUT47), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n787), .B(new_n758), .C1(new_n767), .C2(new_n768), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n785), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT106), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT106), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n791), .B(new_n785), .C1(new_n786), .C2(new_n788), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(KEYINPUT107), .B(G140), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(G42));
  AND2_X1   g609(.A1(new_n767), .A2(new_n768), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n787), .B1(new_n796), .B2(new_n758), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n710), .A2(new_n436), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT108), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n758), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n769), .A2(KEYINPUT47), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n601), .A2(new_n602), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n255), .A3(new_n736), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n804), .A2(new_n449), .A3(new_n776), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(new_n771), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(KEYINPUT51), .A3(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n691), .A2(new_n447), .A3(new_n711), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n805), .A2(KEYINPUT50), .A3(new_n808), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n712), .A2(KEYINPUT116), .A3(new_n745), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n784), .B2(new_n711), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n813), .A2(new_n449), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n776), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n737), .A2(new_n692), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n811), .A2(new_n812), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n688), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n816), .A3(new_n733), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n821), .A2(new_n816), .A3(KEYINPUT117), .A4(new_n733), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n606), .A3(new_n615), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT118), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n807), .A2(new_n820), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n824), .A2(new_n605), .A3(new_n703), .A4(new_n825), .ZN(new_n830));
  XNOR2_X1  g644(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n831));
  INV_X1    g645(.A(new_n371), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n831), .B1(new_n817), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n448), .B1(new_n805), .B2(new_n740), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n817), .A2(new_n832), .A3(new_n831), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n829), .A2(new_n830), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n826), .A2(new_n820), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n802), .A2(new_n806), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(KEYINPUT115), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(KEYINPUT115), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n838), .B1(new_n844), .B2(new_n827), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n675), .A2(new_n706), .A3(new_n743), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n747), .A2(new_n445), .ZN(new_n848));
  INV_X1    g662(.A(new_n730), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT101), .B1(new_n605), .B2(new_n626), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n650), .A2(new_n652), .A3(new_n673), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n848), .A2(new_n851), .A3(new_n632), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n684), .B2(new_n687), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n846), .B1(new_n847), .B2(new_n854), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n632), .A2(new_n848), .A3(new_n851), .A4(new_n852), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n683), .A2(KEYINPUT98), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n685), .A2(new_n686), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n446), .A2(new_n645), .A3(new_n653), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n660), .C1(new_n674), .C2(new_n705), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n859), .A2(KEYINPUT52), .A3(new_n743), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n855), .A2(KEYINPUT113), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT113), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n864), .B(new_n846), .C1(new_n847), .C2(new_n854), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n598), .A2(new_n655), .A3(new_n738), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n596), .B1(new_n606), .B2(new_n703), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n504), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n641), .A2(new_n870), .A3(new_n661), .A4(new_n733), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n654), .A2(new_n740), .A3(new_n722), .ZN(new_n872));
  INV_X1    g686(.A(new_n660), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n867), .A2(new_n868), .A3(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n748), .A2(new_n742), .A3(new_n737), .A4(new_n692), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n756), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT112), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n626), .A2(new_n673), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(new_n576), .A3(new_n624), .A4(new_n625), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n784), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n660), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n654), .A2(new_n661), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n860), .A2(KEYINPUT112), .A3(new_n660), .A4(new_n881), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n877), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n875), .A2(KEYINPUT53), .A3(new_n753), .A4(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT114), .B1(new_n866), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n884), .A2(new_n885), .ZN(new_n889));
  INV_X1    g703(.A(new_n877), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n753), .A3(new_n890), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n660), .A2(new_n724), .B1(new_n604), .B2(new_n870), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n603), .A2(new_n645), .A3(new_n653), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n731), .A2(new_n711), .A3(new_n504), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n893), .A2(new_n597), .B1(new_n804), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n371), .B(new_n712), .C1(new_n636), .C2(new_n616), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n892), .A2(new_n895), .A3(new_n598), .A4(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT53), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n891), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT114), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n865), .A4(new_n863), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n891), .A2(new_n897), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n855), .A2(new_n862), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n898), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n888), .A2(new_n901), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n902), .A2(new_n865), .A3(new_n863), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n898), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n898), .B2(new_n904), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n845), .B(new_n907), .C1(new_n906), .C2(new_n911), .ZN(new_n912));
  OR2_X1    g726(.A1(G952), .A2(G953), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR4_X1   g728(.A1(new_n775), .A2(new_n255), .A3(new_n758), .A4(new_n629), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT49), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n799), .B2(new_n916), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT109), .Z(new_n918));
  NAND2_X1  g732(.A1(new_n799), .A2(new_n916), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n919), .A2(KEYINPUT110), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n691), .B1(new_n919), .B2(KEYINPUT110), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n918), .A2(new_n821), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT111), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n914), .A2(new_n923), .ZN(G75));
  AOI21_X1  g738(.A(KEYINPUT53), .B1(new_n902), .B2(new_n903), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n866), .A2(new_n887), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n900), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n188), .B1(new_n927), .B2(new_n888), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT56), .B1(new_n928), .B2(new_n500), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n470), .A2(new_n484), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n482), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g747(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n934));
  NAND3_X1  g748(.A1(new_n888), .A2(new_n901), .A3(new_n905), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(G902), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n932), .B(new_n934), .C1(new_n936), .C2(new_n501), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n190), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n933), .A2(new_n940), .ZN(G51));
  XNOR2_X1  g755(.A(new_n746), .B(KEYINPUT121), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT57), .Z(new_n943));
  AOI21_X1  g757(.A(new_n906), .B1(new_n927), .B2(new_n888), .ZN(new_n944));
  INV_X1    g758(.A(new_n907), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n709), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n764), .B(KEYINPUT122), .Z(new_n949));
  NAND2_X1  g763(.A1(new_n928), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n938), .B1(new_n948), .B2(new_n950), .ZN(G54));
  AND2_X1   g765(.A1(KEYINPUT58), .A2(G475), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n935), .A2(G902), .A3(new_n590), .A4(new_n952), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(KEYINPUT123), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n935), .A2(G902), .A3(new_n952), .ZN(new_n955));
  INV_X1    g769(.A(new_n590), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n938), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(KEYINPUT123), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n954), .A2(new_n957), .A3(new_n958), .ZN(G60));
  NOR2_X1   g773(.A1(new_n944), .A2(new_n945), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n609), .A2(new_n611), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n613), .B(KEYINPUT59), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n939), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n907), .B1(new_n911), .B2(new_n906), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n961), .B1(new_n965), .B2(new_n962), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT60), .Z(new_n969));
  NAND2_X1  g783(.A1(new_n935), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n252), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n935), .A2(new_n643), .A3(new_n969), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(new_n939), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n971), .A2(KEYINPUT61), .A3(new_n939), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(G66));
  NAND2_X1  g791(.A1(new_n897), .A2(new_n190), .ZN(new_n978));
  OAI21_X1  g792(.A(G953), .B1(new_n453), .B2(new_n475), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n978), .A2(KEYINPUT124), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(KEYINPUT124), .B2(new_n978), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n930), .B1(G898), .B2(new_n190), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n981), .B(new_n982), .Z(G69));
  INV_X1    g797(.A(new_n663), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n770), .A2(new_n371), .A3(new_n632), .A4(new_n851), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n861), .A2(new_n743), .A3(new_n756), .ZN(new_n986));
  AND4_X1   g800(.A1(new_n753), .A2(new_n985), .A3(new_n782), .A4(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n987), .A2(new_n793), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n984), .B1(new_n988), .B2(G953), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n338), .A2(new_n339), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n584), .B(KEYINPUT125), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(G227), .A2(G900), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(G953), .ZN(new_n995));
  INV_X1    g809(.A(new_n992), .ZN(new_n996));
  INV_X1    g810(.A(new_n697), .ZN(new_n997));
  NOR4_X1   g811(.A1(new_n446), .A2(new_n784), .A3(new_n869), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n371), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(KEYINPUT126), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT126), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n998), .A2(new_n1001), .A3(new_n371), .ZN(new_n1002));
  AOI22_X1  g816(.A1(new_n770), .A2(new_n781), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n701), .ZN(new_n1004));
  OAI21_X1  g818(.A(KEYINPUT62), .B1(new_n1004), .B2(new_n847), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OR3_X1    g820(.A1(new_n1004), .A2(KEYINPUT62), .A3(new_n847), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1006), .A2(new_n793), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n996), .B1(new_n1008), .B2(G953), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n993), .A2(new_n995), .A3(new_n1009), .ZN(new_n1010));
  OAI211_X1 g824(.A(G953), .B(new_n994), .C1(new_n989), .C2(new_n996), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(G72));
  NAND4_X1  g826(.A1(new_n1006), .A2(new_n793), .A3(new_n875), .A4(new_n1007), .ZN(new_n1013));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n336), .B1(new_n340), .B2(new_n319), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n938), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n360), .A2(new_n336), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n341), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n910), .A2(new_n1015), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n987), .A2(new_n793), .A3(new_n875), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n1015), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n360), .A2(new_n335), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1018), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT127), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n1018), .A2(KEYINPUT127), .A3(new_n1025), .A4(new_n1021), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(G57));
endmodule


