

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755;

  NOR2_X1 U371 ( .A1(n754), .A2(n755), .ZN(n381) );
  XNOR2_X1 U372 ( .A(n498), .B(n462), .ZN(n486) );
  NOR2_X1 U373 ( .A1(n588), .A2(n675), .ZN(n589) );
  INV_X1 U374 ( .A(n587), .ZN(n675) );
  AND2_X1 U375 ( .A1(n395), .A2(n394), .ZN(n393) );
  XNOR2_X1 U376 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U377 ( .A(n439), .B(n438), .ZN(n557) );
  XNOR2_X1 U378 ( .A(n713), .B(n448), .ZN(n714) );
  XOR2_X1 U379 ( .A(G116), .B(G107), .Z(n500) );
  XNOR2_X1 U380 ( .A(n486), .B(n463), .ZN(n739) );
  XNOR2_X1 U381 ( .A(G137), .B(G134), .ZN(n463) );
  XNOR2_X1 U382 ( .A(n457), .B(G125), .ZN(n512) );
  XNOR2_X1 U383 ( .A(n504), .B(G478), .ZN(n558) );
  XNOR2_X1 U384 ( .A(n539), .B(KEYINPUT67), .ZN(n606) );
  OR2_X1 U385 ( .A1(n677), .A2(n678), .ZN(n539) );
  XNOR2_X1 U386 ( .A(n423), .B(n421), .ZN(n726) );
  XNOR2_X1 U387 ( .A(n483), .B(n422), .ZN(n421) );
  XNOR2_X1 U388 ( .A(n424), .B(n481), .ZN(n423) );
  XNOR2_X1 U389 ( .A(n567), .B(n367), .ZN(n366) );
  INV_X1 U390 ( .A(KEYINPUT101), .ZN(n367) );
  XNOR2_X1 U391 ( .A(n381), .B(KEYINPUT46), .ZN(n380) );
  AND2_X1 U392 ( .A1(n383), .A2(n614), .ZN(n382) );
  INV_X1 U393 ( .A(KEYINPUT48), .ZN(n434) );
  NAND2_X1 U394 ( .A1(n461), .A2(n460), .ZN(n498) );
  XNOR2_X1 U395 ( .A(n444), .B(G122), .ZN(n507) );
  INV_X1 U396 ( .A(G113), .ZN(n444) );
  XNOR2_X1 U397 ( .A(n512), .B(n416), .ZN(n527) );
  INV_X1 U398 ( .A(KEYINPUT10), .ZN(n416) );
  XOR2_X1 U399 ( .A(G131), .B(G140), .Z(n513) );
  INV_X1 U400 ( .A(KEYINPUT105), .ZN(n403) );
  AND2_X1 U401 ( .A1(n431), .A2(n430), .ZN(n604) );
  INV_X1 U402 ( .A(n581), .ZN(n430) );
  XNOR2_X1 U403 ( .A(n433), .B(n432), .ZN(n431) );
  INV_X1 U404 ( .A(KEYINPUT30), .ZN(n432) );
  XNOR2_X1 U405 ( .A(n515), .B(G475), .ZN(n438) );
  OR2_X1 U406 ( .A1(n713), .A2(G902), .ZN(n439) );
  OR2_X1 U407 ( .A1(n723), .A2(G902), .ZN(n414) );
  XNOR2_X1 U408 ( .A(n437), .B(n435), .ZN(n465) );
  XNOR2_X1 U409 ( .A(n436), .B(n482), .ZN(n435) );
  XNOR2_X1 U410 ( .A(n453), .B(n456), .ZN(n437) );
  XNOR2_X1 U411 ( .A(G119), .B(G110), .ZN(n528) );
  XOR2_X1 U412 ( .A(KEYINPUT23), .B(G140), .Z(n529) );
  XNOR2_X1 U413 ( .A(G137), .B(G128), .ZN(n449) );
  XNOR2_X1 U414 ( .A(n527), .B(n415), .ZN(n532) );
  XNOR2_X1 U415 ( .A(n526), .B(KEYINPUT88), .ZN(n415) );
  XNOR2_X1 U416 ( .A(KEYINPUT89), .B(KEYINPUT24), .ZN(n526) );
  XNOR2_X1 U417 ( .A(n509), .B(KEYINPUT12), .ZN(n445) );
  INV_X1 U418 ( .A(n507), .ZN(n443) );
  XOR2_X1 U419 ( .A(KEYINPUT95), .B(KEYINPUT11), .Z(n506) );
  XNOR2_X1 U420 ( .A(G143), .B(G104), .ZN(n505) );
  XNOR2_X1 U421 ( .A(G104), .B(KEYINPUT85), .ZN(n469) );
  XNOR2_X1 U422 ( .A(n598), .B(n399), .ZN(n696) );
  XNOR2_X1 U423 ( .A(n597), .B(n400), .ZN(n399) );
  NOR2_X1 U424 ( .A1(n667), .A2(n668), .ZN(n598) );
  INV_X1 U425 ( .A(KEYINPUT109), .ZN(n400) );
  NAND2_X1 U426 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U427 ( .A(n557), .B(n388), .ZN(n559) );
  INV_X1 U428 ( .A(KEYINPUT97), .ZN(n388) );
  NAND2_X1 U429 ( .A1(n606), .A2(n413), .ZN(n552) );
  INV_X1 U430 ( .A(n538), .ZN(n413) );
  XNOR2_X1 U431 ( .A(n411), .B(n474), .ZN(n602) );
  OR2_X1 U432 ( .A1(n708), .A2(G902), .ZN(n411) );
  XNOR2_X1 U433 ( .A(KEYINPUT22), .B(KEYINPUT74), .ZN(n521) );
  XNOR2_X1 U434 ( .A(n407), .B(n502), .ZN(n720) );
  XNOR2_X1 U435 ( .A(n501), .B(n408), .ZN(n407) );
  XNOR2_X1 U436 ( .A(n726), .B(n425), .ZN(n702) );
  XNOR2_X1 U437 ( .A(n492), .B(n426), .ZN(n425) );
  XNOR2_X1 U438 ( .A(n427), .B(n490), .ZN(n426) );
  NAND2_X1 U439 ( .A1(n360), .A2(G210), .ZN(n362) );
  AND2_X1 U440 ( .A1(n595), .A2(n649), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n620), .B(n596), .ZN(n663) );
  OR2_X1 U442 ( .A1(G237), .A2(G902), .ZN(n494) );
  XNOR2_X1 U443 ( .A(G116), .B(G131), .ZN(n454) );
  XNOR2_X1 U444 ( .A(KEYINPUT77), .B(KEYINPUT92), .ZN(n451) );
  XOR2_X1 U445 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n452) );
  XNOR2_X1 U446 ( .A(n450), .B(KEYINPUT93), .ZN(n436) );
  NOR2_X1 U447 ( .A1(G953), .A2(G237), .ZN(n508) );
  XNOR2_X1 U448 ( .A(KEYINPUT4), .B(KEYINPUT68), .ZN(n462) );
  XOR2_X1 U449 ( .A(KEYINPUT66), .B(G101), .Z(n485) );
  XOR2_X1 U450 ( .A(KEYINPUT3), .B(G119), .Z(n482) );
  XNOR2_X1 U451 ( .A(n507), .B(KEYINPUT16), .ZN(n424) );
  INV_X1 U452 ( .A(n500), .ZN(n422) );
  XNOR2_X1 U453 ( .A(n364), .B(n568), .ZN(n655) );
  INV_X1 U454 ( .A(KEYINPUT45), .ZN(n568) );
  NAND2_X1 U455 ( .A1(n551), .A2(KEYINPUT102), .ZN(n394) );
  INV_X1 U456 ( .A(KEYINPUT0), .ZN(n428) );
  NAND2_X1 U457 ( .A1(n389), .A2(n495), .ZN(n429) );
  NAND2_X1 U458 ( .A1(n625), .A2(n624), .ZN(n742) );
  XNOR2_X1 U459 ( .A(n499), .B(n409), .ZN(n408) );
  XNOR2_X1 U460 ( .A(n503), .B(n410), .ZN(n409) );
  INV_X1 U461 ( .A(KEYINPUT7), .ZN(n410) );
  XOR2_X1 U462 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n491) );
  XNOR2_X1 U463 ( .A(n543), .B(n542), .ZN(n695) );
  INV_X1 U464 ( .A(KEYINPUT39), .ZN(n607) );
  BUF_X1 U465 ( .A(n580), .Z(n620) );
  XNOR2_X1 U466 ( .A(n535), .B(n534), .ZN(n723) );
  XNOR2_X1 U467 ( .A(n530), .B(n449), .ZN(n531) );
  XNOR2_X1 U468 ( .A(n514), .B(n741), .ZN(n713) );
  XNOR2_X1 U469 ( .A(n445), .B(n443), .ZN(n510) );
  INV_X1 U470 ( .A(G475), .ZN(n361) );
  XNOR2_X1 U471 ( .A(n470), .B(n412), .ZN(n708) );
  XNOR2_X1 U472 ( .A(n473), .B(n481), .ZN(n412) );
  NAND2_X1 U473 ( .A1(n360), .A2(G469), .ZN(n359) );
  XNOR2_X1 U474 ( .A(KEYINPUT42), .B(n601), .ZN(n755) );
  XNOR2_X1 U475 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n404) );
  NAND2_X1 U476 ( .A1(n537), .A2(n576), .ZN(n371) );
  NOR2_X1 U477 ( .A1(n675), .A2(KEYINPUT65), .ZN(n441) );
  INV_X1 U478 ( .A(KEYINPUT99), .ZN(n386) );
  OR2_X1 U479 ( .A1(n560), .A2(n559), .ZN(n387) );
  INV_X1 U480 ( .A(n552), .ZN(n555) );
  INV_X1 U481 ( .A(n725), .ZN(n405) );
  XNOR2_X1 U482 ( .A(n629), .B(n354), .ZN(n406) );
  XNOR2_X1 U483 ( .A(n718), .B(n357), .ZN(n721) );
  XNOR2_X1 U484 ( .A(n720), .B(n719), .ZN(n357) );
  NOR2_X1 U485 ( .A1(n725), .A2(n705), .ZN(n706) );
  AND2_X1 U486 ( .A1(n662), .A2(n358), .ZN(n701) );
  NOR2_X1 U487 ( .A1(n700), .A2(G953), .ZN(n358) );
  XNOR2_X1 U488 ( .A(n414), .B(n350), .ZN(n677) );
  XOR2_X1 U489 ( .A(n384), .B(KEYINPUT36), .Z(n349) );
  XOR2_X1 U490 ( .A(n525), .B(n524), .Z(n350) );
  OR2_X1 U491 ( .A1(n587), .A2(n442), .ZN(n351) );
  OR2_X2 U492 ( .A1(n752), .A2(n398), .ZN(n352) );
  XNOR2_X1 U493 ( .A(n587), .B(KEYINPUT6), .ZN(n576) );
  NOR2_X1 U494 ( .A1(n603), .A2(n602), .ZN(n353) );
  INV_X1 U495 ( .A(G146), .ZN(n457) );
  INV_X1 U496 ( .A(n677), .ZN(n564) );
  XOR2_X1 U497 ( .A(n628), .B(KEYINPUT62), .Z(n354) );
  AND2_X1 U498 ( .A1(n550), .A2(KEYINPUT44), .ZN(n355) );
  INV_X1 U499 ( .A(KEYINPUT65), .ZN(n442) );
  INV_X1 U500 ( .A(KEYINPUT84), .ZN(n398) );
  XNOR2_X1 U501 ( .A(G902), .B(KEYINPUT15), .ZN(n626) );
  OR2_X1 U502 ( .A1(n626), .A2(n361), .ZN(n356) );
  NOR2_X2 U503 ( .A1(n725), .A2(n711), .ZN(n712) );
  NOR2_X2 U504 ( .A1(n725), .A2(n716), .ZN(n717) );
  OR2_X2 U505 ( .A1(n627), .A2(n362), .ZN(n704) );
  XNOR2_X1 U506 ( .A(n379), .B(n434), .ZN(n625) );
  NAND2_X1 U507 ( .A1(n587), .A2(n664), .ZN(n433) );
  XNOR2_X2 U508 ( .A(n653), .B(KEYINPUT2), .ZN(n627) );
  NOR2_X1 U509 ( .A1(n653), .A2(KEYINPUT81), .ZN(n654) );
  NOR2_X1 U510 ( .A1(n417), .A2(KEYINPUT84), .ZN(n376) );
  NOR2_X2 U511 ( .A1(n627), .A2(n626), .ZN(n363) );
  OR2_X1 U512 ( .A1(n627), .A2(n359), .ZN(n710) );
  INV_X1 U513 ( .A(n626), .ZN(n360) );
  OR2_X1 U514 ( .A1(n627), .A2(n356), .ZN(n715) );
  NAND2_X1 U515 ( .A1(n363), .A2(G478), .ZN(n718) );
  NAND2_X1 U516 ( .A1(n363), .A2(G472), .ZN(n629) );
  NAND2_X1 U517 ( .A1(n363), .A2(G217), .ZN(n722) );
  NAND2_X1 U518 ( .A1(n368), .A2(n365), .ZN(n364) );
  NOR2_X1 U519 ( .A1(n366), .A2(n355), .ZN(n365) );
  XNOR2_X1 U520 ( .A(n369), .B(n549), .ZN(n368) );
  NAND2_X1 U521 ( .A1(n372), .A2(n750), .ZN(n369) );
  XNOR2_X2 U522 ( .A(n370), .B(n404), .ZN(n752) );
  OR2_X2 U523 ( .A1(n536), .A2(n371), .ZN(n370) );
  XNOR2_X2 U524 ( .A(n522), .B(n521), .ZN(n536) );
  NAND2_X1 U525 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U526 ( .A1(n378), .A2(n377), .ZN(n373) );
  NAND2_X1 U527 ( .A1(n376), .A2(n375), .ZN(n374) );
  INV_X1 U528 ( .A(n419), .ZN(n375) );
  NAND2_X1 U529 ( .A1(n352), .A2(n397), .ZN(n377) );
  NAND2_X1 U530 ( .A1(n396), .A2(n397), .ZN(n378) );
  NAND2_X1 U531 ( .A1(n382), .A2(n380), .ZN(n379) );
  NAND2_X1 U532 ( .A1(n385), .A2(n579), .ZN(n384) );
  XNOR2_X1 U533 ( .A(n616), .B(KEYINPUT111), .ZN(n385) );
  NAND2_X1 U534 ( .A1(n401), .A2(n402), .ZN(n616) );
  XNOR2_X2 U535 ( .A(n387), .B(n386), .ZN(n643) );
  NAND2_X1 U536 ( .A1(n599), .A2(n389), .ZN(n591) );
  XNOR2_X2 U537 ( .A(n578), .B(KEYINPUT19), .ZN(n389) );
  NOR2_X1 U538 ( .A1(n536), .A2(n551), .ZN(n562) );
  NAND2_X1 U539 ( .A1(n393), .A2(n390), .ZN(n420) );
  NOR2_X1 U540 ( .A1(n551), .A2(KEYINPUT102), .ZN(n391) );
  INV_X1 U541 ( .A(n536), .ZN(n392) );
  NAND2_X1 U542 ( .A1(n536), .A2(KEYINPUT102), .ZN(n395) );
  NOR2_X1 U543 ( .A1(n417), .A2(n419), .ZN(n396) );
  NOR2_X1 U544 ( .A1(n419), .A2(n417), .ZN(n638) );
  NAND2_X1 U545 ( .A1(n752), .A2(n398), .ZN(n397) );
  NOR2_X1 U546 ( .A1(n564), .A2(n441), .ZN(n440) );
  INV_X1 U547 ( .A(n643), .ZN(n401) );
  XNOR2_X1 U548 ( .A(n577), .B(n403), .ZN(n402) );
  NAND2_X1 U549 ( .A1(n349), .A2(n551), .ZN(n649) );
  NOR2_X2 U550 ( .A1(n655), .A2(n742), .ZN(n653) );
  NAND2_X1 U551 ( .A1(n406), .A2(n405), .ZN(n630) );
  INV_X1 U552 ( .A(n606), .ZN(n684) );
  NAND2_X1 U553 ( .A1(n418), .A2(n440), .ZN(n417) );
  NAND2_X1 U554 ( .A1(n420), .A2(n442), .ZN(n418) );
  NOR2_X1 U555 ( .A1(n420), .A2(n351), .ZN(n419) );
  XNOR2_X1 U556 ( .A(n512), .B(n491), .ZN(n427) );
  INV_X1 U557 ( .A(n520), .ZN(n538) );
  XNOR2_X2 U558 ( .A(n429), .B(n428), .ZN(n520) );
  NAND2_X2 U559 ( .A1(n580), .A2(n664), .ZN(n578) );
  XNOR2_X2 U560 ( .A(n466), .B(n467), .ZN(n587) );
  XNOR2_X1 U561 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U562 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U563 ( .A(n704), .B(n703), .ZN(n705) );
  BUF_X1 U564 ( .A(n655), .Z(n730) );
  XNOR2_X1 U565 ( .A(n702), .B(n447), .ZN(n703) );
  AND2_X1 U566 ( .A1(G210), .A2(n494), .ZN(n446) );
  XNOR2_X1 U567 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n447) );
  XNOR2_X1 U568 ( .A(KEYINPUT59), .B(KEYINPUT119), .ZN(n448) );
  INV_X1 U569 ( .A(n578), .ZN(n579) );
  INV_X1 U570 ( .A(n652), .ZN(n623) );
  XNOR2_X1 U571 ( .A(n541), .B(KEYINPUT103), .ZN(n542) );
  AND2_X1 U572 ( .A1(n751), .A2(n623), .ZN(n624) );
  XNOR2_X1 U573 ( .A(n465), .B(n470), .ZN(n628) );
  INV_X1 U574 ( .A(n558), .ZN(n560) );
  XNOR2_X1 U575 ( .A(n608), .B(n607), .ZN(n622) );
  NOR2_X1 U576 ( .A1(n496), .A2(G952), .ZN(n725) );
  XNOR2_X1 U577 ( .A(n630), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U578 ( .A(G472), .B(KEYINPUT73), .ZN(n467) );
  NAND2_X1 U579 ( .A1(n508), .A2(G210), .ZN(n450) );
  XNOR2_X1 U580 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U581 ( .A(KEYINPUT78), .B(G113), .Z(n455) );
  XNOR2_X1 U582 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U583 ( .A(G146), .B(n485), .ZN(n464) );
  INV_X1 U584 ( .A(G128), .ZN(n458) );
  NAND2_X1 U585 ( .A1(G143), .A2(n458), .ZN(n461) );
  INV_X1 U586 ( .A(G143), .ZN(n459) );
  NAND2_X1 U587 ( .A1(n459), .A2(G128), .ZN(n460) );
  XNOR2_X1 U588 ( .A(n464), .B(n739), .ZN(n470) );
  NOR2_X1 U589 ( .A1(n628), .A2(G902), .ZN(n466) );
  XNOR2_X1 U590 ( .A(G469), .B(KEYINPUT70), .ZN(n468) );
  XNOR2_X1 U591 ( .A(n468), .B(KEYINPUT69), .ZN(n474) );
  XNOR2_X1 U592 ( .A(n469), .B(G110), .ZN(n481) );
  XOR2_X1 U593 ( .A(G107), .B(n513), .Z(n472) );
  XOR2_X2 U594 ( .A(KEYINPUT64), .B(G953), .Z(n496) );
  NAND2_X1 U595 ( .A1(G227), .A2(n496), .ZN(n471) );
  XNOR2_X1 U596 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U597 ( .A(n602), .B(KEYINPUT1), .ZN(n673) );
  INV_X1 U598 ( .A(n673), .ZN(n551) );
  NAND2_X1 U599 ( .A1(G234), .A2(G237), .ZN(n475) );
  XNOR2_X1 U600 ( .A(n475), .B(KEYINPUT14), .ZN(n476) );
  NAND2_X1 U601 ( .A1(G952), .A2(n476), .ZN(n694) );
  NOR2_X1 U602 ( .A1(G953), .A2(n694), .ZN(n574) );
  NAND2_X1 U603 ( .A1(G902), .A2(n476), .ZN(n569) );
  INV_X1 U604 ( .A(n569), .ZN(n477) );
  INV_X1 U605 ( .A(G953), .ZN(n661) );
  NOR2_X1 U606 ( .A1(G898), .A2(n661), .ZN(n728) );
  NAND2_X1 U607 ( .A1(n477), .A2(n728), .ZN(n478) );
  XOR2_X1 U608 ( .A(KEYINPUT86), .B(n478), .Z(n479) );
  NOR2_X1 U609 ( .A1(n574), .A2(n479), .ZN(n480) );
  XNOR2_X1 U610 ( .A(KEYINPUT87), .B(n480), .ZN(n495) );
  INV_X1 U611 ( .A(n482), .ZN(n483) );
  INV_X1 U612 ( .A(n486), .ZN(n484) );
  NAND2_X1 U613 ( .A1(n484), .A2(n485), .ZN(n489) );
  INV_X1 U614 ( .A(n485), .ZN(n487) );
  NAND2_X1 U615 ( .A1(n487), .A2(n486), .ZN(n488) );
  NAND2_X1 U616 ( .A1(n489), .A2(n488), .ZN(n492) );
  NAND2_X1 U617 ( .A1(G224), .A2(n496), .ZN(n490) );
  NAND2_X1 U618 ( .A1(n702), .A2(n626), .ZN(n493) );
  XNOR2_X2 U619 ( .A(n493), .B(n446), .ZN(n580) );
  NAND2_X1 U620 ( .A1(G214), .A2(n494), .ZN(n664) );
  NAND2_X1 U621 ( .A1(n496), .A2(G234), .ZN(n497) );
  XOR2_X1 U622 ( .A(KEYINPUT8), .B(n497), .Z(n533) );
  NAND2_X1 U623 ( .A1(G217), .A2(n533), .ZN(n502) );
  XNOR2_X1 U624 ( .A(G134), .B(n498), .ZN(n499) );
  XOR2_X1 U625 ( .A(n500), .B(G122), .Z(n501) );
  XNOR2_X1 U626 ( .A(KEYINPUT9), .B(KEYINPUT98), .ZN(n503) );
  NOR2_X1 U627 ( .A1(G902), .A2(n720), .ZN(n504) );
  XNOR2_X1 U628 ( .A(n506), .B(n505), .ZN(n511) );
  NAND2_X1 U629 ( .A1(G214), .A2(n508), .ZN(n509) );
  XNOR2_X1 U630 ( .A(n511), .B(n510), .ZN(n514) );
  XNOR2_X1 U631 ( .A(n513), .B(n527), .ZN(n741) );
  XNOR2_X1 U632 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n515) );
  NAND2_X1 U633 ( .A1(n558), .A2(n557), .ZN(n516) );
  XNOR2_X1 U634 ( .A(n516), .B(KEYINPUT100), .ZN(n667) );
  NAND2_X1 U635 ( .A1(G234), .A2(n626), .ZN(n517) );
  XNOR2_X1 U636 ( .A(KEYINPUT20), .B(n517), .ZN(n523) );
  NAND2_X1 U637 ( .A1(n523), .A2(G221), .ZN(n518) );
  XNOR2_X1 U638 ( .A(KEYINPUT21), .B(n518), .ZN(n678) );
  NOR2_X1 U639 ( .A1(n667), .A2(n678), .ZN(n519) );
  NAND2_X1 U640 ( .A1(n520), .A2(n519), .ZN(n522) );
  XOR2_X1 U641 ( .A(KEYINPUT25), .B(KEYINPUT90), .Z(n525) );
  NAND2_X1 U642 ( .A1(n523), .A2(G217), .ZN(n524) );
  XNOR2_X1 U643 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U644 ( .A(n532), .B(n531), .ZN(n535) );
  NAND2_X1 U645 ( .A1(G221), .A2(n533), .ZN(n534) );
  NOR2_X1 U646 ( .A1(n673), .A2(n564), .ZN(n537) );
  NOR2_X1 U647 ( .A1(n673), .A2(n576), .ZN(n540) );
  NAND2_X1 U648 ( .A1(n606), .A2(n540), .ZN(n543) );
  XOR2_X1 U649 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n541) );
  NOR2_X1 U650 ( .A1(n538), .A2(n695), .ZN(n544) );
  XNOR2_X1 U651 ( .A(n544), .B(KEYINPUT34), .ZN(n546) );
  OR2_X1 U652 ( .A1(n558), .A2(n557), .ZN(n586) );
  INV_X1 U653 ( .A(n586), .ZN(n545) );
  NAND2_X1 U654 ( .A1(n546), .A2(n545), .ZN(n548) );
  INV_X1 U655 ( .A(KEYINPUT35), .ZN(n547) );
  XNOR2_X1 U656 ( .A(n548), .B(n547), .ZN(n750) );
  INV_X1 U657 ( .A(KEYINPUT72), .ZN(n550) );
  NOR2_X1 U658 ( .A1(n550), .A2(KEYINPUT44), .ZN(n549) );
  NAND2_X1 U659 ( .A1(n551), .A2(n587), .ZN(n685) );
  NOR2_X1 U660 ( .A1(n685), .A2(n552), .ZN(n553) );
  XNOR2_X1 U661 ( .A(KEYINPUT31), .B(n553), .ZN(n645) );
  NOR2_X1 U662 ( .A1(n602), .A2(n587), .ZN(n554) );
  NAND2_X1 U663 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U664 ( .A(KEYINPUT94), .B(n556), .ZN(n635) );
  NAND2_X1 U665 ( .A1(n645), .A2(n635), .ZN(n561) );
  NAND2_X1 U666 ( .A1(n560), .A2(n559), .ZN(n646) );
  NAND2_X1 U667 ( .A1(n643), .A2(n646), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n561), .A2(n592), .ZN(n566) );
  NAND2_X1 U669 ( .A1(n562), .A2(n576), .ZN(n563) );
  XNOR2_X1 U670 ( .A(KEYINPUT83), .B(n563), .ZN(n565) );
  NAND2_X1 U671 ( .A1(n565), .A2(n564), .ZN(n631) );
  NAND2_X1 U672 ( .A1(n566), .A2(n631), .ZN(n567) );
  NOR2_X1 U673 ( .A1(G900), .A2(n569), .ZN(n571) );
  INV_X1 U674 ( .A(n496), .ZN(n570) );
  NAND2_X1 U675 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U676 ( .A(KEYINPUT104), .B(n572), .Z(n573) );
  NOR2_X1 U677 ( .A1(n574), .A2(n573), .ZN(n581) );
  NOR2_X1 U678 ( .A1(n581), .A2(n678), .ZN(n575) );
  NAND2_X1 U679 ( .A1(n575), .A2(n677), .ZN(n588) );
  NOR2_X1 U680 ( .A1(n588), .A2(n576), .ZN(n577) );
  NAND2_X1 U681 ( .A1(n606), .A2(n604), .ZN(n582) );
  NOR2_X1 U682 ( .A1(n602), .A2(n582), .ZN(n583) );
  AND2_X1 U683 ( .A1(n583), .A2(n620), .ZN(n584) );
  XOR2_X1 U684 ( .A(KEYINPUT108), .B(n584), .Z(n585) );
  NOR2_X1 U685 ( .A1(n586), .A2(n585), .ZN(n641) );
  XOR2_X1 U686 ( .A(n589), .B(KEYINPUT28), .Z(n590) );
  NOR2_X1 U687 ( .A1(n602), .A2(n590), .ZN(n599) );
  XNOR2_X1 U688 ( .A(n591), .B(KEYINPUT80), .ZN(n610) );
  INV_X1 U689 ( .A(n592), .ZN(n669) );
  NAND2_X1 U690 ( .A1(KEYINPUT75), .A2(n669), .ZN(n593) );
  NOR2_X1 U691 ( .A1(n610), .A2(n593), .ZN(n594) );
  NOR2_X1 U692 ( .A1(n641), .A2(n594), .ZN(n595) );
  XOR2_X1 U693 ( .A(KEYINPUT38), .B(KEYINPUT76), .Z(n596) );
  NAND2_X1 U694 ( .A1(n664), .A2(n663), .ZN(n668) );
  XNOR2_X1 U695 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n597) );
  INV_X1 U696 ( .A(n599), .ZN(n600) );
  NOR2_X1 U697 ( .A1(n696), .A2(n600), .ZN(n601) );
  INV_X1 U698 ( .A(n663), .ZN(n603) );
  AND2_X1 U699 ( .A1(n604), .A2(n353), .ZN(n605) );
  NAND2_X1 U700 ( .A1(n606), .A2(n605), .ZN(n608) );
  NOR2_X1 U701 ( .A1(n622), .A2(n643), .ZN(n609) );
  XNOR2_X1 U702 ( .A(n609), .B(KEYINPUT40), .ZN(n754) );
  INV_X1 U703 ( .A(KEYINPUT75), .ZN(n612) );
  NOR2_X1 U704 ( .A1(n610), .A2(n669), .ZN(n611) );
  NAND2_X1 U705 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U706 ( .A(KEYINPUT47), .B(n613), .Z(n614) );
  NAND2_X1 U707 ( .A1(n664), .A2(n673), .ZN(n615) );
  NOR2_X1 U708 ( .A1(n616), .A2(n615), .ZN(n618) );
  XNOR2_X1 U709 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n617) );
  XNOR2_X1 U710 ( .A(n618), .B(n617), .ZN(n619) );
  NOR2_X1 U711 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U712 ( .A(KEYINPUT107), .B(n621), .ZN(n751) );
  NOR2_X1 U713 ( .A1(n622), .A2(n646), .ZN(n652) );
  XNOR2_X1 U714 ( .A(G101), .B(n631), .ZN(G3) );
  NOR2_X1 U715 ( .A1(n635), .A2(n643), .ZN(n632) );
  XOR2_X1 U716 ( .A(G104), .B(n632), .Z(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n634) );
  XNOR2_X1 U718 ( .A(G107), .B(KEYINPUT27), .ZN(n633) );
  XNOR2_X1 U719 ( .A(n634), .B(n633), .ZN(n637) );
  NOR2_X1 U720 ( .A1(n635), .A2(n646), .ZN(n636) );
  XOR2_X1 U721 ( .A(n637), .B(n636), .Z(G9) );
  XOR2_X1 U722 ( .A(n638), .B(G110), .Z(G12) );
  NOR2_X1 U723 ( .A1(n610), .A2(n646), .ZN(n640) );
  XNOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .ZN(n639) );
  XNOR2_X1 U725 ( .A(n640), .B(n639), .ZN(G30) );
  XOR2_X1 U726 ( .A(n641), .B(G143), .Z(G45) );
  NOR2_X1 U727 ( .A1(n610), .A2(n643), .ZN(n642) );
  XOR2_X1 U728 ( .A(G146), .B(n642), .Z(G48) );
  NOR2_X1 U729 ( .A1(n643), .A2(n645), .ZN(n644) );
  XOR2_X1 U730 ( .A(G113), .B(n644), .Z(G15) );
  NOR2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n648) );
  XNOR2_X1 U732 ( .A(G116), .B(KEYINPUT113), .ZN(n647) );
  XNOR2_X1 U733 ( .A(n648), .B(n647), .ZN(G18) );
  INV_X1 U734 ( .A(n649), .ZN(n650) );
  XNOR2_X1 U735 ( .A(G125), .B(n650), .ZN(n651) );
  XNOR2_X1 U736 ( .A(n651), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U737 ( .A(G134), .B(n652), .Z(G36) );
  XNOR2_X1 U738 ( .A(n654), .B(KEYINPUT2), .ZN(n659) );
  INV_X1 U739 ( .A(n742), .ZN(n656) );
  NAND2_X1 U740 ( .A1(n656), .A2(n730), .ZN(n657) );
  NAND2_X1 U741 ( .A1(KEYINPUT81), .A2(n657), .ZN(n658) );
  NAND2_X1 U742 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U743 ( .A(n660), .B(KEYINPUT82), .ZN(n662) );
  NOR2_X1 U744 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U745 ( .A(n665), .B(KEYINPUT116), .ZN(n666) );
  NOR2_X1 U746 ( .A1(n667), .A2(n666), .ZN(n671) );
  NOR2_X1 U747 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U748 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U749 ( .A1(n672), .A2(n695), .ZN(n691) );
  NAND2_X1 U750 ( .A1(n673), .A2(n684), .ZN(n674) );
  XNOR2_X1 U751 ( .A(n674), .B(KEYINPUT50), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n676), .A2(n675), .ZN(n683) );
  XOR2_X1 U753 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n680) );
  NAND2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U755 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U756 ( .A(n681), .B(KEYINPUT114), .ZN(n682) );
  NOR2_X1 U757 ( .A1(n683), .A2(n682), .ZN(n687) );
  NOR2_X1 U758 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U759 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U760 ( .A(KEYINPUT51), .B(n688), .Z(n689) );
  NOR2_X1 U761 ( .A1(n696), .A2(n689), .ZN(n690) );
  NOR2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U763 ( .A(n692), .B(KEYINPUT52), .ZN(n693) );
  NOR2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n698) );
  NOR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U767 ( .A(n699), .B(KEYINPUT117), .ZN(n700) );
  XNOR2_X1 U768 ( .A(KEYINPUT53), .B(n701), .ZN(G75) );
  XNOR2_X1 U769 ( .A(KEYINPUT56), .B(n706), .ZN(G51) );
  XOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n707) );
  XNOR2_X1 U771 ( .A(KEYINPUT118), .B(n712), .ZN(G54) );
  XNOR2_X1 U772 ( .A(KEYINPUT60), .B(n717), .ZN(G60) );
  XOR2_X1 U773 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n719) );
  NOR2_X1 U774 ( .A1(n725), .A2(n721), .ZN(G63) );
  XNOR2_X1 U775 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U776 ( .A1(n725), .A2(n724), .ZN(G66) );
  XOR2_X1 U777 ( .A(n726), .B(G101), .Z(n727) );
  XNOR2_X1 U778 ( .A(KEYINPUT123), .B(n727), .ZN(n729) );
  NOR2_X1 U779 ( .A1(n729), .A2(n728), .ZN(n737) );
  OR2_X1 U780 ( .A1(G953), .A2(n730), .ZN(n734) );
  NAND2_X1 U781 ( .A1(G953), .A2(G224), .ZN(n731) );
  XNOR2_X1 U782 ( .A(KEYINPUT61), .B(n731), .ZN(n732) );
  NAND2_X1 U783 ( .A1(n732), .A2(G898), .ZN(n733) );
  NAND2_X1 U784 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U785 ( .A(n735), .B(KEYINPUT124), .ZN(n736) );
  XNOR2_X1 U786 ( .A(n737), .B(n736), .ZN(n738) );
  XNOR2_X1 U787 ( .A(KEYINPUT122), .B(n738), .ZN(G69) );
  XOR2_X1 U788 ( .A(n739), .B(KEYINPUT125), .Z(n740) );
  XOR2_X1 U789 ( .A(n741), .B(n740), .Z(n745) );
  XNOR2_X1 U790 ( .A(n742), .B(n745), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n743), .A2(n496), .ZN(n744) );
  XNOR2_X1 U792 ( .A(n744), .B(KEYINPUT126), .ZN(n749) );
  XNOR2_X1 U793 ( .A(G227), .B(n745), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U795 ( .A1(G953), .A2(n747), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(G72) );
  XNOR2_X1 U797 ( .A(G122), .B(n750), .ZN(G24) );
  XNOR2_X1 U798 ( .A(G140), .B(n751), .ZN(G42) );
  XNOR2_X1 U799 ( .A(G119), .B(KEYINPUT127), .ZN(n753) );
  XNOR2_X1 U800 ( .A(n753), .B(n752), .ZN(G21) );
  XOR2_X1 U801 ( .A(G131), .B(n754), .Z(G33) );
  XOR2_X1 U802 ( .A(G137), .B(n755), .Z(G39) );
endmodule

