//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(G137), .A3(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n469), .B1(new_n462), .B2(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n467), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n461), .A2(new_n462), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n475), .B1(new_n478), .B2(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT67), .B1(new_n479), .B2(new_n467), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  INV_X1    g056(.A(G125), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n482), .B1(new_n476), .B2(new_n477), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n481), .B(G2105), .C1(new_n483), .C2(new_n475), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n474), .B1(new_n480), .B2(new_n484), .ZN(G160));
  AOI21_X1  g060(.A(new_n467), .B1(new_n463), .B2(new_n465), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n463), .B2(new_n465), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  AND3_X1   g068(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(KEYINPUT3), .B1(new_n464), .B2(G2104), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n467), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n496), .A2(KEYINPUT4), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G126), .B(G2105), .C1(new_n494), .C2(new_n495), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(G114), .B2(new_n467), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n500), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  XOR2_X1   g089(.A(new_n514), .B(KEYINPUT71), .Z(new_n515));
  AOI21_X1  g090(.A(new_n507), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n516), .B1(new_n524), .B2(new_n525), .ZN(G166));
  INV_X1    g101(.A(new_n518), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  INV_X1    g103(.A(new_n520), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n528), .A2(new_n530), .A3(new_n531), .A4(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n509), .A2(new_n511), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(KEYINPUT72), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(G651), .A3(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(KEYINPUT73), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n527), .A2(G90), .B1(G52), .B2(new_n529), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(KEYINPUT73), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  AOI22_X1  g122(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT74), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n527), .A2(G81), .B1(G43), .B2(new_n529), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND3_X1  g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT75), .ZN(G176));
  XOR2_X1   g133(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n559));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(G188));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  INV_X1    g138(.A(G78), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n537), .A2(new_n563), .B1(new_n564), .B2(new_n508), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI221_X1 g142(.A(KEYINPUT77), .B1(new_n564), .B2(new_n508), .C1(new_n537), .C2(new_n563), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n567), .A2(G651), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n517), .A2(G53), .A3(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n527), .A2(G91), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n574));
  NOR2_X1   g149(.A1(G166), .A2(new_n574), .ZN(new_n575));
  AOI211_X1 g150(.A(KEYINPUT78), .B(new_n516), .C1(new_n524), .C2(new_n525), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n575), .A2(new_n576), .ZN(G303));
  NAND2_X1  g152(.A1(new_n527), .A2(G87), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n529), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  AOI22_X1  g156(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n507), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  INV_X1    g159(.A(G48), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n518), .A2(new_n584), .B1(new_n520), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n507), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT79), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n527), .A2(G85), .B1(G47), .B2(new_n529), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G290));
  AND3_X1   g168(.A1(new_n512), .A2(G92), .A3(new_n517), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT10), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n507), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n529), .A2(KEYINPUT80), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n529), .A2(KEYINPUT80), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n598), .A2(G54), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G171), .B2(new_n602), .ZN(G284));
  OAI21_X1  g179(.A(new_n603), .B1(G171), .B2(new_n602), .ZN(G321));
  NAND2_X1  g180(.A1(G299), .A2(new_n602), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n602), .B2(G168), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n602), .B2(G168), .ZN(G280));
  INV_X1    g183(.A(new_n601), .ZN(new_n609));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n552), .A2(new_n602), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n601), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n616));
  INV_X1    g191(.A(new_n486), .ZN(new_n617));
  INV_X1    g192(.A(G123), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  INV_X1    g195(.A(G111), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G2105), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n488), .B2(G135), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n486), .A2(KEYINPUT81), .A3(G123), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n619), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n472), .A2(new_n478), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n630), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT84), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT15), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2435), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(G2435), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT85), .Z(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n649), .A2(new_n651), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n642), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n654), .ZN(new_n656));
  INV_X1    g231(.A(new_n642), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n656), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n638), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n657), .B1(new_n656), .B2(new_n652), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n653), .A2(new_n654), .A3(new_n642), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n661), .A3(new_n637), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n662), .A3(G14), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n665), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n634), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n667), .A2(new_n668), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT18), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n678), .A3(new_n681), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n684), .B(new_n687), .C1(new_n678), .C2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT89), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n695), .B(new_n696), .Z(G229));
  NAND2_X1  g272(.A1(new_n609), .A2(G16), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G4), .B2(G16), .ZN(new_n699));
  INV_X1    g274(.A(G1348), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n486), .A2(G128), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n488), .A2(G140), .ZN(new_n704));
  OAI21_X1  g279(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n467), .A2(G116), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(KEYINPUT92), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(KEYINPUT92), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n712), .A2(G26), .ZN(new_n714));
  OAI21_X1  g289(.A(KEYINPUT28), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(KEYINPUT28), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n702), .B1(new_n717), .B2(G2067), .ZN(new_n718));
  INV_X1    g293(.A(G2067), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n715), .A2(new_n719), .A3(new_n716), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n699), .A2(new_n700), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G19), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n553), .B2(new_n722), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G1341), .Z(new_n725));
  NAND4_X1  g300(.A1(new_n718), .A2(new_n720), .A3(new_n721), .A4(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT93), .Z(new_n727));
  NAND3_X1  g302(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT25), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n488), .A2(G139), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n729), .B(new_n730), .C1(new_n467), .C2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT94), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G29), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G29), .B2(G33), .ZN(new_n735));
  INV_X1    g310(.A(G2072), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(G299), .A2(G16), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT98), .B(KEYINPUT23), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n722), .A2(G20), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G1956), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n627), .A2(G29), .A3(new_n628), .ZN(new_n745));
  NOR2_X1   g320(.A1(G29), .A2(G35), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G162), .B2(G29), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G2090), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n737), .A2(new_n744), .A3(new_n745), .A4(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(KEYINPUT24), .A2(G34), .ZN(new_n753));
  NAND2_X1  g328(.A1(KEYINPUT24), .A2(G34), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n753), .A2(new_n712), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G160), .B2(new_n712), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2084), .ZN(new_n757));
  OAI22_X1  g332(.A1(new_n735), .A2(new_n736), .B1(new_n750), .B2(new_n749), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n712), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n712), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT31), .B(G11), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT30), .B(G28), .Z(new_n764));
  OAI211_X1 g339(.A(new_n762), .B(new_n763), .C1(G29), .C2(new_n764), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n752), .A2(new_n757), .A3(new_n758), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n722), .A2(G22), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G166), .B2(new_n722), .ZN(new_n768));
  INV_X1    g343(.A(G1971), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G23), .ZN(new_n771));
  AND3_X1   g346(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT33), .B(G1976), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G6), .A2(G16), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n587), .B2(G16), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT32), .B(G1981), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n770), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT34), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n722), .A2(G24), .ZN(new_n782));
  INV_X1    g357(.A(G290), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n722), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1986), .ZN(new_n785));
  AND2_X1   g360(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n486), .A2(G119), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n488), .A2(G131), .ZN(new_n788));
  OAI21_X1  g363(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n467), .A2(G107), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n787), .B(new_n788), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G25), .B(new_n791), .S(G29), .Z(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT35), .B(G1991), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n781), .A2(new_n785), .A3(new_n786), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT91), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n795), .A2(new_n797), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n727), .B(new_n766), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G5), .B2(G16), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n801), .A2(G5), .A3(G16), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n802), .B(new_n803), .C1(G301), .C2(new_n722), .ZN(new_n804));
  INV_X1    g379(.A(G1961), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(G168), .A2(G16), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G16), .B2(G21), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT95), .B(G1966), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G29), .A2(G32), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n486), .A2(G129), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n488), .A2(G141), .ZN(new_n814));
  NAND3_X1  g389(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT26), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n472), .A2(G105), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n813), .A2(new_n814), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n812), .B1(new_n819), .B2(G29), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT27), .B(G1996), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n800), .A2(new_n806), .A3(new_n811), .A4(new_n822), .ZN(G311));
  INV_X1    g398(.A(G311), .ZN(G150));
  AOI22_X1  g399(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n507), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT100), .B(G55), .Z(new_n828));
  OAI22_X1  g403(.A1(new_n518), .A2(new_n827), .B1(new_n520), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n552), .B1(new_n834), .B2(new_n830), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n834), .B2(new_n830), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n552), .A2(KEYINPUT101), .A3(new_n831), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n601), .A2(new_n610), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT39), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n838), .B(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n833), .B1(new_n843), .B2(G860), .ZN(G145));
  XNOR2_X1  g419(.A(new_n629), .B(G162), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G160), .ZN(new_n846));
  INV_X1    g421(.A(new_n733), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n710), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n711), .A2(new_n733), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n819), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n818), .A3(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n499), .A2(new_n498), .ZN(new_n854));
  AOI211_X1 g429(.A(new_n497), .B(G2105), .C1(new_n463), .C2(new_n465), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT4), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n501), .A2(KEYINPUT102), .A3(new_n504), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT102), .B1(new_n501), .B2(new_n504), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  INV_X1    g437(.A(G126), .ZN(new_n863));
  AOI211_X1 g438(.A(new_n863), .B(new_n467), .C1(new_n463), .C2(new_n465), .ZN(new_n864));
  INV_X1    g439(.A(G114), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n502), .B1(new_n865), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n862), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n501), .A2(KEYINPUT102), .A3(new_n504), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n851), .A2(new_n857), .A3(new_n869), .A4(new_n852), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n861), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n488), .A2(G142), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT103), .Z(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n467), .A2(G118), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n486), .A2(new_n876), .A3(G130), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n486), .B2(G130), .ZN(new_n878));
  OAI221_X1 g453(.A(new_n873), .B1(new_n874), .B2(new_n875), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n632), .B(new_n791), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n879), .B(new_n880), .Z(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n871), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n861), .A2(new_n881), .A3(new_n870), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n846), .B1(new_n885), .B2(KEYINPUT105), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n885), .A2(new_n846), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g467(.A1(new_n836), .A2(new_n837), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n613), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n609), .B1(new_n895), .B2(G299), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n895), .B2(G299), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n601), .A2(new_n895), .A3(G299), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT41), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(KEYINPUT107), .A3(new_n902), .ZN(new_n903));
  OR3_X1    g478(.A1(new_n899), .A2(KEYINPUT107), .A3(KEYINPUT41), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n894), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n894), .A2(new_n899), .ZN(new_n906));
  XNOR2_X1  g481(.A(G166), .B(G288), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(G305), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n783), .ZN(new_n909));
  OR3_X1    g484(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n905), .B2(new_n906), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(G868), .B2(new_n830), .ZN(G295));
  OAI21_X1  g491(.A(new_n915), .B1(G868), .B2(new_n830), .ZN(G331));
  OAI21_X1  g492(.A(G171), .B1(KEYINPUT109), .B2(G286), .ZN(new_n918));
  AND2_X1   g493(.A1(G286), .A2(KEYINPUT109), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(G301), .A2(KEYINPUT109), .A3(G286), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n893), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n918), .A2(new_n919), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n838), .B1(new_n924), .B2(new_n921), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n926), .A2(new_n899), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n904), .A3(new_n903), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n909), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G37), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n909), .B1(new_n927), .B2(new_n928), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n909), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n900), .B(KEYINPUT111), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n902), .B(KEYINPUT110), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n935), .A2(new_n936), .B1(new_n923), .B2(new_n925), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n926), .A2(new_n899), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n939), .A2(new_n940), .A3(new_n930), .A4(new_n929), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n933), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n940), .B1(new_n931), .B2(new_n932), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n939), .A2(KEYINPUT43), .A3(new_n930), .A4(new_n929), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n944), .B1(new_n943), .B2(new_n947), .ZN(G397));
  NAND3_X1  g523(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n949));
  OAI21_X1  g524(.A(G8), .B1(new_n575), .B2(new_n576), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT55), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n860), .A2(KEYINPUT45), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G40), .ZN(new_n956));
  AOI211_X1 g531(.A(new_n956), .B(new_n474), .C1(new_n480), .C2(new_n484), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n954), .B1(new_n500), .B2(new_n505), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n955), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n769), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n860), .A2(new_n963), .A3(new_n954), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n958), .A2(KEYINPUT50), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n957), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n962), .B1(G2090), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n953), .A2(G8), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(G305), .A2(G1981), .ZN(new_n969));
  INV_X1    g544(.A(G1981), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n587), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n860), .A2(G160), .A3(G40), .A4(new_n954), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n975), .A2(G8), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n969), .A2(KEYINPUT49), .A3(new_n971), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n772), .A2(new_n979), .A3(G1976), .ZN(new_n980));
  INV_X1    g555(.A(G1976), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT114), .B1(G288), .B2(new_n981), .ZN(new_n982));
  AND4_X1   g557(.A1(G8), .A2(new_n980), .A3(new_n975), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n772), .A2(G1976), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT52), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(KEYINPUT115), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n983), .B(KEYINPUT115), .C1(KEYINPUT52), .C2(new_n984), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n978), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n968), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n963), .B1(new_n860), .B2(new_n954), .ZN(new_n992));
  NAND2_X1  g567(.A1(G160), .A2(G40), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n864), .A2(new_n866), .ZN(new_n995));
  AOI21_X1  g570(.A(G1384), .B1(new_n857), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n963), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n869), .B2(new_n857), .ZN(new_n998));
  OAI211_X1 g573(.A(KEYINPUT116), .B(new_n957), .C1(new_n998), .C2(new_n963), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n994), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n1000), .A2(G2090), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n962), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n953), .B1(new_n1002), .B2(G8), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n990), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1966), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT45), .B1(new_n860), .B2(new_n954), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT45), .B(new_n954), .C1(new_n500), .C2(new_n505), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(G40), .A3(G160), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G2084), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n964), .A2(new_n1011), .A3(new_n957), .A4(new_n965), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(G8), .A3(G286), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(G168), .A3(new_n1012), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(KEYINPUT120), .A3(G8), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT121), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(KEYINPUT51), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1015), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1014), .B(new_n1018), .C1(new_n1019), .C2(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n955), .A2(new_n957), .A3(new_n960), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT53), .B1(new_n1024), .B2(new_n761), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n805), .B2(new_n966), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n761), .A2(KEYINPUT53), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(G301), .B(KEYINPUT54), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1007), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n955), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1033), .A2(new_n474), .A3(new_n1028), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1034), .B(G40), .C1(new_n467), .C2(new_n479), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1030), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n1026), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1023), .A2(new_n1031), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT61), .ZN(new_n1039));
  XNOR2_X1  g614(.A(G299), .B(KEYINPUT57), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1000), .A2(new_n743), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT56), .B(G2072), .ZN(new_n1043));
  AND4_X1   g618(.A1(new_n957), .A2(new_n955), .A3(new_n960), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n1044), .B(new_n1040), .C1(new_n1000), .C2(new_n743), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1039), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1042), .A2(new_n1045), .A3(new_n1041), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1044), .B1(new_n1000), .B2(new_n743), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1040), .B(KEYINPUT118), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1049), .B(KEYINPUT61), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(KEYINPUT59), .ZN(new_n1054));
  INV_X1    g629(.A(G1996), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n955), .A2(new_n1055), .A3(new_n957), .A4(new_n960), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT58), .B(G1341), .Z(new_n1057));
  NAND2_X1  g632(.A1(new_n975), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1054), .B1(new_n1059), .B2(new_n553), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1054), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n552), .B(new_n1061), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1053), .A2(KEYINPUT59), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n975), .A2(G2067), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1065), .A2(new_n1066), .B1(new_n966), .B2(new_n700), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT117), .B1(new_n975), .B2(G2067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(KEYINPUT60), .A3(new_n609), .A4(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n860), .A2(new_n963), .A3(new_n954), .ZN(new_n1070));
  OAI211_X1 g645(.A(G40), .B(G160), .C1(new_n996), .C2(new_n963), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n700), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n998), .A2(new_n957), .A3(new_n1065), .A4(new_n719), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT60), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n601), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1072), .A2(new_n1068), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n609), .A2(KEYINPUT60), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1063), .A2(new_n1064), .B1(new_n1069), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1048), .A2(new_n1052), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n601), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(new_n1049), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1038), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n967), .A2(G8), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(new_n949), .A3(new_n952), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n968), .A2(new_n989), .A3(KEYINPUT63), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1013), .A2(G8), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(G286), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1005), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1090), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT63), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n989), .A2(G8), .A3(new_n953), .A4(new_n967), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n978), .A2(G1976), .A3(G288), .ZN(new_n1096));
  INV_X1    g671(.A(new_n971), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n976), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT122), .B1(new_n1092), .B2(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1094), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1038), .A2(new_n1084), .B1(new_n1090), .B2(new_n1088), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1101), .B(new_n1102), .C1(new_n1103), .C2(new_n1005), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1023), .A2(KEYINPUT62), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT123), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1023), .A2(new_n1107), .A3(KEYINPUT62), .ZN(new_n1108));
  AOI21_X1  g683(.A(G301), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1023), .A2(KEYINPUT62), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1109), .A2(new_n1004), .A3(new_n1029), .A4(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1100), .A2(new_n1104), .A3(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n710), .B(G2067), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1032), .A2(new_n993), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(new_n1115), .B(KEYINPUT113), .Z(new_n1116));
  INV_X1    g691(.A(new_n1114), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n818), .B(new_n1055), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n791), .B(new_n793), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G1986), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n783), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT112), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1123), .B2(new_n783), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1122), .B1(new_n1114), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1112), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n791), .A2(new_n793), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1119), .A2(new_n1130), .B1(G2067), .B2(new_n710), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1131), .A2(KEYINPUT124), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(KEYINPUT124), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1114), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1125), .A2(new_n1117), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1135), .B(KEYINPUT48), .Z(new_n1136));
  NAND2_X1  g711(.A1(new_n1121), .A2(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1113), .A2(new_n818), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT46), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1138), .A2(new_n1114), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI22_X1  g716(.A1(new_n1117), .A2(G1996), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1114), .A2(KEYINPUT125), .A3(KEYINPUT46), .A4(new_n1055), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1145));
  XNOR2_X1  g720(.A(new_n1144), .B(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1134), .A2(new_n1137), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1128), .A2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g723(.A(G229), .ZN(new_n1150));
  OR2_X1    g724(.A1(G227), .A2(new_n459), .ZN(new_n1151));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n1152));
  OR2_X1    g726(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g727(.A1(new_n663), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g728(.A(new_n1154), .B1(new_n889), .B2(new_n890), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1156));
  AND4_X1   g730(.A1(new_n1150), .A2(new_n1155), .A3(new_n942), .A4(new_n1156), .ZN(G308));
  NAND4_X1  g731(.A1(new_n1155), .A2(new_n942), .A3(new_n1150), .A4(new_n1156), .ZN(G225));
endmodule


