//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1227, new_n1228,
    new_n1229, new_n1230;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n451), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G113), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(new_n462), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n467), .B2(G125), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT69), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n462), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n475), .B1(new_n465), .B2(new_n466), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n474), .B(G2105), .C1(new_n476), .C2(new_n463), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n470), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n471), .A2(G136), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n469), .B1(new_n465), .B2(new_n466), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  MUX2_X1   g057(.A(G100), .B(G112), .S(G2105), .Z(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2104), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(G162));
  INV_X1    g060(.A(G126), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n465), .B2(new_n466), .ZN(new_n487));
  AND2_X1   g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  OAI21_X1  g063(.A(G2105), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(KEYINPUT4), .A2(G138), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n465), .B2(new_n466), .ZN(new_n491));
  NAND2_X1  g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n469), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n469), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n489), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI211_X1 g078(.A(G50), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  XNOR2_X1  g080(.A(new_n504), .B(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(KEYINPUT5), .B1(KEYINPUT71), .B2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n509), .A2(new_n510), .B1(new_n503), .B2(new_n502), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n506), .A2(new_n514), .A3(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND2_X1  g094(.A1(KEYINPUT71), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(new_n508), .ZN(new_n523));
  AND2_X1   g098(.A1(G63), .A2(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n502), .A2(new_n503), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n502), .A2(new_n503), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(G89), .A3(new_n523), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n523), .A2(KEYINPUT72), .A3(new_n524), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n527), .A2(new_n531), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT73), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT7), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n535), .A2(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(new_n532), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT74), .B(G90), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n541), .A2(new_n542), .B1(new_n515), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n523), .A2(G64), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n544), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n545), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n532), .A2(G81), .A3(new_n523), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  OAI211_X1 g128(.A(G43), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n551), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT77), .ZN(new_n564));
  XOR2_X1   g139(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(G188));
  INV_X1    g142(.A(G78), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT78), .B1(new_n568), .B2(new_n529), .ZN(new_n569));
  OR3_X1    g144(.A1(new_n568), .A2(new_n529), .A3(KEYINPUT78), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n569), .B(new_n570), .C1(new_n511), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  OAI211_X1 g148(.A(G53), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n516), .A2(G91), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  NAND2_X1  g154(.A1(new_n516), .A2(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n530), .A2(G49), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n515), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n532), .A2(new_n523), .A3(KEYINPUT79), .A4(G86), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g163(.A(G48), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(G61), .B1(new_n509), .B2(new_n510), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n590), .B1(new_n593), .B2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT80), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n588), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G305));
  AOI22_X1  g175(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(new_n545), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n530), .A2(G47), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n532), .A2(G85), .A3(new_n523), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n605), .B1(new_n603), .B2(new_n604), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n602), .B1(new_n607), .B2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n511), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n515), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n532), .A2(new_n523), .A3(G92), .A4(new_n614), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  MUX2_X1   g195(.A(new_n620), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g196(.A(new_n620), .B(G301), .S(G868), .Z(G321));
  NOR2_X1   g197(.A1(G299), .A2(G868), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(G868), .B2(G168), .ZN(G297));
  XNOR2_X1  g199(.A(G297), .B(KEYINPUT83), .ZN(G280));
  INV_X1    g200(.A(new_n620), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND3_X1  g203(.A1(new_n626), .A2(KEYINPUT84), .A3(new_n627), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n620), .B2(G559), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g210(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n469), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT13), .Z(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  MUX2_X1   g217(.A(G99), .B(G111), .S(G2105), .Z(new_n643));
  AOI22_X1  g218(.A1(G123), .A2(new_n481), .B1(new_n643), .B2(G2104), .ZN(new_n644));
  INV_X1    g219(.A(G135), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n467), .A2(new_n469), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2096), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n641), .A2(new_n642), .A3(new_n648), .ZN(G156));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  INV_X1    g225(.A(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n652), .A2(G2427), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(G2427), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(G2430), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(G2430), .A3(new_n654), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n663), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT86), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n670));
  NAND4_X1  g245(.A1(new_n664), .A2(new_n670), .A3(new_n665), .A4(new_n667), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(G14), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n664), .A2(new_n665), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n673), .B1(new_n674), .B2(new_n666), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G401));
  XNOR2_X1  g252(.A(G2067), .B(G2678), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2072), .B(G2078), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  OR3_X1    g256(.A1(new_n680), .A2(KEYINPUT87), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(KEYINPUT87), .B1(new_n680), .B2(new_n681), .ZN(new_n683));
  INV_X1    g258(.A(new_n678), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n679), .B(KEYINPUT17), .Z(new_n685));
  OAI211_X1 g260(.A(new_n682), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n685), .A2(new_n684), .A3(new_n681), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n681), .A2(new_n678), .A3(new_n679), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT18), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G2096), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT88), .B(G2100), .Z(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G227));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT19), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1956), .B(G2474), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT89), .ZN(new_n701));
  XOR2_X1   g276(.A(G1961), .B(G1966), .Z(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT20), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n701), .A2(new_n702), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(new_n698), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(new_n705), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n704), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n709), .A2(new_n711), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(G1991), .B(G1996), .Z(new_n715));
  XNOR2_X1  g290(.A(G1981), .B(G1986), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n715), .B(new_n716), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n717), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n712), .B2(new_n713), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(G229));
  NAND2_X1  g297(.A1(new_n626), .A2(G16), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G4), .B2(G16), .ZN(new_n724));
  INV_X1    g299(.A(G1348), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G5), .A2(G16), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT99), .Z(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G171), .B2(G16), .ZN(new_n729));
  INV_X1    g304(.A(G1961), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n724), .A2(new_n725), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  AND2_X1   g308(.A1(KEYINPUT24), .A2(G34), .ZN(new_n734));
  NOR2_X1   g309(.A1(KEYINPUT24), .A2(G34), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n478), .B2(new_n733), .ZN(new_n737));
  INV_X1    g312(.A(G2084), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n726), .A2(new_n731), .A3(new_n732), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n733), .A2(G35), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT101), .Z(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n733), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT102), .B(KEYINPUT29), .Z(new_n744));
  XOR2_X1   g319(.A(new_n743), .B(new_n744), .Z(new_n745));
  INV_X1    g320(.A(G2090), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT31), .B(G11), .Z(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT30), .B(G28), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n733), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n733), .A2(G32), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT26), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n471), .A2(G141), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n481), .A2(G129), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n472), .A2(G105), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n753), .A2(new_n754), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n751), .B1(new_n757), .B2(G29), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n750), .B1(new_n733), .B2(new_n647), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n758), .B2(new_n759), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n733), .A2(G26), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT28), .ZN(new_n763));
  OAI211_X1 g338(.A(G140), .B(new_n469), .C1(new_n495), .C2(new_n496), .ZN(new_n764));
  OAI211_X1 g339(.A(G128), .B(G2105), .C1(new_n495), .C2(new_n496), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(G2104), .B1(new_n469), .B2(G116), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G104), .B2(G2105), .ZN(new_n769));
  INV_X1    g344(.A(G104), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n770), .A2(new_n469), .A3(KEYINPUT95), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n767), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n766), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n763), .B1(new_n773), .B2(new_n733), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT96), .B(G2067), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G27), .A2(G29), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G164), .B2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G2078), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n747), .A2(new_n761), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n740), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n467), .A2(G127), .ZN(new_n783));
  NAND2_X1  g358(.A1(G115), .A2(G2104), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n469), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT97), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n469), .A2(G2104), .ZN(new_n789));
  INV_X1    g364(.A(G103), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n791), .A2(new_n792), .B1(new_n471), .B2(G139), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n786), .A2(new_n787), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n787), .B1(new_n786), .B2(new_n793), .ZN(new_n796));
  OAI21_X1  g371(.A(G29), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G33), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(G29), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G2072), .Z(new_n800));
  NOR2_X1   g375(.A1(new_n745), .A2(new_n746), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT103), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G16), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G20), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT23), .Z(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G299), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1956), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n782), .A2(new_n800), .A3(new_n803), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G19), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n559), .B2(G16), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1341), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n737), .A2(new_n738), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT100), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(G16), .A2(G21), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G168), .B2(G16), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT98), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1966), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n809), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT104), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(KEYINPUT104), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT32), .B(G1981), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n599), .A2(G16), .ZN(new_n826));
  OR2_X1    g401(.A1(G6), .A2(G16), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n826), .A2(KEYINPUT93), .A3(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(KEYINPUT93), .B1(new_n826), .B2(new_n827), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n825), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n830), .ZN(new_n832));
  INV_X1    g407(.A(new_n825), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n832), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT34), .ZN(new_n836));
  NOR2_X1   g411(.A1(G16), .A2(G22), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G166), .B2(G16), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G1971), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n804), .A2(G23), .ZN(new_n840));
  INV_X1    g415(.A(G288), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n841), .B2(new_n804), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT33), .B(G1976), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n835), .A2(new_n836), .A3(new_n845), .ZN(new_n846));
  MUX2_X1   g421(.A(G24), .B(G290), .S(G16), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G1986), .ZN(new_n848));
  NOR2_X1   g423(.A1(G25), .A2(G29), .ZN(new_n849));
  OAI211_X1 g424(.A(G131), .B(new_n469), .C1(new_n495), .C2(new_n496), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT91), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n467), .A2(KEYINPUT91), .A3(G131), .A4(new_n469), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT92), .ZN(new_n855));
  MUX2_X1   g430(.A(G95), .B(G107), .S(G2105), .Z(new_n856));
  AOI22_X1  g431(.A1(G119), .A2(new_n481), .B1(new_n856), .B2(G2104), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n855), .B1(new_n854), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n849), .B1(new_n860), .B2(G29), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G1991), .Z(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n861), .B(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n848), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n846), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n836), .B1(new_n835), .B2(new_n845), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n823), .B(new_n824), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n867), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n823), .A2(new_n824), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n869), .A2(new_n846), .A3(new_n865), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n821), .A2(new_n822), .B1(new_n872), .B2(new_n873), .ZN(G311));
  NAND2_X1  g449(.A1(new_n822), .A2(new_n821), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n873), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(G150));
  INV_X1    g452(.A(G55), .ZN(new_n878));
  INV_X1    g453(.A(G93), .ZN(new_n879));
  OAI22_X1  g454(.A1(new_n541), .A2(new_n878), .B1(new_n515), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n523), .A2(G67), .ZN(new_n881));
  NAND2_X1  g456(.A1(G80), .A2(G543), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n545), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G860), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT37), .ZN(new_n887));
  INV_X1    g462(.A(new_n884), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n558), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n884), .B(new_n551), .C1(new_n557), .C2(new_n556), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT38), .Z(new_n892));
  NOR2_X1   g467(.A1(new_n620), .A2(new_n627), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT105), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n892), .B(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n896), .A2(KEYINPUT39), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n885), .B1(new_n896), .B2(KEYINPUT39), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n887), .B1(new_n897), .B2(new_n898), .ZN(G145));
  INV_X1    g474(.A(new_n757), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n495), .A2(new_n496), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n492), .B1(new_n901), .B2(new_n490), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n902), .A2(new_n469), .B1(new_n498), .B2(new_n497), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n773), .B1(new_n903), .B2(new_n489), .ZN(new_n904));
  INV_X1    g479(.A(new_n772), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(new_n764), .A3(new_n765), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n500), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n900), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n500), .A2(new_n906), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n903), .A2(new_n773), .A3(new_n489), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n910), .A3(new_n757), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n791), .A2(new_n792), .ZN(new_n912));
  INV_X1    g487(.A(G139), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(new_n646), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT106), .B1(new_n914), .B2(new_n785), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n908), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  OAI211_X1 g491(.A(KEYINPUT97), .B(KEYINPUT106), .C1(new_n914), .C2(new_n785), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n917), .A2(new_n794), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n908), .B2(new_n911), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n471), .A2(G142), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n481), .A2(G130), .ZN(new_n921));
  MUX2_X1   g496(.A(G106), .B(G118), .S(G2105), .Z(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(G2104), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n858), .B2(new_n859), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n854), .A2(new_n857), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT92), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n854), .A2(new_n857), .A3(new_n855), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n924), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n638), .B(KEYINPUT107), .Z(new_n931));
  AND3_X1   g506(.A1(new_n926), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n926), .B2(new_n930), .ZN(new_n933));
  OAI22_X1  g508(.A1(new_n916), .A2(new_n919), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(G160), .A2(G162), .ZN(new_n935));
  INV_X1    g510(.A(G162), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n478), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n935), .A2(new_n647), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n647), .B1(new_n935), .B2(new_n937), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n926), .A2(new_n930), .ZN(new_n941));
  INV_X1    g516(.A(new_n931), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n917), .A2(new_n794), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n909), .A2(new_n910), .A3(new_n757), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n757), .B1(new_n909), .B2(new_n910), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n908), .A2(new_n911), .A3(new_n915), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n926), .A2(new_n930), .A3(new_n931), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n943), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n934), .A2(new_n940), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G37), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n934), .A2(new_n950), .ZN(new_n955));
  INV_X1    g530(.A(new_n940), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI211_X1 g532(.A(KEYINPUT108), .B(new_n940), .C1(new_n934), .C2(new_n950), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n953), .B(KEYINPUT109), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g539(.A1(new_n888), .A2(G868), .ZN(new_n965));
  AOI21_X1  g540(.A(G303), .B1(new_n596), .B2(new_n598), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(G290), .A2(G288), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n841), .B(new_n602), .C1(new_n608), .C2(new_n607), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n596), .A2(G303), .A3(new_n598), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n967), .A2(new_n968), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n969), .ZN(new_n972));
  INV_X1    g547(.A(new_n970), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(new_n966), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n632), .B(new_n891), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n620), .A2(G299), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n572), .A2(G651), .B1(new_n516), .B2(G91), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n978), .A2(new_n613), .A3(new_n575), .A4(new_n619), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n976), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT110), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT41), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n977), .B2(new_n979), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n977), .A2(new_n984), .A3(new_n979), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n985), .B1(KEYINPUT111), .B2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n980), .A2(KEYINPUT111), .A3(KEYINPUT41), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n976), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n976), .A2(new_n991), .A3(new_n981), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n983), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT42), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(KEYINPUT42), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n975), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n996), .ZN(new_n998));
  INV_X1    g573(.A(new_n975), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n994), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n965), .B1(new_n1001), .B2(G868), .ZN(G295));
  AOI21_X1  g577(.A(new_n965), .B1(new_n1001), .B2(G868), .ZN(G331));
  NAND2_X1  g578(.A1(G168), .A2(G171), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n535), .A2(new_n539), .B1(new_n548), .B2(new_n544), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n891), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n889), .A2(new_n1004), .A3(new_n890), .A4(new_n1005), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n987), .B2(new_n988), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n981), .A3(new_n1008), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n975), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n952), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n975), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n985), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n986), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1009), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n1011), .ZN(new_n1020));
  AOI21_X1  g595(.A(G37), .B1(new_n1020), .B2(new_n999), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT43), .B1(new_n1021), .B2(new_n1012), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(KEYINPUT44), .ZN(new_n1024));
  OR3_X1    g599(.A1(new_n1013), .A2(KEYINPUT43), .A3(new_n1015), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1021), .A2(new_n1012), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT112), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1027), .B2(new_n1014), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1024), .B1(new_n1028), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g604(.A(KEYINPUT49), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n588), .A2(new_n594), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n516), .A2(G86), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n594), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1030), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT118), .B(G8), .Z(new_n1036));
  NAND4_X1  g611(.A1(new_n470), .A2(G40), .A3(new_n473), .A4(new_n477), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1384), .B1(new_n903), .B2(new_n489), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n588), .A2(new_n594), .A3(new_n1031), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n594), .A2(new_n1033), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT49), .B(new_n1041), .C1(new_n1042), .C2(new_n1031), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1035), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n580), .A2(G1976), .A3(new_n581), .A4(new_n582), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1040), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1036), .ZN(new_n1049));
  INV_X1    g624(.A(G1384), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n500), .A2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1049), .B(new_n1045), .C1(new_n1037), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT52), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1044), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(KEYINPUT117), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(KEYINPUT117), .B2(new_n1055), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n500), .A2(KEYINPUT50), .A3(new_n1050), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT50), .B1(new_n500), .B2(new_n1050), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n746), .B(new_n1038), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT115), .B(G1971), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT45), .B1(new_n500), .B2(new_n1050), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(new_n1037), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT113), .B(G1384), .Z(new_n1067));
  NAND3_X1  g642(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1064), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1049), .B1(new_n1063), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1054), .B1(new_n1059), .B2(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1069), .A2(KEYINPUT116), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1062), .B1(new_n1069), .B2(KEYINPUT116), .ZN(new_n1073));
  OAI211_X1 g648(.A(G8), .B(new_n1058), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT45), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1051), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1077), .A2(new_n1038), .A3(new_n779), .A4(new_n1068), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1038), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n730), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1039), .A2(KEYINPUT45), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1066), .A2(KEYINPUT53), .A3(new_n779), .A4(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G171), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1075), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n738), .B(new_n1038), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(G1966), .B1(new_n1066), .B2(new_n1083), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1051), .A2(new_n1076), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1093), .A2(new_n1065), .A3(new_n1037), .ZN(new_n1094));
  OAI211_X1 g669(.A(KEYINPUT123), .B(new_n1089), .C1(new_n1094), .C2(G1966), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1092), .A2(G8), .A3(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G168), .A2(new_n1036), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1092), .A2(new_n1097), .A3(new_n1095), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(KEYINPUT51), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(new_n1036), .ZN(new_n1104));
  OR3_X1    g679(.A1(new_n1104), .A2(KEYINPUT51), .A3(new_n1097), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1102), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1087), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1101), .A2(new_n1109), .A3(new_n1105), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n500), .A2(new_n1067), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1076), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n473), .A2(KEYINPUT53), .A3(G40), .A4(new_n779), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n468), .A2(new_n469), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1115), .A3(new_n1068), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1080), .A2(new_n1082), .A3(G301), .A4(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT54), .B1(new_n1086), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g695(.A(KEYINPUT124), .B(KEYINPUT54), .C1(new_n1086), .C2(new_n1117), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .A4(G301), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT54), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1080), .A2(new_n1082), .A3(new_n1124), .A4(new_n1116), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(G171), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1080), .A2(new_n1082), .A3(new_n1116), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT125), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1123), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1120), .A2(new_n1121), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1956), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1081), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT56), .B(G2072), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1066), .A2(new_n1068), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n1135));
  XNOR2_X1  g710(.A(G299), .B(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1081), .A2(new_n725), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1037), .A2(new_n1051), .ZN(new_n1139));
  INV_X1    g714(.A(G2067), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n620), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1136), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1137), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(new_n626), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT60), .B1(new_n1149), .B2(new_n1142), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1077), .A2(new_n1038), .A3(new_n1068), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT58), .B(G1341), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1151), .A2(G1996), .B1(new_n1139), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n559), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(KEYINPUT122), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1153), .B(new_n559), .C1(KEYINPUT122), .C2(new_n1155), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1143), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1160), .A2(KEYINPUT61), .A3(new_n1137), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1150), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  OR3_X1    g737(.A1(new_n1148), .A2(KEYINPUT60), .A3(new_n620), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1137), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(new_n1143), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1163), .B1(new_n1165), .B2(KEYINPUT61), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1146), .B(new_n1147), .C1(new_n1162), .C2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1110), .A2(new_n1130), .A3(new_n1167), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1044), .A2(new_n1046), .A3(new_n841), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1041), .B(KEYINPUT120), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1040), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1054), .B(KEYINPUT119), .Z(new_n1172));
  OAI21_X1  g747(.A(new_n1171), .B1(new_n1172), .B2(new_n1074), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1104), .A2(G168), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(G8), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1059), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1054), .B(KEYINPUT119), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1176), .A2(new_n1074), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1175), .B1(new_n1075), .B2(new_n1174), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1173), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1108), .A2(new_n1168), .A3(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1112), .A2(new_n1037), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1184), .A2(KEYINPUT114), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(KEYINPUT114), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n757), .B(G1996), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n906), .A2(G2067), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n773), .A2(new_n1140), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n863), .B1(new_n858), .B2(new_n859), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n860), .A2(new_n862), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(G290), .B(G1986), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1188), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1183), .A2(new_n1198), .ZN(new_n1199));
  OR3_X1    g774(.A1(new_n1187), .A2(G1986), .A3(G290), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT48), .ZN(new_n1201));
  OR2_X1    g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1188), .A2(new_n1196), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1187), .A2(new_n1193), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1191), .B1(new_n1206), .B2(new_n1195), .ZN(new_n1207));
  AND2_X1   g782(.A1(new_n1207), .A2(KEYINPUT126), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1188), .B1(new_n1207), .B2(KEYINPUT126), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1205), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1187), .A2(G1996), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT46), .Z(new_n1212));
  OAI21_X1  g787(.A(new_n1188), .B1(new_n757), .B2(new_n1192), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1214), .A2(KEYINPUT47), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1214), .A2(KEYINPUT47), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1210), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1199), .A2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g793(.A(new_n459), .B1(new_n693), .B2(new_n694), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n676), .A2(new_n721), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g795(.A(new_n1221), .ZN(new_n1222));
  AND4_X1   g796(.A1(KEYINPUT127), .A2(new_n963), .A3(new_n1023), .A4(new_n1222), .ZN(new_n1223));
  AOI21_X1  g797(.A(new_n1221), .B1(new_n961), .B2(new_n962), .ZN(new_n1224));
  AOI21_X1  g798(.A(KEYINPUT127), .B1(new_n1224), .B2(new_n1023), .ZN(new_n1225));
  NOR2_X1   g799(.A1(new_n1223), .A2(new_n1225), .ZN(G308));
  NAND3_X1  g800(.A1(new_n963), .A2(new_n1023), .A3(new_n1222), .ZN(new_n1227));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n1228));
  NAND2_X1  g802(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g803(.A1(new_n1224), .A2(KEYINPUT127), .A3(new_n1023), .ZN(new_n1230));
  NAND2_X1  g804(.A1(new_n1229), .A2(new_n1230), .ZN(G225));
endmodule


