//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  XNOR2_X1  g010(.A(G125), .B(G140), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n201));
  INV_X1    g015(.A(G953), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G237), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT69), .A2(G953), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n203), .A2(G214), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT69), .A2(G953), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT69), .A2(G953), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n211), .A2(G143), .A3(G214), .A4(new_n204), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT88), .A2(KEYINPUT18), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n208), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n206), .A2(new_n207), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n206), .A2(new_n207), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n200), .B(new_n215), .C1(new_n218), .C2(new_n214), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n208), .A2(new_n212), .A3(new_n213), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n213), .B1(new_n208), .B2(new_n212), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT17), .ZN(new_n223));
  OAI211_X1 g037(.A(KEYINPUT17), .B(G131), .C1(new_n216), .C2(new_n217), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT79), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT16), .ZN(new_n226));
  OR3_X1    g040(.A1(new_n193), .A2(KEYINPUT16), .A3(G140), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n193), .A2(KEYINPUT16), .A3(G140), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT79), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n198), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n225), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n229), .B1(new_n197), .B2(KEYINPUT16), .ZN(new_n233));
  OAI211_X1 g047(.A(G146), .B(new_n232), .C1(new_n233), .C2(new_n225), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n224), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n190), .B(new_n219), .C1(new_n223), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT91), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n218), .A2(new_n238), .A3(new_n220), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(new_n231), .A3(new_n234), .A4(new_n224), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n240), .A2(new_n241), .A3(new_n190), .A4(new_n219), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT19), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n192), .A2(new_n194), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT90), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT89), .B1(new_n197), .B2(new_n244), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT89), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n195), .A2(new_n248), .A3(KEYINPUT19), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n246), .A2(new_n198), .A3(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n251), .B(new_n234), .C1(new_n222), .C2(new_n221), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n190), .B1(new_n252), .B2(new_n219), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT92), .B1(new_n243), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n256));
  AOI211_X1 g070(.A(new_n256), .B(new_n253), .C1(new_n237), .C2(new_n242), .ZN(new_n257));
  NOR2_X1   g071(.A1(G475), .A2(G902), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n258), .B(KEYINPUT93), .Z(new_n259));
  NOR3_X1   g073(.A1(new_n255), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT20), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n187), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n243), .A2(new_n254), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n256), .ZN(new_n264));
  INV_X1    g078(.A(new_n259), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n243), .A2(KEYINPUT92), .A3(new_n254), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n259), .A2(KEYINPUT20), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n262), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G902), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n190), .B1(new_n240), .B2(new_n219), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(KEYINPUT95), .ZN(new_n274));
  INV_X1    g088(.A(new_n243), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G475), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(G210), .B1(G237), .B2(G902), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n279), .B(KEYINPUT86), .Z(new_n280));
  OAI21_X1  g094(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n282));
  INV_X1    g096(.A(G107), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(G104), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n189), .A2(G107), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n281), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G101), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT4), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n284), .A2(new_n285), .ZN(new_n291));
  INV_X1    g105(.A(G101), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n291), .A2(KEYINPUT82), .A3(new_n292), .A4(new_n281), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n281), .A2(new_n284), .A3(new_n292), .A4(new_n285), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT82), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n288), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n287), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n290), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G116), .ZN(new_n301));
  INV_X1    g115(.A(G116), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT2), .B(G113), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n306), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n283), .A2(G104), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n285), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n293), .A2(new_n296), .B1(G101), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n305), .A2(KEYINPUT5), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n301), .A2(KEYINPUT5), .ZN(new_n316));
  INV_X1    g130(.A(G113), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n315), .A2(new_n318), .B1(new_n305), .B2(new_n307), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n299), .A2(new_n311), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G122), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n314), .B(new_n319), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(KEYINPUT8), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(KEYINPUT0), .A2(G128), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n198), .A2(G143), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n207), .A2(KEYINPUT65), .A3(G146), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT65), .B1(new_n207), .B2(G146), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n327), .B(new_n328), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n207), .A2(G146), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  OR2_X1    g147(.A1(KEYINPUT0), .A2(G128), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n326), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n193), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n207), .A2(G146), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n339));
  OAI21_X1  g153(.A(G128), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n333), .ZN(new_n341));
  INV_X1    g155(.A(G128), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(KEYINPUT1), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n328), .B(new_n343), .C1(new_n329), .C2(new_n330), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n337), .B1(G125), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G224), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT7), .B1(new_n347), .B2(G953), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT84), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n348), .B1(new_n336), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n345), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n193), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(new_n349), .A3(new_n337), .A4(new_n348), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n325), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT85), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n322), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n323), .A2(new_n324), .B1(new_n351), .B2(new_n354), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(KEYINPUT85), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n272), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n314), .A2(new_n319), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n294), .A2(new_n295), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n294), .A2(new_n295), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT4), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n289), .B1(new_n365), .B2(new_n287), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n362), .B1(new_n366), .B2(new_n310), .ZN(new_n367));
  INV_X1    g181(.A(new_n321), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n322), .A3(KEYINPUT6), .ZN(new_n370));
  OR3_X1    g184(.A1(new_n320), .A2(KEYINPUT6), .A3(new_n321), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n347), .A2(G953), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n346), .B(new_n372), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n280), .B1(new_n361), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n359), .A2(KEYINPUT85), .B1(new_n321), .B2(new_n320), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n356), .A2(new_n357), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n280), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n375), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(KEYINPUT87), .B(new_n280), .C1(new_n361), .C2(new_n374), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G214), .B1(G237), .B2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT9), .B(G234), .ZN(new_n389));
  OAI21_X1  g203(.A(G221), .B1(new_n389), .B2(G902), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n390), .B(KEYINPUT81), .Z(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G469), .ZN(new_n393));
  INV_X1    g207(.A(G134), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G137), .ZN(new_n395));
  INV_X1    g209(.A(G137), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT66), .B1(new_n396), .B2(G134), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT11), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n395), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT66), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n394), .B2(G137), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(KEYINPUT11), .ZN(new_n402));
  OAI21_X1  g216(.A(G131), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT67), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n396), .A2(G134), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n401), .B2(KEYINPUT11), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n397), .A2(new_n398), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n213), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n403), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(KEYINPUT67), .B(G131), .C1(new_n399), .C2(new_n402), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n313), .A2(G101), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n363), .B2(new_n364), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n352), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n332), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n207), .A2(KEYINPUT65), .A3(G146), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n338), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n342), .B1(new_n328), .B2(KEYINPUT1), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n344), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n420), .B(new_n412), .C1(new_n363), .C2(new_n364), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n411), .B1(new_n414), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT12), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n331), .A2(new_n335), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT68), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT68), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n331), .A2(new_n335), .A3(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT10), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n352), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n299), .A2(new_n428), .B1(new_n314), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT83), .B1(new_n421), .B2(new_n429), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n421), .A2(KEYINPUT83), .A3(new_n429), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n431), .B(new_n411), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n211), .A2(G227), .ZN(new_n435));
  XOR2_X1   g249(.A(G110), .B(G140), .Z(new_n436));
  XNOR2_X1  g250(.A(new_n435), .B(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n423), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n411), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n433), .A2(new_n432), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n299), .A2(new_n428), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n430), .A2(new_n314), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n440), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n438), .B1(new_n445), .B2(new_n434), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n393), .B(new_n272), .C1(new_n439), .C2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n434), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT12), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n422), .B(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n437), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n445), .A2(new_n434), .A3(new_n438), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(G469), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n393), .A2(new_n272), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n392), .B1(new_n448), .B2(new_n457), .ZN(new_n458));
  XOR2_X1   g272(.A(KEYINPUT77), .B(G217), .Z(new_n459));
  INV_X1    g273(.A(G234), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n460), .B2(G902), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n211), .A2(G221), .A3(G234), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT22), .B(G137), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n462), .B(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n342), .A2(KEYINPUT23), .A3(G119), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n300), .A2(G128), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n300), .A2(G128), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(KEYINPUT23), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G110), .ZN(new_n470));
  INV_X1    g284(.A(G110), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT24), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT24), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G110), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(G119), .B(G128), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT78), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n475), .B2(new_n476), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n470), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n231), .B2(new_n234), .ZN(new_n481));
  OAI22_X1  g295(.A1(new_n469), .A2(G110), .B1(new_n476), .B2(new_n475), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n234), .A2(new_n482), .A3(new_n199), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n465), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n231), .A2(new_n234), .ZN(new_n485));
  INV_X1    g299(.A(new_n480), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n234), .A2(new_n482), .A3(new_n199), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n464), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT25), .ZN(new_n490));
  AOI21_X1  g304(.A(G902), .B1(new_n490), .B2(KEYINPUT80), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n484), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n490), .A2(KEYINPUT80), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n461), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n493), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n484), .A2(new_n489), .A3(new_n495), .A4(new_n491), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n484), .A2(new_n489), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n461), .A2(new_n272), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n458), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n342), .A2(G143), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n207), .A2(G128), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(new_n394), .ZN(new_n508));
  XNOR2_X1  g322(.A(G116), .B(G122), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n283), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n302), .A2(KEYINPUT14), .A3(G122), .ZN(new_n511));
  INV_X1    g325(.A(new_n509), .ZN(new_n512));
  OAI211_X1 g326(.A(G107), .B(new_n511), .C1(new_n512), .C2(KEYINPUT14), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n508), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n506), .B1(KEYINPUT13), .B2(new_n505), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT13), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n342), .B2(G143), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n394), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT96), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n507), .A2(new_n394), .ZN(new_n520));
  INV_X1    g334(.A(new_n510), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n509), .A2(new_n283), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n514), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n389), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(new_n459), .A3(new_n202), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n524), .B(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT97), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n272), .ZN(new_n529));
  INV_X1    g343(.A(G478), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(KEYINPUT15), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n529), .B(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n202), .A2(G952), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n460), .B2(new_n204), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  AOI211_X1 g349(.A(new_n272), .B(new_n211), .C1(G234), .C2(G237), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT98), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT21), .B(G898), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n532), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n278), .A2(new_n388), .A3(new_n504), .A4(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n409), .A2(new_n425), .A3(new_n410), .A4(new_n427), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n394), .A2(G137), .ZN(new_n543));
  OAI21_X1  g357(.A(G131), .B1(new_n543), .B2(new_n405), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n345), .A2(new_n408), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n310), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT28), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n542), .A2(new_n548), .A3(new_n310), .A4(new_n545), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n542), .A2(new_n545), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n547), .A2(new_n549), .B1(new_n550), .B2(new_n311), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT75), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n211), .A2(G210), .A3(new_n204), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT27), .ZN(new_n554));
  XOR2_X1   g368(.A(KEYINPUT26), .B(G101), .Z(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT29), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n551), .A2(new_n552), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n272), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n552), .B1(new_n551), .B2(new_n558), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT76), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n424), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n409), .A2(new_n410), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n545), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n547), .A2(new_n549), .B1(new_n311), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(new_n556), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n556), .A2(new_n546), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n542), .A2(KEYINPUT30), .A3(new_n545), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n311), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n557), .B1(new_n567), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n551), .A2(new_n558), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT75), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT76), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n272), .A4(new_n559), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n562), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G472), .ZN(new_n581));
  INV_X1    g395(.A(new_n556), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT71), .B1(new_n566), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n547), .A2(new_n549), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n565), .A2(new_n311), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT71), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n556), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT70), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n556), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n573), .A2(new_n546), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT31), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n573), .A2(KEYINPUT31), .A3(new_n546), .A4(new_n590), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n583), .A2(new_n588), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(G472), .A2(G902), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT72), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT32), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n581), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT73), .B1(new_n595), .B2(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n588), .A2(new_n583), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n593), .A2(new_n594), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT73), .ZN(new_n605));
  INV_X1    g419(.A(new_n597), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT32), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n601), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT74), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n601), .A2(new_n607), .A3(KEYINPUT74), .A4(new_n608), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n600), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n541), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT99), .B(G101), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G3));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n524), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n526), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n524), .A2(new_n617), .A3(new_n526), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(KEYINPUT33), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT101), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n620), .A2(new_n624), .A3(KEYINPUT33), .A4(new_n621), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n527), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n530), .A2(G902), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n623), .A2(new_n625), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n527), .A2(new_n272), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n530), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n271), .B2(new_n277), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n380), .B1(new_n379), .B2(new_n381), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n386), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n539), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(G472), .B1(new_n595), .B2(G902), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n601), .A2(new_n640), .A3(new_n607), .ZN(new_n641));
  INV_X1    g455(.A(new_n504), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT34), .B(G104), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  NAND3_X1  g459(.A1(new_n264), .A2(new_n266), .A3(new_n269), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT102), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n255), .A2(new_n257), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n649), .A3(new_n269), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n262), .A2(new_n268), .A3(new_n647), .A4(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n638), .A2(new_n277), .A3(new_n532), .A4(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n652), .A2(new_n642), .A3(new_n641), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NAND3_X1  g469(.A1(new_n278), .A2(new_n388), .A3(new_n540), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT103), .B1(new_n481), .B2(new_n483), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n487), .A2(new_n659), .A3(new_n488), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n465), .A2(KEYINPUT36), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n661), .B1(new_n658), .B2(new_n660), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n501), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n497), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT104), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n497), .A2(new_n667), .A3(new_n664), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n669), .B(new_n392), .C1(new_n448), .C2(new_n457), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n641), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n657), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT105), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT37), .B(G110), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NAND2_X1  g489(.A1(new_n611), .A2(new_n612), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n580), .A2(G472), .B1(new_n598), .B2(KEYINPUT32), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n535), .B1(new_n537), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n651), .A2(new_n277), .A3(new_n532), .A4(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n457), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n391), .B1(new_n683), .B2(new_n447), .ZN(new_n684));
  INV_X1    g498(.A(new_n637), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n669), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n678), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  INV_X1    g503(.A(G472), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n573), .A2(new_n546), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n582), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n550), .A2(new_n311), .ZN(new_n693));
  AOI21_X1  g507(.A(G902), .B1(new_n569), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n690), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n598), .B2(KEYINPUT32), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n676), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n680), .B(KEYINPUT39), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n684), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT40), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n385), .B(KEYINPUT38), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n271), .A2(new_n277), .ZN(new_n702));
  INV_X1    g516(.A(new_n669), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n702), .A2(new_n386), .A3(new_n532), .A4(new_n703), .ZN(new_n704));
  OR4_X1    g518(.A1(new_n697), .A2(new_n700), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  NAND3_X1  g520(.A1(new_n702), .A2(new_n632), .A3(new_n681), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n686), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n678), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  OAI21_X1  g524(.A(new_n272), .B1(new_n439), .B2(new_n446), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n392), .A3(new_n447), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n503), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n634), .A2(new_n638), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n613), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT41), .B(G113), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  INV_X1    g532(.A(new_n714), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n652), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n678), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NOR2_X1   g536(.A1(new_n713), .A2(new_n637), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n278), .A2(new_n540), .A3(new_n669), .A4(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n613), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n300), .ZN(G21));
  OAI211_X1 g540(.A(new_n386), .B(new_n532), .C1(new_n635), .C2(new_n636), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n713), .A2(new_n539), .ZN(new_n729));
  INV_X1    g543(.A(new_n503), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n551), .A2(new_n582), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n603), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n606), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n640), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n702), .A2(new_n728), .A3(new_n729), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n737));
  AOI21_X1  g551(.A(G902), .B1(new_n602), .B2(new_n603), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n669), .B(new_n733), .C1(new_n738), .C2(new_n690), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n723), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n737), .B1(new_n707), .B2(new_n741), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n739), .A2(new_n713), .A3(new_n637), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n634), .A3(KEYINPUT106), .A4(new_n681), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  AOI21_X1  g560(.A(new_n387), .B1(new_n383), .B2(new_n384), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n684), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n613), .A2(new_n503), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n707), .A2(KEYINPUT42), .ZN(new_n750));
  AOI211_X1 g564(.A(new_n680), .B(new_n633), .C1(new_n271), .C2(new_n277), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n747), .A2(new_n684), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n608), .B1(new_n595), .B2(new_n597), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n503), .B1(new_n677), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n749), .A2(new_n750), .B1(KEYINPUT42), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  NOR4_X1   g571(.A1(new_n613), .A2(new_n503), .A3(new_n682), .A4(new_n748), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n394), .ZN(G36));
  XNOR2_X1  g573(.A(new_n702), .B(KEYINPUT108), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(KEYINPUT43), .A3(new_n632), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n702), .B2(new_n633), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n641), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n703), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT44), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n452), .A2(new_n453), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n393), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n769), .B2(new_n768), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n455), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n447), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n392), .ZN(new_n778));
  INV_X1    g592(.A(new_n698), .ZN(new_n779));
  INV_X1    g593(.A(new_n747), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n767), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n764), .A2(KEYINPUT44), .A3(new_n766), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT109), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G137), .ZN(G39));
  NAND4_X1  g599(.A1(new_n613), .A2(new_n751), .A3(new_n503), .A4(new_n747), .ZN(new_n786));
  INV_X1    g600(.A(new_n778), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT47), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n778), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n786), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n191), .ZN(G42));
  NAND2_X1  g606(.A1(new_n712), .A2(new_n447), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(KEYINPUT49), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(KEYINPUT49), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n632), .A2(new_n392), .A3(new_n730), .A4(new_n386), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n697), .A2(new_n760), .A3(new_n701), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n713), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n701), .A2(new_n387), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT114), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(KEYINPUT115), .B2(KEYINPUT50), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n534), .B1(new_n761), .B2(new_n763), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n734), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n805), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n764), .A2(new_n535), .A3(new_n799), .A4(new_n747), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT116), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT116), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n739), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n503), .A2(new_n534), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n697), .A2(new_n799), .A3(new_n747), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT117), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n278), .A3(new_n633), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n809), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n809), .A2(new_n814), .A3(KEYINPUT118), .A4(new_n818), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n788), .B(new_n790), .C1(new_n392), .C2(new_n793), .ZN(new_n823));
  INV_X1    g637(.A(new_n804), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n747), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n821), .A2(new_n822), .A3(KEYINPUT51), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n723), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n533), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n634), .B2(new_n817), .ZN(new_n829));
  INV_X1    g643(.A(new_n754), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n811), .B2(new_n812), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT48), .ZN(new_n833));
  XOR2_X1   g647(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n834));
  OAI211_X1 g648(.A(new_n829), .B(new_n833), .C1(new_n831), .C2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n825), .A2(new_n814), .A3(new_n809), .A4(new_n818), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n826), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n751), .A2(new_n640), .A3(new_n733), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n532), .A2(new_n680), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n651), .A2(new_n277), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT110), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT110), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n651), .A2(new_n844), .A3(new_n277), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n840), .B1(new_n846), .B2(new_n613), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n748), .A2(new_n703), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n758), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n634), .B1(new_n278), .B2(new_n532), .ZN(new_n850));
  INV_X1    g664(.A(new_n539), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n388), .A2(new_n504), .A3(new_n851), .A4(new_n765), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n671), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n735), .B1(new_n656), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n651), .A2(new_n277), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n532), .A3(new_n638), .A4(new_n714), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n613), .B1(new_n858), .B2(new_n724), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n613), .B1(new_n541), .B2(new_n715), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n849), .A2(new_n756), .A3(new_n856), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT106), .B1(new_n751), .B2(new_n743), .ZN(new_n865));
  AND4_X1   g679(.A1(KEYINPUT106), .A2(new_n743), .A3(new_n634), .A4(new_n681), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n688), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n665), .A2(new_n680), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n702), .A2(new_n684), .A3(new_n728), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n670), .A2(new_n637), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n751), .A2(new_n870), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n697), .A2(new_n869), .B1(new_n871), .B2(new_n613), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n864), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n742), .A2(new_n744), .B1(new_n678), .B2(new_n687), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n676), .A2(new_n696), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n392), .B(new_n868), .C1(new_n448), .C2(new_n457), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n727), .B(new_n876), .C1(new_n277), .C2(new_n271), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n708), .A2(new_n678), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n874), .A2(KEYINPUT111), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n862), .B1(new_n863), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n873), .A2(new_n879), .A3(KEYINPUT52), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(KEYINPUT53), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT52), .B1(new_n867), .B2(new_n872), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n885), .B2(KEYINPUT53), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n874), .A2(KEYINPUT111), .A3(new_n878), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT111), .B1(new_n874), .B2(new_n878), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n863), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n847), .A2(new_n848), .ZN(new_n891));
  INV_X1    g705(.A(new_n758), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n756), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n861), .A2(new_n856), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n890), .A2(new_n895), .A3(new_n882), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT112), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n881), .A2(KEYINPUT53), .A3(new_n884), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n896), .A2(KEYINPUT112), .A3(new_n897), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n899), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n887), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n904), .A2(KEYINPUT113), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(KEYINPUT113), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n839), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(G952), .A2(G953), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n798), .B1(new_n907), .B2(new_n908), .ZN(G75));
  NAND2_X1  g723(.A1(new_n370), .A2(new_n371), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(new_n373), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT55), .Z(new_n912));
  NAND2_X1  g726(.A1(new_n902), .A2(new_n901), .ZN(new_n913));
  OAI211_X1 g727(.A(G902), .B(new_n280), .C1(new_n913), .C2(new_n898), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n915), .B2(KEYINPUT56), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  INV_X1    g731(.A(new_n912), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n211), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n916), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n916), .A2(KEYINPUT120), .A3(new_n919), .A4(new_n921), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(G51));
  OAI21_X1  g740(.A(KEYINPUT54), .B1(new_n913), .B2(new_n898), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n903), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(KEYINPUT121), .B(KEYINPUT54), .C1(new_n913), .C2(new_n898), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n455), .B(KEYINPUT57), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n446), .B2(new_n439), .ZN(new_n933));
  AND4_X1   g747(.A1(KEYINPUT53), .A2(new_n890), .A3(new_n895), .A4(new_n884), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT53), .B1(new_n881), .B2(new_n882), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(KEYINPUT112), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n272), .B1(new_n936), .B2(new_n899), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n773), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n920), .B1(new_n933), .B2(new_n938), .ZN(G54));
  NAND3_X1  g753(.A1(new_n937), .A2(KEYINPUT58), .A3(G475), .ZN(new_n940));
  INV_X1    g754(.A(new_n648), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n920), .ZN(G60));
  NAND3_X1  g758(.A1(new_n623), .A2(new_n625), .A3(new_n627), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT59), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n929), .A2(new_n930), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n921), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n905), .A2(new_n906), .A3(new_n948), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n950), .B1(new_n951), .B2(new_n945), .ZN(G63));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT60), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n936), .B2(new_n899), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n499), .ZN(new_n957));
  INV_X1    g771(.A(new_n955), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n662), .A2(new_n663), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT122), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n958), .B(new_n960), .C1(new_n913), .C2(new_n898), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n921), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n953), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n958), .B1(new_n913), .B2(new_n898), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n965), .A2(new_n966), .A3(new_n498), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n965), .B2(new_n498), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n961), .A2(KEYINPUT61), .A3(new_n921), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT123), .B1(new_n956), .B2(new_n499), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n965), .A2(new_n966), .A3(new_n498), .ZN(new_n973));
  AND4_X1   g787(.A1(new_n964), .A2(new_n970), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n963), .B1(new_n971), .B2(new_n974), .ZN(G66));
  OAI21_X1  g789(.A(G953), .B1(new_n538), .B2(new_n347), .ZN(new_n976));
  INV_X1    g790(.A(new_n894), .ZN(new_n977));
  INV_X1    g791(.A(new_n211), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n910), .B1(G898), .B2(new_n211), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G69));
  NAND2_X1  g795(.A1(new_n571), .A2(new_n572), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n246), .A2(new_n250), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n978), .A2(G900), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n278), .A2(new_n727), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n787), .A2(new_n698), .A3(new_n986), .A4(new_n754), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n987), .A2(new_n756), .A3(new_n892), .ZN(new_n988));
  INV_X1    g802(.A(new_n791), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n874), .A2(new_n709), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n988), .A2(new_n989), .A3(new_n784), .A4(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n984), .B(new_n985), .C1(new_n991), .C2(new_n978), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n705), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT125), .Z(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n850), .A2(new_n699), .A3(new_n780), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(new_n678), .A3(new_n730), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT126), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n791), .A2(new_n999), .ZN(new_n1000));
  AND4_X1   g814(.A1(new_n784), .A2(new_n995), .A3(new_n996), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1001), .A2(new_n978), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n992), .B1(new_n1002), .B2(new_n984), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n211), .B1(G227), .B2(G900), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1004), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n992), .B(new_n1006), .C1(new_n1002), .C2(new_n984), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(G72));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  OAI21_X1  g824(.A(new_n1010), .B1(new_n991), .B2(new_n894), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n920), .B1(new_n1011), .B2(new_n574), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1010), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(new_n1001), .B2(new_n977), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1012), .B1(new_n1014), .B2(new_n692), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n574), .A2(new_n1013), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n886), .A2(new_n692), .A3(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT127), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1015), .A2(new_n1018), .ZN(G57));
endmodule


