//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT66), .B(KEYINPUT0), .Z(new_n217));
  XNOR2_X1  g0017(.A(new_n216), .B(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n203), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n214), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n212), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n206), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n218), .B(new_n230), .C1(new_n232), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n225), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n231), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n212), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n256), .A2(new_n258), .B1(G150), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n253), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n252), .ZN(new_n264));
  INV_X1    g0064(.A(G50), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(new_n211), .B2(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G50), .B2(new_n262), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G222), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  OAI221_X1 g0075(.A(new_n272), .B1(new_n273), .B2(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  INV_X1    g0081(.A(new_n231), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(new_n277), .ZN(new_n283));
  XOR2_X1   g0083(.A(KEYINPUT68), .B(G45), .Z(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G41), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n283), .B(new_n211), .C1(new_n284), .C2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n278), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G226), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n280), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G179), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI211_X1 g0096(.A(new_n269), .B(new_n295), .C1(new_n296), .C2(new_n294), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(G200), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n294), .A2(new_n301), .B1(new_n269), .B2(KEYINPUT9), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n297), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n256), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n221), .A2(KEYINPUT15), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT15), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G87), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT69), .B1(new_n312), .B2(new_n257), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n312), .A2(KEYINPUT69), .A3(new_n257), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n252), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n273), .B1(new_n211), .B2(G20), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n264), .A2(new_n317), .B1(new_n273), .B2(new_n263), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G107), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n274), .A2(new_n220), .B1(new_n320), .B2(new_n270), .ZN(new_n321));
  INV_X1    g0121(.A(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n326), .A2(new_n225), .A3(G1698), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n279), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT67), .B(G41), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT68), .B(G45), .ZN(new_n330));
  AOI21_X1  g0130(.A(G1), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(new_n283), .B1(new_n292), .B2(G244), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n319), .B1(new_n333), .B2(G200), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n328), .A2(G190), .A3(new_n332), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n328), .A2(new_n336), .A3(new_n332), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n333), .A2(new_n296), .B1(new_n316), .B2(new_n318), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n334), .A2(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n306), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT7), .B1(new_n326), .B2(new_n212), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  AOI211_X1 g0142(.A(new_n342), .B(G20), .C1(new_n323), .C2(new_n325), .ZN(new_n343));
  OAI21_X1  g0143(.A(G68), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G58), .A2(G68), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n204), .A2(new_n205), .A3(new_n345), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(KEYINPUT16), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n342), .B1(new_n270), .B2(G20), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n326), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n203), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n346), .A2(G20), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n259), .A2(G159), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n349), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n348), .A2(new_n356), .A3(new_n252), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT73), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n348), .A2(new_n356), .A3(KEYINPUT73), .A4(new_n252), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n264), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n211), .A2(G20), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n256), .A2(new_n363), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n362), .A2(new_n364), .B1(new_n262), .B2(new_n256), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n323), .A2(new_n325), .A3(G226), .A4(G1698), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n323), .A2(new_n325), .A3(G223), .A4(new_n271), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G87), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n279), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT74), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n292), .A2(G232), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n290), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT74), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n370), .A2(new_n375), .A3(new_n279), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n372), .A2(new_n374), .A3(new_n301), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  INV_X1    g0178(.A(new_n371), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n290), .A2(new_n373), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n361), .A2(new_n366), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT17), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n344), .A2(new_n347), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n253), .B1(new_n386), .B2(new_n349), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT73), .B1(new_n387), .B2(new_n348), .ZN(new_n388));
  INV_X1    g0188(.A(new_n360), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n366), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n376), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n290), .A2(new_n373), .A3(new_n336), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n375), .B1(new_n370), .B2(new_n279), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(G169), .B1(new_n374), .B2(new_n371), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT75), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT75), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n372), .A2(new_n374), .A3(new_n336), .A4(new_n376), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n296), .B1(new_n379), .B2(new_n380), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT18), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n390), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n365), .B1(new_n359), .B2(new_n360), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT75), .B1(new_n394), .B2(new_n395), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n398), .A2(new_n399), .A3(new_n397), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT18), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(KEYINPUT17), .A3(new_n382), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n385), .A2(new_n403), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n331), .A2(new_n283), .B1(new_n292), .B2(G238), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT13), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n323), .A2(new_n325), .A3(G232), .A4(G1698), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n323), .A2(new_n325), .A3(G226), .A4(new_n271), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G97), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n279), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n411), .A2(new_n412), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n412), .B1(new_n411), .B2(new_n417), .ZN(new_n420));
  OAI21_X1  g0220(.A(G200), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n420), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(G190), .A3(new_n418), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n264), .A2(G68), .A3(new_n363), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n273), .B2(new_n257), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT11), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n426), .A2(new_n427), .A3(new_n252), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n426), .B2(new_n252), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n263), .A2(new_n203), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT71), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n432), .B1(new_n431), .B2(new_n433), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n431), .A2(KEYINPUT12), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n421), .A2(new_n423), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT72), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT72), .A4(new_n438), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n438), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT14), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n445), .B(G169), .C1(new_n419), .C2(new_n420), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n422), .A2(new_n418), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n336), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n445), .B1(new_n447), .B2(G169), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n340), .A2(new_n410), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n320), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT25), .B1(new_n263), .B2(new_n320), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n211), .A2(G33), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n262), .A2(new_n456), .A3(new_n231), .A4(new_n251), .ZN(new_n457));
  OAI22_X1  g0257(.A1(new_n454), .A2(new_n455), .B1(new_n320), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT83), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n323), .A2(new_n325), .A3(new_n212), .A4(G87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT22), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT22), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n270), .A2(new_n463), .A3(new_n212), .A4(G87), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n212), .A2(G33), .A3(G116), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(new_n320), .A3(G20), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT23), .B1(new_n212), .B2(G107), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT82), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n466), .B(new_n468), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n320), .A2(G20), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT82), .B1(new_n472), .B2(KEYINPUT23), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT24), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n465), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n460), .B1(new_n479), .B2(new_n252), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n465), .A2(new_n477), .A3(new_n474), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n477), .B1(new_n465), .B2(new_n474), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n460), .B(new_n252), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n459), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT5), .B1(new_n286), .B2(new_n288), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT5), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n211), .B(G45), .C1(new_n487), .C2(G41), .ZN(new_n488));
  OAI211_X1 g0288(.A(G264), .B(new_n278), .C1(new_n486), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n488), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n283), .B(new_n490), .C1(KEYINPUT5), .C2(new_n329), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G250), .A2(G1698), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n227), .B2(G1698), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n493), .A2(new_n270), .B1(G33), .B2(G294), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n489), .B(new_n491), .C1(new_n494), .C2(new_n278), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT84), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n227), .A2(G1698), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(G250), .B2(G1698), .ZN(new_n498));
  INV_X1    g0298(.A(G294), .ZN(new_n499));
  OAI22_X1  g0299(.A1(new_n498), .A2(new_n326), .B1(new_n322), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n279), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT84), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(new_n491), .A4(new_n489), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n496), .A2(G169), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n495), .A2(new_n336), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT85), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n496), .A2(new_n507), .A3(G169), .A4(new_n503), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n485), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT86), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n252), .B1(new_n481), .B2(new_n482), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT83), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n458), .B1(new_n513), .B2(new_n483), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n495), .A2(new_n378), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n496), .A2(new_n503), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(G190), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n510), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n511), .B1(new_n510), .B2(new_n518), .ZN(new_n520));
  OR2_X1    g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n522), .B(new_n212), .C1(G33), .C2(new_n226), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G20), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n252), .A3(new_n525), .ZN(new_n526));
  OR2_X1    g0326(.A1(KEYINPUT80), .A2(KEYINPUT20), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g0328(.A(KEYINPUT80), .B(KEYINPUT20), .Z(new_n529));
  AOI22_X1  g0329(.A1(new_n526), .A2(new_n529), .B1(new_n524), .B2(new_n263), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT79), .ZN(new_n531));
  INV_X1    g0331(.A(new_n457), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n532), .B2(G116), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n457), .A2(KEYINPUT79), .A3(new_n524), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n528), .B(new_n530), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G303), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n278), .B1(new_n326), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(G257), .A2(G1698), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n271), .A2(G264), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n270), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G270), .B(new_n278), .C1(new_n486), .C2(new_n488), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(new_n491), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n535), .A2(KEYINPUT21), .A3(G169), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT81), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n543), .A2(G169), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT81), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT21), .A4(new_n535), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n535), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT21), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n541), .A2(new_n542), .A3(new_n491), .A4(G179), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n550), .A2(new_n551), .B1(new_n535), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT6), .ZN(new_n556));
  AND2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G97), .A2(G107), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n320), .A2(KEYINPUT6), .A3(G97), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G20), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n259), .A2(G77), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n320), .B1(new_n350), .B2(new_n351), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n252), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n532), .A2(G97), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n262), .A2(G97), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n566), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n323), .A2(new_n325), .A3(G244), .A4(new_n271), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT4), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n323), .A2(new_n325), .A3(G250), .A4(G1698), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .A4(new_n522), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n279), .ZN(new_n579));
  OAI211_X1 g0379(.A(G257), .B(new_n278), .C1(new_n486), .C2(new_n488), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n580), .A2(new_n491), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n296), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(new_n491), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n279), .B2(new_n578), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n336), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n572), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n588));
  OAI21_X1  g0388(.A(G107), .B1(new_n341), .B2(new_n343), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n561), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n588), .B1(new_n591), .B2(new_n252), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n579), .A2(new_n581), .A3(G190), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n592), .B(new_n593), .C1(new_n378), .C2(new_n585), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n323), .A2(new_n325), .A3(G244), .A4(G1698), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n323), .A2(new_n325), .A3(G238), .A4(new_n271), .ZN(new_n596));
  NAND2_X1  g0396(.A1(G33), .A2(G116), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n279), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n211), .A2(G45), .ZN(new_n600));
  NAND2_X1  g0400(.A1(KEYINPUT77), .A2(G250), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n282), .A2(new_n277), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(G45), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(G1), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n604), .B(new_n281), .C1(KEYINPUT77), .C2(new_n222), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n599), .A2(new_n301), .A3(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n598), .A2(new_n279), .B1(new_n605), .B2(new_n602), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n607), .B1(G200), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n457), .A2(new_n221), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n311), .A2(new_n262), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT19), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n212), .B1(new_n415), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n558), .A2(new_n221), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n323), .A2(new_n325), .A3(new_n212), .A4(G68), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n613), .B1(new_n257), .B2(new_n226), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI211_X1 g0419(.A(KEYINPUT78), .B(new_n612), .C1(new_n619), .C2(new_n252), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT78), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n252), .ZN(new_n622));
  INV_X1    g0422(.A(new_n612), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n609), .B(new_n611), .C1(new_n620), .C2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n312), .A2(new_n457), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n624), .B2(new_n620), .ZN(new_n628));
  AOI221_X4 g0428(.A(G179), .B1(new_n605), .B2(new_n602), .C1(new_n598), .C2(new_n279), .ZN(new_n629));
  AOI21_X1  g0429(.A(G169), .B1(new_n599), .B2(new_n606), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n587), .A2(new_n594), .A3(new_n625), .A4(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n543), .A2(new_n301), .ZN(new_n634));
  AOI211_X1 g0434(.A(new_n535), .B(new_n634), .C1(G200), .C2(new_n543), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n555), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n452), .A2(new_n521), .A3(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n632), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n622), .A2(new_n623), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT78), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n622), .A2(new_n621), .A3(new_n623), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n626), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n608), .A2(new_n336), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(G169), .B2(new_n608), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n611), .B1(new_n624), .B2(new_n620), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n599), .A2(new_n301), .A3(new_n606), .ZN(new_n647));
  AOI21_X1  g0447(.A(G200), .B1(new_n599), .B2(new_n606), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n643), .A2(new_n645), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n639), .B1(new_n650), .B2(new_n587), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n610), .B1(new_n641), .B2(new_n642), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n652), .A2(new_n609), .B1(new_n628), .B2(new_n631), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n579), .A2(new_n581), .A3(new_n336), .ZN(new_n654));
  AOI21_X1  g0454(.A(G169), .B1(new_n579), .B2(new_n581), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n654), .A2(new_n592), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n653), .A2(KEYINPUT26), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n638), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n555), .B1(new_n485), .B2(new_n509), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n587), .A2(new_n594), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n518), .A2(new_n653), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n658), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n452), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n403), .A2(new_n408), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n385), .A2(new_n409), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n450), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n338), .A2(new_n337), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n443), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n664), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n304), .A2(new_n305), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n297), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n663), .A2(new_n673), .ZN(G369));
  INV_X1    g0474(.A(G330), .ZN(new_n675));
  OR3_X1    g0475(.A1(new_n555), .A2(KEYINPUT88), .A3(new_n635), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT88), .B1(new_n555), .B2(new_n635), .ZN(new_n677));
  INV_X1    g0477(.A(new_n535), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(G213), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n676), .B(new_n677), .C1(new_n678), .C2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n555), .A2(new_n535), .A3(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT87), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT89), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n686), .A2(new_n688), .A3(KEYINPUT89), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n675), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n521), .B1(new_n514), .B2(new_n685), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n485), .A2(new_n509), .A3(new_n684), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n510), .A2(new_n684), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n549), .A2(new_n554), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n684), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n698), .B1(new_n521), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(G399));
  NAND2_X1  g0502(.A1(new_n215), .A2(new_n329), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n615), .A2(G116), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n233), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n662), .A2(new_n685), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT92), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT92), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n662), .A2(new_n711), .A3(new_n685), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT93), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n653), .A2(KEYINPUT95), .A3(KEYINPUT26), .A4(new_n656), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n632), .A2(KEYINPUT94), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT94), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n628), .A2(new_n631), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n633), .B1(new_n514), .B2(new_n517), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n699), .A2(new_n510), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT95), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n651), .A2(new_n725), .A3(new_n657), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n684), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT29), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n709), .A2(KEYINPUT93), .A3(new_n710), .A4(new_n712), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n715), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n636), .B(new_n685), .C1(new_n519), .C2(new_n520), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n684), .A2(KEYINPUT31), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n608), .A2(new_n489), .A3(new_n501), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n582), .A2(new_n733), .A3(new_n552), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(KEYINPUT30), .ZN(new_n735));
  INV_X1    g0535(.A(new_n733), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(KEYINPUT30), .A3(new_n585), .A4(new_n553), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n543), .A2(new_n336), .ZN(new_n738));
  INV_X1    g0538(.A(new_n608), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n738), .A2(new_n582), .A3(new_n495), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n732), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT90), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(KEYINPUT90), .B(new_n732), .C1(new_n735), .C2(new_n741), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT91), .B1(new_n734), .B2(KEYINPUT30), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n736), .A2(new_n585), .A3(new_n553), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT91), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n747), .A2(new_n751), .A3(new_n737), .A4(new_n740), .ZN(new_n752));
  AOI21_X1  g0552(.A(KEYINPUT31), .B1(new_n752), .B2(new_n684), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n746), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n731), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n730), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n707), .B1(new_n758), .B2(G1), .ZN(G364));
  AND2_X1   g0559(.A1(new_n212), .A2(G13), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n211), .B1(new_n760), .B2(G45), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n703), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n215), .A2(new_n270), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n764), .A2(new_n209), .B1(G116), .B2(new_n215), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n215), .A2(new_n326), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT96), .Z(new_n767));
  AOI22_X1  g0567(.A1(new_n249), .A2(G45), .B1(new_n234), .B2(new_n330), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n231), .B1(G20), .B2(new_n296), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT97), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n763), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n301), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n336), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n270), .B1(new_n780), .B2(new_n226), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n212), .A2(new_n336), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n301), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n265), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n212), .A2(G179), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G190), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G159), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n781), .B(new_n786), .C1(KEYINPUT32), .C2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT98), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n782), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n212), .A2(new_n336), .A3(KEYINPUT98), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n777), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n788), .B1(new_n794), .B2(new_n795), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G58), .A2(new_n797), .B1(new_n799), .B2(G77), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n787), .A2(new_n301), .A3(G200), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G107), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n783), .A2(G190), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n805), .A2(new_n203), .B1(new_n791), .B2(KEYINPUT32), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n221), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n792), .A2(new_n800), .A3(new_n803), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n270), .B1(new_n790), .B2(G329), .ZN(new_n811));
  INV_X1    g0611(.A(G326), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n785), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n797), .B2(G322), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n799), .A2(G311), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n780), .A2(new_n499), .B1(new_n807), .B2(new_n536), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT33), .B(G317), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n816), .B1(new_n804), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n802), .A2(G283), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n814), .A2(new_n815), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n810), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n776), .B1(new_n821), .B2(new_n773), .ZN(new_n822));
  INV_X1    g0622(.A(new_n772), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n689), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n693), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n762), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n691), .A2(new_n675), .A3(new_n692), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT100), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  INV_X1    g0630(.A(KEYINPUT104), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n669), .A2(new_n831), .A3(new_n684), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT104), .B1(new_n668), .B2(new_n685), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n319), .A2(new_n684), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n832), .A2(new_n833), .B1(new_n339), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n709), .A2(new_n712), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n832), .A2(new_n833), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n339), .A2(new_n834), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n662), .A2(new_n685), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n763), .B1(new_n841), .B2(new_n756), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n756), .B2(new_n841), .ZN(new_n843));
  INV_X1    g0643(.A(new_n773), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n771), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n763), .B1(G77), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n802), .A2(G68), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n270), .B1(new_n789), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n807), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(G50), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n847), .B(new_n851), .C1(new_n202), .C2(new_n780), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT103), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G137), .A2(new_n784), .B1(new_n804), .B2(G150), .ZN(new_n854));
  INV_X1    g0654(.A(G143), .ZN(new_n855));
  INV_X1    g0655(.A(G159), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n854), .B1(new_n855), .B2(new_n796), .C1(new_n856), .C2(new_n798), .ZN(new_n857));
  XNOR2_X1  g0657(.A(KEYINPUT102), .B(KEYINPUT34), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n857), .B(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(G311), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n326), .B1(new_n789), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G97), .B2(new_n779), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n862), .B1(new_n524), .B2(new_n798), .C1(new_n499), .C2(new_n796), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n802), .A2(G87), .ZN(new_n864));
  XNOR2_X1  g0664(.A(KEYINPUT101), .B(G283), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n804), .A2(new_n866), .B1(new_n850), .B2(G107), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n864), .B(new_n867), .C1(new_n536), .C2(new_n785), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n853), .A2(new_n859), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n846), .B1(new_n869), .B2(new_n773), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n839), .B2(new_n771), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n843), .A2(new_n871), .ZN(G384));
  OR2_X1    g0672(.A1(new_n561), .A2(KEYINPUT35), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n561), .A2(KEYINPUT35), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n873), .A2(G116), .A3(new_n232), .A4(new_n874), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT36), .Z(new_n876));
  NAND3_X1  g0676(.A1(new_n234), .A2(G77), .A3(new_n345), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n265), .A2(G68), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n211), .B(G13), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n356), .A2(new_n252), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n881), .A2(KEYINPUT105), .ZN(new_n882));
  INV_X1    g0682(.A(new_n348), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n881), .B2(KEYINPUT105), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n365), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n383), .B1(new_n407), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n682), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n390), .A2(new_n401), .ZN(new_n889));
  INV_X1    g0689(.A(new_n682), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n390), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g0691(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n892));
  NAND4_X1  g0692(.A1(new_n889), .A2(new_n891), .A3(new_n383), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n410), .A2(new_n887), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n668), .A2(new_n684), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n840), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n444), .A2(new_n684), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n443), .A2(new_n450), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n443), .B2(new_n450), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n899), .A2(new_n908), .B1(new_n664), .B2(new_n890), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n897), .A2(new_n898), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n404), .A2(new_n407), .ZN(new_n913));
  AOI221_X4 g0713(.A(new_n365), .B1(new_n381), .B2(new_n377), .C1(new_n359), .C2(new_n360), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n892), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n915), .A2(KEYINPUT107), .A3(new_n916), .A4(new_n891), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n889), .A2(new_n891), .A3(new_n383), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT107), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n404), .B2(new_n682), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n916), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n891), .B1(new_n665), .B2(new_n664), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n912), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT39), .B1(new_n925), .B2(new_n896), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n911), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n667), .A2(new_n685), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n909), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n715), .A2(new_n452), .A3(new_n728), .A4(new_n729), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n673), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n930), .B(new_n932), .Z(new_n933));
  AND3_X1   g0733(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(new_n753), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n731), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n452), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT108), .Z(new_n938));
  OAI21_X1  g0738(.A(new_n839), .B1(new_n904), .B2(new_n905), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n731), .B2(new_n935), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n940), .B(new_n941), .C1(new_n897), .C2(new_n898), .ZN(new_n942));
  INV_X1    g0742(.A(new_n905), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n443), .A2(new_n450), .A3(new_n903), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n835), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n936), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n896), .B2(new_n925), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n942), .B1(new_n947), .B2(new_n941), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n675), .B1(new_n938), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n938), .B2(new_n948), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n933), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n211), .B2(new_n760), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n933), .A2(new_n950), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n880), .B1(new_n952), .B2(new_n953), .ZN(G367));
  XNOR2_X1  g0754(.A(new_n761), .B(KEYINPUT112), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT111), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n521), .A2(new_n700), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n957), .A2(KEYINPUT110), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n696), .B2(new_n700), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n957), .A2(KEYINPUT110), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n693), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n825), .A2(new_n959), .A3(new_n960), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n758), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT45), .ZN(new_n965));
  INV_X1    g0765(.A(new_n701), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n660), .B1(new_n592), .B2(new_n685), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n656), .A2(new_n684), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n965), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n701), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n966), .A2(KEYINPUT44), .A3(new_n970), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT44), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n701), .B2(new_n969), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n697), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n973), .A2(new_n697), .A3(new_n977), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n956), .B1(new_n964), .B2(new_n982), .ZN(new_n983));
  AND4_X1   g0783(.A1(new_n756), .A2(new_n962), .A3(new_n730), .A4(new_n963), .ZN(new_n984));
  INV_X1    g0784(.A(new_n981), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n697), .B1(new_n973), .B2(new_n977), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n987), .A3(KEYINPUT111), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n757), .B1(new_n983), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n703), .B(KEYINPUT41), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n955), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n646), .A2(new_n684), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT109), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n650), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n638), .B2(new_n993), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT43), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n521), .A2(new_n700), .A3(new_n969), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT42), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n587), .B1(new_n967), .B2(new_n510), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n998), .A2(KEYINPUT42), .B1(new_n685), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n997), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n995), .A2(new_n996), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n697), .A2(new_n970), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n991), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n767), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n774), .B1(new_n215), .B2(new_n312), .C1(new_n1008), .C2(new_n242), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n763), .ZN(new_n1010));
  INV_X1    g0810(.A(G317), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n326), .B1(new_n789), .B2(new_n1011), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n785), .A2(new_n860), .B1(new_n801), .B2(new_n226), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(G107), .C2(new_n779), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n807), .A2(new_n524), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n805), .A2(new_n499), .B1(KEYINPUT46), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(KEYINPUT46), .B2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(KEYINPUT113), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G303), .A2(new_n797), .B1(new_n799), .B2(new_n866), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1014), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1017), .A2(KEYINPUT113), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n804), .A2(G159), .B1(new_n850), .B2(G58), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n855), .B2(new_n785), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n801), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n326), .B1(new_n1024), .B2(G77), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1023), .B1(KEYINPUT114), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(KEYINPUT114), .B2(new_n1025), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n780), .A2(new_n203), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G137), .B2(new_n790), .ZN(new_n1029));
  INV_X1    g0829(.A(G150), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1029), .B1(new_n798), .B2(new_n265), .C1(new_n1030), .C2(new_n796), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1020), .A2(new_n1021), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT47), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1010), .B1(new_n1033), .B2(new_n773), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n995), .A2(new_n772), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1007), .A2(new_n1036), .ZN(G387));
  AND2_X1   g0837(.A1(new_n962), .A2(new_n963), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n955), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n696), .A2(new_n823), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G311), .A2(new_n804), .B1(new_n784), .B2(G322), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n536), .B2(new_n798), .C1(new_n1011), .C2(new_n796), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G294), .A2(new_n850), .B1(new_n779), .B2(new_n866), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT49), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n326), .B1(new_n789), .B2(new_n812), .C1(new_n524), .C2(new_n801), .ZN(new_n1052));
  OR3_X1    g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n856), .A2(new_n785), .B1(new_n805), .B2(new_n255), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n780), .A2(new_n312), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n799), .A2(G68), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n270), .B1(new_n789), .B2(new_n1030), .C1(new_n273), .C2(new_n807), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n797), .B2(G50), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n802), .A2(G97), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n844), .B1(new_n1053), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n775), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n603), .B1(new_n203), .B2(new_n273), .C1(new_n704), .C2(KEYINPUT115), .ZN(new_n1064));
  XOR2_X1   g0864(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n1065));
  OR3_X1    g0865(.A1(new_n1065), .A2(G50), .A3(new_n255), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(G50), .B2(new_n255), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n704), .A2(KEYINPUT115), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n767), .B1(new_n1064), .B2(new_n1069), .C1(new_n239), .C2(new_n330), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(G107), .B2(new_n215), .C1(new_n704), .C2(new_n764), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n762), .B(new_n1062), .C1(new_n1063), .C2(new_n1071), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT117), .Z(new_n1073));
  INV_X1    g0873(.A(new_n703), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n964), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1038), .A2(new_n758), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1040), .B1(new_n1041), .B2(new_n1073), .C1(new_n1075), .C2(new_n1076), .ZN(G393));
  OAI21_X1  g0877(.A(new_n774), .B1(new_n226), .B2(new_n215), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n767), .B2(new_n246), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n797), .A2(G159), .B1(G150), .B2(new_n784), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT51), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n799), .A2(new_n256), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n270), .B1(new_n789), .B2(new_n855), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G68), .B2(new_n850), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n804), .A2(G50), .B1(new_n779), .B2(G77), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n864), .A2(new_n1082), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n797), .A2(G311), .B1(G317), .B2(new_n784), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT52), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n270), .B1(new_n790), .B2(G322), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n807), .B2(new_n865), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n799), .A2(G294), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n804), .A2(G303), .B1(new_n779), .B2(G116), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n803), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1081), .A2(new_n1086), .B1(new_n1088), .B2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n762), .B(new_n1079), .C1(new_n1095), .C2(new_n773), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n969), .B2(new_n823), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n982), .B2(new_n955), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n983), .A2(new_n988), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n703), .B1(new_n964), .B2(new_n982), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G390));
  OAI21_X1  g0902(.A(new_n763), .B1(new_n256), .B2(new_n845), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n927), .A2(new_n771), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n270), .B(new_n808), .C1(G294), .C2(new_n790), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n226), .B2(new_n798), .C1(new_n524), .C2(new_n796), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n804), .A2(G107), .B1(new_n779), .B2(G77), .ZN(new_n1107));
  INV_X1    g0907(.A(G283), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n847), .B(new_n1107), .C1(new_n1108), .C2(new_n785), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n801), .A2(new_n265), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n326), .B(new_n1110), .C1(G125), .C2(new_n790), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT119), .Z(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n799), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1111), .B(new_n1114), .C1(new_n848), .C2(new_n796), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n807), .A2(new_n1030), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n784), .A2(G128), .B1(new_n779), .B2(G159), .ZN(new_n1119));
  INV_X1    g0919(.A(G137), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1119), .C1(new_n1120), .C2(new_n805), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1106), .A2(new_n1109), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1103), .B(new_n1104), .C1(new_n773), .C2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n675), .B1(new_n731), .B2(new_n935), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n945), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n929), .B1(new_n902), .B2(new_n907), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n915), .A2(new_n891), .B1(new_n916), .B2(new_n920), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n918), .A2(new_n921), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n410), .A2(new_n390), .A3(new_n890), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT38), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n910), .B1(new_n1132), .B2(new_n897), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n894), .A2(new_n895), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n912), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1135), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1127), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n716), .A2(new_n720), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1138), .B(new_n726), .C1(new_n659), .C2(new_n661), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(new_n685), .A3(new_n839), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n901), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n907), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n925), .A2(new_n896), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n928), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1126), .B1(new_n1137), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n755), .A2(G330), .A3(new_n945), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1142), .A2(new_n1143), .A3(new_n928), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n927), .C2(new_n1127), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1149), .A2(new_n955), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1123), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n452), .A2(new_n1124), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n931), .A2(new_n673), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n675), .B1(new_n731), .B2(new_n754), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n907), .B1(new_n1154), .B2(new_n839), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n902), .B1(new_n1126), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1141), .B1(new_n1154), .B2(new_n945), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1124), .A2(new_n839), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n906), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT118), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n900), .B1(new_n727), .B2(new_n839), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1146), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n907), .B1(new_n1124), .B2(new_n839), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT118), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1156), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1153), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n1149), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1153), .A2(new_n1166), .A3(new_n1148), .A4(new_n1145), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n1074), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1151), .A2(new_n1170), .ZN(G378));
  INV_X1    g0971(.A(new_n930), .ZN(new_n1172));
  XOR2_X1   g0972(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n306), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n269), .A2(new_n682), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT124), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n306), .A2(new_n1174), .ZN(new_n1180));
  OR3_X1    g0980(.A1(new_n1176), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1179), .B1(new_n1176), .B2(new_n1180), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n942), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n941), .B1(new_n1143), .B2(new_n940), .ZN(new_n1185));
  OAI211_X1 g0985(.A(G330), .B(new_n1183), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1183), .B1(new_n948), .B2(G330), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1172), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1183), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1143), .A2(new_n940), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT40), .B1(new_n1135), .B2(new_n896), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1191), .A2(KEYINPUT40), .B1(new_n1192), .B2(new_n940), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1190), .B1(new_n1193), .B2(new_n675), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(new_n930), .A3(new_n1186), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1189), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1190), .A2(new_n770), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n763), .B1(G50), .B2(new_n845), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n801), .A2(new_n202), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n805), .A2(new_n226), .B1(new_n273), .B2(new_n807), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G116), .C2(new_n784), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n329), .B(new_n326), .C1(new_n789), .C2(new_n1108), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1202), .B(new_n1028), .C1(G107), .C2(new_n797), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(new_n312), .C2(new_n798), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT122), .Z(new_n1205));
  INV_X1    g1005(.A(KEYINPUT58), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n265), .B1(G33), .B2(G41), .C1(new_n289), .C2(new_n270), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT121), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1113), .A2(new_n850), .B1(new_n797), .B2(G128), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n848), .B2(new_n805), .C1(new_n1120), .C2(new_n798), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n784), .A2(G125), .B1(new_n779), .B2(G150), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT123), .Z(new_n1214));
  NOR2_X1   g1014(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1216), .A2(KEYINPUT59), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(KEYINPUT59), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1024), .A2(G159), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G33), .B(G41), .C1(new_n790), .C2(G124), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1210), .B1(new_n1206), .B2(new_n1205), .C1(new_n1217), .C2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1198), .B1(new_n1222), .B2(new_n773), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1196), .A2(new_n1039), .B1(new_n1197), .B2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1195), .A2(new_n1189), .B1(new_n1169), .B2(new_n1153), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1074), .B1(new_n1225), .B2(KEYINPUT57), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT57), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1169), .B2(new_n1153), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1189), .A2(new_n1229), .A3(new_n1195), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1194), .A2(KEYINPUT125), .A3(new_n930), .A4(new_n1186), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1228), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1224), .B1(new_n1226), .B2(new_n1232), .ZN(G375));
  OAI21_X1  g1033(.A(new_n763), .B1(G68), .B2(new_n845), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n270), .B(new_n1055), .C1(G303), .C2(new_n790), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n320), .B2(new_n798), .C1(new_n1108), .C2(new_n796), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n802), .A2(G77), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n784), .A2(G294), .B1(new_n850), .B2(G97), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(new_n524), .C2(new_n805), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1113), .A2(new_n804), .B1(new_n799), .B2(G150), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n326), .B(new_n1199), .C1(G128), .C2(new_n790), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(new_n1120), .C2(new_n796), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n784), .A2(G132), .B1(new_n850), .B2(G159), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n265), .B2(new_n780), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1236), .A2(new_n1239), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1234), .B1(new_n1245), .B2(new_n773), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n907), .B2(new_n771), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1157), .A2(new_n1159), .A3(KEYINPUT118), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1164), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n906), .B1(new_n756), .B2(new_n835), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1125), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1248), .A2(new_n1249), .B1(new_n1251), .B2(new_n902), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1247), .B1(new_n1252), .B2(new_n955), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n931), .A2(new_n673), .A3(new_n1152), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(new_n990), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1253), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(G381));
  NOR3_X1   g1059(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n1101), .A3(new_n1258), .ZN(new_n1261));
  OR4_X1    g1061(.A1(G387), .A2(new_n1261), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1062(.A(G378), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n683), .A2(G213), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G407), .B(G213), .C1(G375), .C2(new_n1266), .ZN(G409));
  NAND2_X1  g1067(.A1(G387), .A2(new_n1101), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(new_n829), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1007), .A2(new_n1036), .A3(G390), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1269), .ZN(new_n1272));
  AOI21_X1  g1072(.A(G390), .B1(new_n1007), .B2(new_n1036), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1036), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1274), .B(new_n1101), .C1(new_n991), .C2(new_n1006), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1272), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1271), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G378), .B(new_n1224), .C1(new_n1226), .C2(new_n1232), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1230), .A2(new_n1231), .A3(new_n1039), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1169), .A2(new_n1153), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n990), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1196), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1197), .A2(new_n1223), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1280), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1263), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1265), .B1(new_n1279), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1265), .A2(G2897), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1252), .A2(KEYINPUT60), .A3(new_n1254), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1074), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT60), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1257), .B1(new_n1255), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1253), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(G384), .ZN(new_n1296));
  INV_X1    g1096(.A(G384), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1297), .B(new_n1253), .C1(new_n1292), .C2(new_n1294), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1289), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1167), .A2(KEYINPUT60), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1291), .B1(new_n1257), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1297), .B1(new_n1301), .B2(new_n1253), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1295), .A2(G384), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1288), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1299), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1278), .B1(new_n1287), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(KEYINPUT126), .B(new_n1278), .C1(new_n1287), .C2(new_n1305), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1279), .A2(new_n1286), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1312));
  OR2_X1    g1112(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1311), .A2(new_n1264), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1313), .B1(new_n1287), .B2(new_n1312), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1277), .B1(new_n1310), .B2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1277), .A2(new_n1306), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1287), .A2(new_n1312), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1321), .B(KEYINPUT63), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1319), .A2(new_n1323), .ZN(G405));
  NAND2_X1  g1124(.A1(G375), .A2(new_n1263), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1279), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n1312), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1327), .B(new_n1277), .ZN(G402));
endmodule


