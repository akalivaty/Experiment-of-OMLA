//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(G101), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G131), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n195), .A2(new_n198), .A3(new_n201), .A4(new_n196), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT64), .B1(new_n206), .B2(G143), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(new_n204), .A3(G146), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n205), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n204), .A2(G146), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n210), .A2(new_n211), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n203), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n197), .A2(G134), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n194), .A2(G137), .ZN(new_n219));
  OAI21_X1  g033(.A(G131), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n202), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  OAI21_X1  g036(.A(G128), .B1(new_n205), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n212), .A2(new_n213), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n226), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n210), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n221), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  OR2_X1    g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n232), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n217), .A2(new_n229), .A3(new_n235), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n236), .A2(KEYINPUT28), .ZN(new_n237));
  INV_X1    g051(.A(new_n235), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n228), .A2(new_n225), .ZN(new_n239));
  INV_X1    g053(.A(new_n221), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n203), .A2(new_n216), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n238), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT28), .B1(new_n243), .B2(new_n236), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n192), .B1(new_n237), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT30), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT65), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(KEYINPUT65), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n249), .B(new_n250), .C1(new_n217), .C2(new_n229), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT65), .A4(new_n247), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n236), .B1(new_n253), .B2(new_n235), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT31), .B1(new_n254), .B2(new_n192), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n238), .B1(new_n251), .B2(new_n252), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT31), .ZN(new_n257));
  INV_X1    g071(.A(new_n192), .ZN(new_n258));
  NOR4_X1   g072(.A1(new_n256), .A2(new_n257), .A3(new_n236), .A4(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n246), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G472), .A2(G902), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n260), .A2(KEYINPUT32), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT32), .B1(new_n260), .B2(new_n261), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n187), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n261), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT32), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n187), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G472), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT67), .B1(new_n254), .B2(new_n192), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n237), .A2(new_n244), .A3(new_n192), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n274), .B(new_n258), .C1(new_n256), .C2(new_n236), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n271), .A2(new_n272), .A3(new_n273), .A4(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n273), .A2(new_n272), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT69), .B(G902), .Z(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n270), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n269), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G119), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G128), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n226), .A2(G119), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT24), .B(G110), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G110), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n293), .B1(G119), .B2(new_n226), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n284), .A2(KEYINPUT23), .A3(G128), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n292), .B(new_n285), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n287), .A2(new_n288), .A3(KEYINPUT71), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n291), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT70), .B(G125), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT16), .ZN(new_n300));
  INV_X1    g114(.A(G140), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(G125), .A2(G140), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n303), .B1(new_n299), .B2(G140), .ZN(new_n304));
  OAI211_X1 g118(.A(G146), .B(new_n302), .C1(new_n304), .C2(new_n300), .ZN(new_n305));
  XNOR2_X1  g119(.A(G125), .B(G140), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n206), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n298), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n286), .A2(KEYINPUT23), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n293), .A2(new_n226), .A3(G119), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n309), .A2(new_n310), .B1(new_n284), .B2(G128), .ZN(new_n311));
  OAI22_X1  g125(.A1(new_n311), .A2(new_n292), .B1(new_n287), .B2(new_n288), .ZN(new_n312));
  INV_X1    g126(.A(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(G140), .ZN(new_n317));
  INV_X1    g131(.A(new_n303), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n300), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND4_X1   g133(.A1(new_n300), .A2(new_n314), .A3(new_n316), .A4(new_n301), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n206), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n312), .B1(new_n321), .B2(new_n305), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT73), .B1(new_n308), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n312), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n317), .A2(new_n318), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT16), .ZN(new_n326));
  AOI21_X1  g140(.A(G146), .B1(new_n326), .B2(new_n302), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n319), .A2(new_n206), .A3(new_n320), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n298), .A2(new_n305), .A3(new_n307), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G137), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT72), .ZN(new_n334));
  INV_X1    g148(.A(G221), .ZN(new_n335));
  INV_X1    g149(.A(G234), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n335), .A2(new_n336), .A3(G953), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n334), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n323), .A2(new_n332), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n329), .A2(new_n331), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(KEYINPUT73), .A3(new_n338), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n280), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G217), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(new_n344), .B2(G234), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n350), .A2(G902), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n343), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n283), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n203), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n208), .B1(new_n204), .B2(G146), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n206), .A2(KEYINPUT64), .A3(G143), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n212), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n359), .B1(new_n362), .B2(new_n223), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n210), .A2(KEYINPUT76), .A3(new_n227), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n228), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G104), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G107), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n366), .A2(G107), .ZN(new_n369));
  OAI21_X1  g183(.A(G101), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT3), .B1(new_n366), .B2(G107), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n372));
  INV_X1    g186(.A(G107), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(G104), .ZN(new_n374));
  INV_X1    g188(.A(G101), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n371), .A2(new_n374), .A3(new_n375), .A4(new_n367), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT10), .B1(new_n365), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n239), .A2(new_n378), .A3(KEYINPUT10), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n371), .A2(new_n374), .A3(new_n367), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n376), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n384), .A3(G101), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n216), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT79), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n362), .A2(new_n359), .A3(new_n223), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT76), .B1(new_n210), .B2(new_n227), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n390), .A2(new_n391), .B1(new_n227), .B2(new_n210), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n389), .B1(new_n392), .B2(new_n377), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n393), .A2(new_n394), .A3(new_n386), .A4(new_n380), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n358), .B1(new_n388), .B2(new_n395), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n379), .A2(new_n203), .A3(new_n387), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G140), .ZN(new_n398));
  INV_X1    g212(.A(G227), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G953), .ZN(new_n400));
  XOR2_X1   g214(.A(new_n398), .B(new_n400), .Z(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n396), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n397), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n239), .A2(new_n378), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n365), .B2(new_n378), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n358), .B1(new_n406), .B2(KEYINPUT78), .ZN(new_n407));
  INV_X1    g221(.A(new_n239), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n377), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n392), .B2(new_n377), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT12), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n390), .A2(new_n391), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n377), .B1(new_n414), .B2(new_n228), .ZN(new_n415));
  OAI211_X1 g229(.A(KEYINPUT12), .B(new_n203), .C1(new_n415), .C2(new_n405), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n410), .A2(KEYINPUT77), .A3(KEYINPUT12), .A4(new_n203), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n404), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n401), .B(KEYINPUT75), .Z(new_n422));
  AOI21_X1  g236(.A(new_n403), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G469), .ZN(new_n424));
  NAND2_X1  g238(.A1(G469), .A2(G902), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n397), .A2(new_n402), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n426), .B1(new_n413), .B2(new_n420), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n402), .B1(new_n396), .B2(new_n397), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G469), .ZN(new_n430));
  AND4_X1   g244(.A1(KEYINPUT80), .A2(new_n429), .A3(new_n430), .A4(new_n344), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n280), .B1(new_n427), .B2(new_n428), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT80), .B1(new_n432), .B2(new_n430), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n424), .B(new_n425), .C1(new_n431), .C2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n216), .A2(new_n299), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n408), .B2(new_n299), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n438), .A2(KEYINPUT7), .ZN(new_n439));
  INV_X1    g253(.A(G116), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G119), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G113), .B1(new_n442), .B2(KEYINPUT5), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n443), .A2(KEYINPUT81), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n232), .A2(KEYINPUT5), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n443), .B2(KEYINPUT81), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n234), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n378), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G122), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT8), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n445), .B(G113), .C1(KEYINPUT5), .C2(new_n442), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n234), .A3(new_n377), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n235), .A2(new_n385), .A3(new_n383), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n378), .A2(new_n234), .A3(new_n451), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n439), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n458));
  INV_X1    g272(.A(G953), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G224), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n438), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT7), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n438), .A2(KEYINPUT82), .A3(KEYINPUT7), .A4(new_n460), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n438), .A2(new_n460), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n457), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G902), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n461), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n454), .A2(new_n455), .ZN(new_n470));
  INV_X1    g284(.A(new_n449), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n474), .A3(new_n471), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n469), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n467), .A2(new_n468), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G210), .B1(G237), .B2(G902), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n467), .A2(new_n468), .A3(new_n478), .A4(new_n476), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n436), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT9), .B(G234), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n335), .B1(new_n484), .B2(new_n468), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n434), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G237), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n459), .A3(G214), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT84), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(G143), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n190), .A2(G214), .B1(new_n490), .B2(G143), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n492), .B1(new_n493), .B2(new_n491), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(KEYINPUT85), .ZN(new_n495));
  AND2_X1   g309(.A1(KEYINPUT18), .A2(G131), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n495), .B(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n307), .B1(new_n325), .B2(new_n206), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(G131), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n492), .B(new_n201), .C1(new_n493), .C2(new_n491), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT90), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n321), .B(new_n305), .C1(new_n501), .C2(new_n500), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(G113), .B(G122), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(G104), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(KEYINPUT89), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n499), .B(new_n510), .C1(new_n504), .C2(new_n505), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n468), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G475), .ZN(new_n514));
  INV_X1    g328(.A(G475), .ZN(new_n515));
  INV_X1    g329(.A(new_n508), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n317), .A2(KEYINPUT19), .A3(new_n318), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT19), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n306), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT87), .B1(new_n520), .B2(G146), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT87), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n517), .A2(new_n522), .A3(new_n206), .A4(new_n519), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n305), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT88), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n500), .A2(new_n502), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT86), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n527), .A2(KEYINPUT86), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n521), .A2(KEYINPUT88), .A3(new_n305), .A4(new_n523), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n526), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n516), .B1(new_n531), .B2(new_n499), .ZN(new_n532));
  INV_X1    g346(.A(new_n511), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n515), .B(new_n468), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n534), .A2(KEYINPUT20), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n514), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(G128), .B(G143), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT13), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n204), .A2(G128), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n541), .A2(KEYINPUT13), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(G134), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n194), .ZN(new_n545));
  INV_X1    g359(.A(G122), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G116), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n440), .A2(G122), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n373), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n373), .B1(new_n547), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n226), .A2(G143), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n541), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G134), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n555), .A2(new_n545), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT14), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n547), .A2(new_n548), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G107), .B1(new_n548), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n549), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI22_X1  g374(.A1(new_n544), .A2(new_n552), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n483), .A2(new_n349), .A3(G953), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n543), .B(new_n545), .C1(new_n551), .C2(new_n550), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n555), .A2(new_n545), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n566), .B(new_n549), .C1(new_n558), .C2(new_n559), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n567), .A3(new_n562), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n344), .ZN(new_n570));
  INV_X1    g384(.A(G478), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n571), .A2(KEYINPUT15), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n570), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G952), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(G953), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n336), .B2(new_n488), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n459), .B(new_n344), .C1(G234), .C2(G237), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT21), .B(G898), .Z(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n538), .A2(new_n574), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n357), .A2(new_n487), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G101), .ZN(G3));
  AND2_X1   g399(.A1(new_n434), .A2(new_n486), .ZN(new_n586));
  INV_X1    g400(.A(new_n356), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n260), .A2(new_n344), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G472), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n589), .A2(new_n265), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n586), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n561), .A2(new_n563), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n562), .B1(new_n565), .B2(new_n567), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT91), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT33), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n564), .B(new_n568), .C1(KEYINPUT91), .C2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(G478), .B(new_n344), .C1(new_n597), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT92), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n569), .B(KEYINPUT33), .C1(new_n595), .C2(new_n593), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n599), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT92), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(new_n605), .A3(G478), .A4(new_n344), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n570), .A2(new_n571), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n602), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT93), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n602), .A2(new_n606), .A3(KEYINPUT93), .A4(new_n607), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n538), .ZN(new_n613));
  INV_X1    g427(.A(new_n482), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n613), .A2(new_n614), .A3(new_n582), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n591), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT34), .B(G104), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  NOR2_X1   g433(.A1(new_n614), .A2(new_n582), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT94), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n513), .A2(new_n621), .A3(G475), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n509), .B2(new_n511), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT94), .B1(new_n623), .B2(new_n515), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n573), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n534), .B(new_n535), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n620), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n591), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT35), .B(G107), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NOR2_X1   g445(.A1(new_n339), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n341), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n353), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n352), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n590), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n487), .A3(new_n583), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT96), .B(KEYINPUT37), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n292), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n639), .B(new_n641), .ZN(G12));
  INV_X1    g456(.A(new_n635), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n253), .A2(new_n235), .ZN(new_n644));
  INV_X1    g458(.A(new_n236), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n645), .A3(new_n192), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n257), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n254), .A2(KEYINPUT31), .A3(new_n192), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n245), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n261), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n266), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n260), .A2(KEYINPUT32), .A3(new_n261), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n267), .B1(new_n653), .B2(new_n187), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n276), .A2(KEYINPUT68), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n276), .A2(KEYINPUT68), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n281), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G472), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n643), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n579), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n577), .B1(new_n660), .B2(G900), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n625), .A2(new_n626), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n487), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT97), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n226), .ZN(G30));
  OAI21_X1  g480(.A(new_n258), .B1(new_n243), .B2(new_n236), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT98), .B1(new_n646), .B2(new_n667), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n668), .A2(G902), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n646), .A2(KEYINPUT98), .A3(new_n667), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(KEYINPUT99), .B1(new_n654), .B2(new_n671), .ZN(new_n672));
  AND4_X1   g486(.A1(KEYINPUT99), .A2(new_n264), .A3(new_n268), .A4(new_n671), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n635), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n532), .A2(new_n533), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT20), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n515), .A4(new_n468), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n534), .A2(new_n535), .ZN(new_n679));
  AOI22_X1  g493(.A1(new_n678), .A2(new_n679), .B1(G475), .B2(new_n513), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n573), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n661), .B(KEYINPUT39), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n586), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT40), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n682), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n480), .A2(new_n481), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT38), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n436), .B1(new_n684), .B2(KEYINPUT40), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n675), .A2(new_n687), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n204), .ZN(G45));
  AND3_X1   g506(.A1(new_n612), .A2(new_n538), .A3(new_n661), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n487), .A2(new_n659), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NAND2_X1  g509(.A1(new_n432), .A2(new_n430), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT80), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n432), .A2(KEYINPUT80), .A3(new_n430), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n432), .A2(new_n430), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n486), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n357), .A2(new_n615), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT100), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n704), .B(new_n706), .ZN(G15));
  NAND3_X1  g521(.A1(new_n357), .A2(new_n627), .A3(new_n703), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NAND4_X1  g523(.A1(new_n700), .A2(new_n482), .A3(new_n486), .A4(new_n701), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n659), .A3(new_n583), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  NAND3_X1  g527(.A1(new_n538), .A2(new_n482), .A3(new_n574), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT103), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n538), .A2(new_n482), .A3(new_n716), .A4(new_n574), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n702), .A2(new_n582), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n237), .A2(new_n244), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n720), .A2(KEYINPUT101), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(KEYINPUT101), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n258), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n647), .A2(new_n648), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n650), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n589), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n588), .A2(KEYINPUT102), .A3(G472), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n718), .A2(new_n719), .A3(new_n587), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  INV_X1    g545(.A(new_n725), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT102), .B1(new_n588), .B2(G472), .ZN(new_n733));
  AOI211_X1 g547(.A(new_n726), .B(new_n270), .C1(new_n260), .C2(new_n344), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n635), .B(new_n732), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n612), .A2(new_n538), .A3(new_n661), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n710), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT104), .B(G125), .Z(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G27));
  XNOR2_X1  g553(.A(new_n425), .B(KEYINPUT105), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n424), .B(new_n740), .C1(new_n431), .C2(new_n433), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n486), .A2(new_n435), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n688), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n357), .A2(new_n693), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n653), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n356), .B1(new_n658), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n744), .A2(new_n749), .A3(KEYINPUT42), .A4(new_n693), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n750), .A2(KEYINPUT107), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(KEYINPUT107), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n747), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND3_X1  g568(.A1(new_n357), .A2(new_n663), .A3(new_n744), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n357), .A2(new_n757), .A3(new_n744), .A4(new_n663), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  OAI21_X1  g574(.A(G469), .B1(new_n423), .B2(KEYINPUT45), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n423), .A2(KEYINPUT45), .ZN(new_n764));
  OAI211_X1 g578(.A(KEYINPUT109), .B(G469), .C1(new_n423), .C2(KEYINPUT45), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT46), .B1(new_n766), .B2(new_n740), .ZN(new_n767));
  INV_X1    g581(.A(new_n700), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(KEYINPUT46), .A3(new_n740), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n486), .A3(new_n683), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n612), .A2(new_n680), .A3(KEYINPUT43), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT43), .B1(new_n612), .B2(new_n680), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n590), .B1(new_n776), .B2(KEYINPUT110), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n777), .B(new_n635), .C1(KEYINPUT110), .C2(new_n776), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n772), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n480), .A2(new_n435), .A3(new_n481), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n779), .B(new_n781), .C1(new_n773), .C2(new_n778), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  NAND2_X1  g597(.A1(new_n771), .A2(new_n486), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT47), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n486), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n736), .A2(new_n587), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n283), .A3(new_n781), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  XNOR2_X1  g605(.A(new_n573), .B(KEYINPUT111), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n680), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n613), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n794), .A2(new_n620), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(new_n587), .A3(new_n586), .A4(new_n590), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n639), .A2(new_n584), .A3(new_n730), .A4(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n704), .A2(new_n708), .A3(new_n712), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n792), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n781), .A2(new_n626), .A3(new_n661), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n659), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n622), .A2(new_n624), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n586), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n798), .A2(new_n800), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n753), .A2(new_n759), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n735), .A2(new_n736), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n744), .A2(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n352), .A2(new_n634), .A3(new_n661), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT112), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n352), .A2(new_n815), .A3(new_n634), .A4(new_n661), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n741), .A2(new_n817), .A3(new_n486), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n818), .B(new_n718), .C1(new_n672), .C2(new_n673), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n711), .A2(new_n810), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n664), .A3(new_n694), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT52), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n635), .B(new_n663), .C1(new_n269), .C2(new_n282), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n434), .A2(new_n482), .A3(new_n486), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n693), .A2(new_n729), .A3(new_n635), .ZN(new_n826));
  OAI22_X1  g640(.A1(new_n824), .A2(new_n825), .B1(new_n826), .B2(new_n710), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n635), .B1(new_n269), .B2(new_n282), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n828), .A2(new_n825), .A3(new_n736), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT113), .B1(new_n830), .B2(new_n819), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n821), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n823), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n812), .A2(KEYINPUT53), .A3(new_n822), .A4(new_n834), .ZN(new_n835));
  XOR2_X1   g649(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n797), .A2(new_n799), .A3(new_n806), .A4(new_n811), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n753), .A2(new_n759), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n821), .A2(new_n832), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n643), .B(new_n662), .C1(new_n654), .C2(new_n658), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n737), .B1(new_n487), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(KEYINPUT113), .A3(new_n694), .A4(new_n819), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n841), .A2(new_n844), .A3(KEYINPUT52), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT52), .B1(new_n841), .B2(new_n844), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT114), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n841), .A2(new_n844), .A3(KEYINPUT52), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n834), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n840), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n835), .B(new_n837), .C1(new_n851), .C2(KEYINPUT53), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(KEYINPUT53), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n812), .A2(new_n822), .A3(new_n834), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n853), .B1(KEYINPUT54), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n729), .A2(new_n587), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT116), .B1(new_n776), .B2(new_n577), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n862), .B(new_n578), .C1(new_n774), .C2(new_n775), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n860), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n864), .A2(new_n781), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n786), .A2(KEYINPUT117), .A3(new_n787), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n700), .A2(new_n701), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n485), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT117), .B1(new_n786), .B2(new_n787), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n867), .A2(new_n743), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n861), .B2(new_n863), .ZN(new_n873));
  INV_X1    g687(.A(new_n735), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n872), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n674), .A2(new_n876), .A3(new_n587), .A4(new_n578), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n680), .A2(new_n610), .A3(new_n611), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT50), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT118), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n702), .B(new_n860), .C1(new_n861), .C2(new_n863), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n689), .A2(new_n435), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND4_X1   g699(.A1(new_n703), .A2(new_n864), .A3(new_n882), .A4(new_n884), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n875), .B(new_n880), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT51), .B1(new_n871), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n786), .A2(new_n787), .A3(new_n868), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n865), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT51), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n576), .B1(new_n892), .B2(new_n887), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n873), .A2(new_n749), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT48), .Z(new_n895));
  NOR2_X1   g709(.A1(new_n877), .A2(new_n613), .ZN(new_n896));
  NOR4_X1   g710(.A1(new_n889), .A2(new_n893), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n864), .A2(new_n711), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n859), .A2(KEYINPUT119), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n858), .A2(KEYINPUT54), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n897), .A3(new_n852), .A4(new_n898), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n575), .A2(new_n459), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT49), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n673), .B(new_n672), .C1(new_n906), .C2(new_n867), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n612), .A2(new_n680), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n867), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n689), .B(new_n742), .C1(new_n910), .C2(KEYINPUT49), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n907), .A2(new_n587), .A3(new_n909), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n905), .A2(new_n912), .ZN(G75));
  AND2_X1   g727(.A1(new_n473), .A2(new_n475), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(new_n469), .Z(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n835), .B1(new_n851), .B2(KEYINPUT53), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n280), .A3(new_n479), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT55), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(KEYINPUT56), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n918), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n918), .A2(new_n921), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT55), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n915), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n459), .A2(G952), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n924), .A2(new_n928), .A3(new_n930), .ZN(G51));
  NAND2_X1  g745(.A1(new_n740), .A2(KEYINPUT57), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n740), .A2(KEYINPUT57), .ZN(new_n933));
  INV_X1    g747(.A(new_n917), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n837), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n932), .B(new_n933), .C1(new_n935), .C2(new_n853), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n429), .ZN(new_n937));
  OR3_X1    g751(.A1(new_n934), .A2(new_n344), .A3(new_n766), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n929), .B1(new_n937), .B2(new_n938), .ZN(G54));
  AND2_X1   g753(.A1(KEYINPUT58), .A2(G475), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n917), .A2(new_n280), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n676), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n929), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n917), .A2(new_n280), .A3(new_n676), .A4(new_n940), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT122), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(KEYINPUT122), .B(new_n943), .C1(new_n945), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(G60));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT59), .Z(new_n953));
  OAI211_X1 g767(.A(new_n599), .B(new_n603), .C1(new_n859), .C2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n953), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n604), .B(new_n955), .C1(new_n935), .C2(new_n853), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n954), .A2(new_n930), .A3(new_n956), .ZN(G63));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT123), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT60), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n633), .B(KEYINPUT124), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n917), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n963), .A3(new_n930), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT61), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n917), .A2(new_n960), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n930), .B(new_n962), .C1(new_n966), .C2(new_n343), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G66));
  AOI21_X1  g782(.A(new_n459), .B1(new_n580), .B2(G224), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n798), .A2(new_n800), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n459), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT126), .ZN(new_n972));
  INV_X1    g786(.A(G898), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n914), .B1(new_n973), .B2(G953), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n972), .B(new_n974), .ZN(G69));
  INV_X1    g789(.A(new_n830), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n691), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT62), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n782), .A2(new_n790), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n685), .A2(new_n357), .A3(new_n781), .A4(new_n794), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n459), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n253), .B(new_n520), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n459), .A2(G900), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n772), .B1(new_n717), .B2(new_n715), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n976), .B1(new_n986), .B2(new_n749), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n979), .A2(new_n839), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n985), .B1(new_n988), .B2(new_n459), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n984), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n459), .B1(G227), .B2(G900), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT127), .Z(new_n992));
  XNOR2_X1  g806(.A(new_n990), .B(new_n992), .ZN(G72));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n981), .B2(new_n970), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n996), .B(new_n192), .C1(new_n236), .C2(new_n256), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n995), .B1(new_n988), .B2(new_n970), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n258), .A3(new_n254), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n997), .A2(new_n930), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n271), .A2(new_n646), .A3(new_n275), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n858), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1000), .B1(new_n995), .B2(new_n1002), .ZN(G57));
endmodule


