

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754;

  XNOR2_X2 U363 ( .A(n393), .B(G134), .ZN(n543) );
  XNOR2_X2 U364 ( .A(n413), .B(G128), .ZN(n393) );
  NAND2_X2 U365 ( .A1(n354), .A2(n423), .ZN(n361) );
  NAND2_X1 U366 ( .A1(n654), .A2(n752), .ZN(n634) );
  NAND2_X1 U367 ( .A1(n456), .A2(n455), .ZN(n460) );
  OR2_X1 U368 ( .A1(n631), .A2(n632), .ZN(n434) );
  XNOR2_X1 U369 ( .A(n562), .B(KEYINPUT19), .ZN(n600) );
  NAND2_X1 U370 ( .A1(n368), .A2(n687), .ZN(n562) );
  XNOR2_X1 U371 ( .A(n565), .B(KEYINPUT1), .ZN(n674) );
  NAND2_X1 U372 ( .A1(n389), .A2(n386), .ZN(n565) );
  XNOR2_X1 U373 ( .A(n425), .B(n347), .ZN(n368) );
  AND2_X1 U374 ( .A1(n391), .A2(n390), .ZN(n389) );
  XNOR2_X1 U375 ( .A(n735), .B(G146), .ZN(n552) );
  XNOR2_X1 U376 ( .A(n543), .B(n410), .ZN(n735) );
  NAND2_X1 U377 ( .A1(n483), .A2(n482), .ZN(n499) );
  XNOR2_X1 U378 ( .A(n407), .B(G953), .ZN(n504) );
  INV_X1 U379 ( .A(G143), .ZN(n413) );
  INV_X1 U380 ( .A(KEYINPUT64), .ZN(n407) );
  BUF_X1 U381 ( .A(n747), .Z(n342) );
  XNOR2_X2 U382 ( .A(n361), .B(KEYINPUT2), .ZN(n343) );
  XNOR2_X1 U383 ( .A(n361), .B(KEYINPUT2), .ZN(n360) );
  XNOR2_X1 U384 ( .A(n403), .B(KEYINPUT20), .ZN(n511) );
  INV_X1 U385 ( .A(n751), .ZN(n385) );
  AND2_X1 U386 ( .A1(n457), .A2(n618), .ZN(n454) );
  NAND2_X1 U387 ( .A1(n392), .A2(G902), .ZN(n390) );
  BUF_X1 U388 ( .A(n565), .Z(n401) );
  XNOR2_X1 U389 ( .A(G902), .B(KEYINPUT15), .ZN(n489) );
  AND2_X1 U390 ( .A1(n741), .A2(n636), .ZN(n451) );
  NOR2_X1 U391 ( .A1(G953), .A2(G237), .ZN(n517) );
  XOR2_X1 U392 ( .A(G122), .B(G104), .Z(n525) );
  INV_X1 U393 ( .A(n669), .ZN(n383) );
  AND2_X1 U394 ( .A1(n348), .A2(n583), .ZN(n378) );
  AND2_X1 U395 ( .A1(n584), .A2(n383), .ZN(n376) );
  AND2_X1 U396 ( .A1(n457), .A2(n458), .ZN(n443) );
  XNOR2_X1 U397 ( .A(n730), .B(n486), .ZN(n549) );
  XNOR2_X1 U398 ( .A(n365), .B(n364), .ZN(n363) );
  XNOR2_X1 U399 ( .A(n367), .B(n366), .ZN(n365) );
  XNOR2_X1 U400 ( .A(KEYINPUT18), .B(KEYINPUT81), .ZN(n367) );
  BUF_X1 U401 ( .A(n674), .Z(n405) );
  XNOR2_X1 U402 ( .A(n510), .B(n345), .ZN(n370) );
  XOR2_X1 U403 ( .A(n563), .B(KEYINPUT6), .Z(n623) );
  XNOR2_X1 U404 ( .A(n479), .B(n478), .ZN(n521) );
  XOR2_X1 U405 ( .A(KEYINPUT3), .B(G116), .Z(n478) );
  XNOR2_X1 U406 ( .A(n477), .B(n476), .ZN(n479) );
  INV_X1 U407 ( .A(G119), .ZN(n476) );
  XNOR2_X1 U408 ( .A(KEYINPUT23), .B(KEYINPUT97), .ZN(n501) );
  XNOR2_X1 U409 ( .A(n437), .B(n500), .ZN(n441) );
  XNOR2_X1 U410 ( .A(n499), .B(n438), .ZN(n437) );
  INV_X1 U411 ( .A(G140), .ZN(n438) );
  XNOR2_X1 U412 ( .A(G119), .B(G128), .ZN(n507) );
  XNOR2_X1 U413 ( .A(n579), .B(n408), .ZN(n586) );
  INV_X1 U414 ( .A(KEYINPUT39), .ZN(n408) );
  OR2_X1 U415 ( .A1(n372), .A2(n346), .ZN(n576) );
  INV_X1 U416 ( .A(KEYINPUT28), .ZN(n373) );
  XNOR2_X1 U417 ( .A(n406), .B(n536), .ZN(n568) );
  NOR2_X1 U418 ( .A1(n716), .A2(G902), .ZN(n406) );
  NOR2_X1 U419 ( .A1(n398), .A2(n723), .ZN(n397) );
  NOR2_X1 U420 ( .A1(n472), .A2(n444), .ZN(n398) );
  NAND2_X1 U421 ( .A1(n395), .A2(n717), .ZN(n394) );
  NOR2_X1 U422 ( .A1(n637), .A2(n449), .ZN(n448) );
  INV_X1 U423 ( .A(G210), .ZN(n449) );
  XNOR2_X1 U424 ( .A(n643), .B(n642), .ZN(n644) );
  XOR2_X1 U425 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n527) );
  NAND2_X1 U426 ( .A1(n553), .A2(n388), .ZN(n387) );
  INV_X1 U427 ( .A(G902), .ZN(n388) );
  NOR2_X1 U428 ( .A1(n461), .A2(KEYINPUT89), .ZN(n458) );
  INV_X1 U429 ( .A(G146), .ZN(n481) );
  XNOR2_X1 U430 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n512), .B(KEYINPUT21), .ZN(n556) );
  XNOR2_X1 U432 ( .A(G113), .B(G101), .ZN(n477) );
  NAND2_X1 U433 ( .A1(G234), .A2(G237), .ZN(n492) );
  OR2_X1 U434 ( .A1(G237), .A2(G902), .ZN(n491) );
  XNOR2_X1 U435 ( .A(n736), .B(n349), .ZN(n531) );
  XNOR2_X1 U436 ( .A(G113), .B(G143), .ZN(n524) );
  XNOR2_X1 U437 ( .A(n521), .B(n520), .ZN(n422) );
  NAND2_X1 U438 ( .A1(n378), .A2(n376), .ZN(n375) );
  INV_X1 U439 ( .A(G953), .ZN(n724) );
  XNOR2_X1 U440 ( .A(G116), .B(G107), .ZN(n537) );
  NOR2_X1 U441 ( .A1(n637), .A2(n445), .ZN(n444) );
  INV_X1 U442 ( .A(G475), .ZN(n445) );
  XNOR2_X1 U443 ( .A(n414), .B(n549), .ZN(n551) );
  XNOR2_X1 U444 ( .A(n550), .B(n475), .ZN(n414) );
  XNOR2_X1 U445 ( .A(n488), .B(n729), .ZN(n641) );
  XNOR2_X1 U446 ( .A(n487), .B(n549), .ZN(n488) );
  XNOR2_X1 U447 ( .A(n424), .B(n363), .ZN(n487) );
  BUF_X1 U448 ( .A(n686), .Z(n703) );
  INV_X1 U449 ( .A(n615), .ZN(n468) );
  NAND2_X1 U450 ( .A1(n465), .A2(n473), .ZN(n464) );
  NOR2_X1 U451 ( .A1(n560), .A2(n559), .ZN(n578) );
  AND2_X1 U452 ( .A1(n450), .A2(n446), .ZN(n357) );
  NOR2_X1 U453 ( .A1(n637), .A2(n447), .ZN(n446) );
  INV_X1 U454 ( .A(G472), .ZN(n447) );
  BUF_X1 U455 ( .A(n504), .Z(n743) );
  XNOR2_X1 U456 ( .A(n485), .B(G107), .ZN(n730) );
  XNOR2_X1 U457 ( .A(G104), .B(G110), .ZN(n485) );
  XNOR2_X1 U458 ( .A(n521), .B(n404), .ZN(n729) );
  XNOR2_X1 U459 ( .A(KEYINPUT16), .B(G122), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n440), .B(n439), .ZN(n722) );
  XNOR2_X1 U461 ( .A(n509), .B(n503), .ZN(n439) );
  AND2_X1 U462 ( .A1(n450), .A2(n356), .ZN(n355) );
  NOR2_X1 U463 ( .A1(n586), .A2(n580), .ZN(n581) );
  XNOR2_X1 U464 ( .A(n555), .B(KEYINPUT113), .ZN(n751) );
  XNOR2_X1 U465 ( .A(n630), .B(KEYINPUT32), .ZN(n426) );
  OR2_X1 U466 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U467 ( .A(n580), .B(KEYINPUT107), .ZN(n660) );
  NOR2_X1 U468 ( .A1(n576), .A2(n566), .ZN(n567) );
  NOR2_X1 U469 ( .A1(n563), .A2(n672), .ZN(n427) );
  INV_X1 U470 ( .A(n660), .ZN(n663) );
  INV_X1 U471 ( .A(KEYINPUT87), .ZN(n412) );
  INV_X1 U472 ( .A(KEYINPUT60), .ZN(n470) );
  NAND2_X1 U473 ( .A1(n396), .A2(n394), .ZN(n400) );
  AND2_X1 U474 ( .A1(n399), .A2(n397), .ZN(n396) );
  INV_X1 U475 ( .A(KEYINPUT56), .ZN(n416) );
  NOR2_X1 U476 ( .A1(G953), .A2(n708), .ZN(n710) );
  XNOR2_X2 U477 ( .A(n523), .B(n522), .ZN(n563) );
  AND2_X1 U478 ( .A1(n450), .A2(n350), .ZN(n344) );
  XNOR2_X1 U479 ( .A(KEYINPUT25), .B(KEYINPUT98), .ZN(n345) );
  XOR2_X1 U480 ( .A(n401), .B(KEYINPUT111), .Z(n346) );
  XNOR2_X1 U481 ( .A(n490), .B(KEYINPUT85), .ZN(n347) );
  AND2_X1 U482 ( .A1(n385), .A2(n384), .ZN(n348) );
  XOR2_X1 U483 ( .A(n530), .B(n528), .Z(n349) );
  XNOR2_X1 U484 ( .A(n629), .B(n426), .ZN(n752) );
  AND2_X1 U485 ( .A1(n472), .A2(n444), .ZN(n350) );
  XNOR2_X1 U486 ( .A(KEYINPUT59), .B(KEYINPUT67), .ZN(n351) );
  XOR2_X1 U487 ( .A(n639), .B(KEYINPUT114), .Z(n352) );
  INV_X1 U488 ( .A(n717), .ZN(n472) );
  XNOR2_X1 U489 ( .A(n716), .B(n351), .ZN(n717) );
  NOR2_X1 U490 ( .A1(n743), .A2(G952), .ZN(n723) );
  INV_X1 U491 ( .A(n723), .ZN(n471) );
  OR2_X1 U492 ( .A1(n711), .A2(n387), .ZN(n386) );
  XNOR2_X1 U493 ( .A(n552), .B(n422), .ZN(n638) );
  XNOR2_X1 U494 ( .A(n552), .B(n551), .ZN(n711) );
  XNOR2_X1 U495 ( .A(n441), .B(n442), .ZN(n440) );
  INV_X1 U496 ( .A(n441), .ZN(n736) );
  NAND2_X1 U497 ( .A1(n504), .A2(G224), .ZN(n364) );
  XNOR2_X1 U498 ( .A(n714), .B(n715), .ZN(n402) );
  NAND2_X1 U499 ( .A1(n353), .A2(G469), .ZN(n714) );
  NAND2_X1 U500 ( .A1(n353), .A2(G217), .ZN(n721) );
  NAND2_X1 U501 ( .A1(n353), .A2(G478), .ZN(n719) );
  AND2_X2 U502 ( .A1(n355), .A2(n343), .ZN(n353) );
  NAND2_X1 U503 ( .A1(n354), .A2(n451), .ZN(n450) );
  NAND2_X1 U504 ( .A1(n354), .A2(n724), .ZN(n728) );
  XNOR2_X2 U505 ( .A(n436), .B(KEYINPUT45), .ZN(n354) );
  NAND2_X1 U506 ( .A1(n360), .A2(n450), .ZN(n395) );
  NAND2_X1 U507 ( .A1(n343), .A2(n344), .ZN(n399) );
  INV_X1 U508 ( .A(n637), .ZN(n356) );
  NAND2_X1 U509 ( .A1(n360), .A2(n357), .ZN(n453) );
  NAND2_X1 U510 ( .A1(n343), .A2(n358), .ZN(n645) );
  AND2_X1 U511 ( .A1(n450), .A2(n448), .ZN(n358) );
  NAND2_X1 U512 ( .A1(n359), .A2(G221), .ZN(n442) );
  NAND2_X1 U513 ( .A1(n359), .A2(G217), .ZN(n539) );
  XNOR2_X2 U514 ( .A(n505), .B(n506), .ZN(n359) );
  NOR2_X2 U515 ( .A1(n362), .A2(n674), .ZN(n608) );
  NOR2_X1 U516 ( .A1(n362), .A2(n401), .ZN(n614) );
  NAND2_X1 U517 ( .A1(n362), .A2(n405), .ZN(n675) );
  XNOR2_X2 U518 ( .A(n369), .B(KEYINPUT69), .ZN(n362) );
  INV_X1 U519 ( .A(n368), .ZN(n592) );
  XNOR2_X1 U520 ( .A(n592), .B(KEYINPUT38), .ZN(n688) );
  NAND2_X1 U521 ( .A1(n578), .A2(n368), .ZN(n561) );
  NOR2_X2 U522 ( .A1(n624), .A2(n556), .ZN(n369) );
  XNOR2_X2 U523 ( .A(n371), .B(n370), .ZN(n624) );
  OR2_X2 U524 ( .A1(n722), .A2(G902), .ZN(n371) );
  XNOR2_X1 U525 ( .A(n400), .B(n470), .ZN(G60) );
  XNOR2_X1 U526 ( .A(n374), .B(n373), .ZN(n372) );
  AND2_X1 U527 ( .A1(n564), .A2(n563), .ZN(n374) );
  NAND2_X1 U528 ( .A1(n377), .A2(n375), .ZN(n594) );
  NAND2_X1 U529 ( .A1(n379), .A2(n383), .ZN(n377) );
  NAND2_X1 U530 ( .A1(n382), .A2(n380), .ZN(n379) );
  NAND2_X1 U531 ( .A1(n381), .A2(n585), .ZN(n380) );
  NAND2_X1 U532 ( .A1(n583), .A2(n385), .ZN(n381) );
  OR2_X1 U533 ( .A1(n584), .A2(n384), .ZN(n382) );
  INV_X1 U534 ( .A(n585), .ZN(n384) );
  NAND2_X1 U535 ( .A1(n711), .A2(n392), .ZN(n391) );
  INV_X1 U536 ( .A(n553), .ZN(n392) );
  XNOR2_X1 U537 ( .A(n484), .B(n393), .ZN(n424) );
  NOR2_X1 U538 ( .A1(n402), .A2(n723), .ZN(G54) );
  NAND2_X1 U539 ( .A1(n637), .A2(G234), .ZN(n403) );
  NAND2_X1 U540 ( .A1(n504), .A2(G234), .ZN(n505) );
  NOR2_X1 U541 ( .A1(n587), .A2(n562), .ZN(n547) );
  NAND2_X1 U542 ( .A1(n409), .A2(KEYINPUT89), .ZN(n456) );
  NAND2_X1 U543 ( .A1(n619), .A2(n454), .ZN(n409) );
  INV_X1 U544 ( .A(n516), .ZN(n410) );
  NAND2_X1 U545 ( .A1(n600), .A2(n601), .ZN(n602) );
  NAND2_X1 U546 ( .A1(n411), .A2(n672), .ZN(n457) );
  XNOR2_X1 U547 ( .A(n607), .B(n412), .ZN(n411) );
  NAND2_X1 U548 ( .A1(n415), .A2(n434), .ZN(n433) );
  NAND2_X1 U549 ( .A1(n418), .A2(n635), .ZN(n415) );
  NAND2_X1 U550 ( .A1(n747), .A2(KEYINPUT44), .ZN(n619) );
  XNOR2_X1 U551 ( .A(n453), .B(n352), .ZN(n452) );
  XNOR2_X1 U552 ( .A(n417), .B(n416), .ZN(G51) );
  NAND2_X1 U553 ( .A1(n646), .A2(n471), .ZN(n417) );
  XNOR2_X1 U554 ( .A(n633), .B(KEYINPUT68), .ZN(n418) );
  NAND2_X1 U555 ( .A1(n614), .A2(n419), .ZN(n559) );
  XNOR2_X1 U556 ( .A(n557), .B(n558), .ZN(n419) );
  NOR2_X1 U557 ( .A1(n420), .A2(n723), .ZN(G66) );
  XNOR2_X1 U558 ( .A(n722), .B(n721), .ZN(n420) );
  NOR2_X1 U559 ( .A1(n421), .A2(n723), .ZN(G63) );
  XNOR2_X1 U560 ( .A(n719), .B(n720), .ZN(n421) );
  NOR2_X1 U561 ( .A1(n741), .A2(n636), .ZN(n423) );
  NAND2_X1 U562 ( .A1(n641), .A2(n637), .ZN(n425) );
  NAND2_X1 U563 ( .A1(n634), .A2(KEYINPUT44), .ZN(n631) );
  NAND2_X1 U564 ( .A1(n622), .A2(n427), .ZN(n654) );
  XNOR2_X2 U565 ( .A(n428), .B(n609), .ZN(n686) );
  NAND2_X1 U566 ( .A1(n429), .A2(n623), .ZN(n428) );
  XNOR2_X1 U567 ( .A(n459), .B(KEYINPUT106), .ZN(n429) );
  XNOR2_X2 U568 ( .A(n608), .B(KEYINPUT78), .ZN(n459) );
  NAND2_X1 U569 ( .A1(n432), .A2(n430), .ZN(n436) );
  NAND2_X1 U570 ( .A1(n460), .A2(n431), .ZN(n430) );
  AND2_X1 U571 ( .A1(n631), .A2(n632), .ZN(n431) );
  NOR2_X1 U572 ( .A1(n435), .A2(n433), .ZN(n432) );
  NOR2_X1 U573 ( .A1(n460), .A2(n632), .ZN(n435) );
  NAND2_X1 U574 ( .A1(n619), .A2(n443), .ZN(n455) );
  NOR2_X1 U575 ( .A1(n466), .A2(n464), .ZN(n463) );
  XNOR2_X2 U576 ( .A(n489), .B(KEYINPUT92), .ZN(n637) );
  NAND2_X1 U577 ( .A1(n452), .A2(n471), .ZN(n640) );
  INV_X1 U578 ( .A(n457), .ZN(n647) );
  NAND2_X1 U579 ( .A1(n459), .A2(n563), .ZN(n681) );
  INV_X1 U580 ( .A(n618), .ZN(n461) );
  NAND2_X1 U581 ( .A1(n463), .A2(n462), .ZN(n469) );
  NAND2_X1 U582 ( .A1(n686), .A2(n611), .ZN(n462) );
  NAND2_X1 U583 ( .A1(n615), .A2(n611), .ZN(n465) );
  NOR2_X1 U584 ( .A1(n686), .A2(n467), .ZN(n466) );
  NAND2_X1 U585 ( .A1(n468), .A2(n610), .ZN(n467) );
  XNOR2_X2 U586 ( .A(n469), .B(KEYINPUT35), .ZN(n747) );
  XNOR2_X1 U587 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X2 U588 ( .A(n602), .B(KEYINPUT0), .ZN(n615) );
  XOR2_X1 U589 ( .A(n612), .B(KEYINPUT82), .Z(n473) );
  XOR2_X1 U590 ( .A(KEYINPUT66), .B(KEYINPUT22), .Z(n474) );
  XOR2_X1 U591 ( .A(n548), .B(KEYINPUT80), .Z(n475) );
  INV_X1 U592 ( .A(KEYINPUT5), .ZN(n518) );
  XNOR2_X1 U593 ( .A(n519), .B(n518), .ZN(n520) );
  INV_X1 U594 ( .A(n690), .ZN(n603) );
  INV_X1 U595 ( .A(KEYINPUT88), .ZN(n632) );
  INV_X1 U596 ( .A(n623), .ZN(n626) );
  INV_X1 U597 ( .A(G125), .ZN(n480) );
  NAND2_X1 U598 ( .A1(G146), .A2(n480), .ZN(n483) );
  NAND2_X1 U599 ( .A1(n481), .A2(G125), .ZN(n482) );
  INV_X1 U600 ( .A(n499), .ZN(n484) );
  XNOR2_X1 U601 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n486) );
  NAND2_X1 U602 ( .A1(n491), .A2(G210), .ZN(n490) );
  NAND2_X1 U603 ( .A1(G214), .A2(n491), .ZN(n687) );
  XNOR2_X1 U604 ( .A(n492), .B(KEYINPUT14), .ZN(n493) );
  NAND2_X1 U605 ( .A1(G952), .A2(n493), .ZN(n702) );
  NOR2_X1 U606 ( .A1(G953), .A2(n702), .ZN(n598) );
  NAND2_X1 U607 ( .A1(n493), .A2(G902), .ZN(n494) );
  XNOR2_X1 U608 ( .A(n494), .B(KEYINPUT93), .ZN(n595) );
  INV_X1 U609 ( .A(n595), .ZN(n495) );
  NOR2_X1 U610 ( .A1(n743), .A2(n495), .ZN(n496) );
  XOR2_X1 U611 ( .A(KEYINPUT108), .B(n496), .Z(n497) );
  NOR2_X1 U612 ( .A1(G900), .A2(n497), .ZN(n498) );
  NOR2_X1 U613 ( .A1(n598), .A2(n498), .ZN(n560) );
  XOR2_X1 U614 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n500) );
  XOR2_X1 U615 ( .A(KEYINPUT96), .B(KEYINPUT24), .Z(n502) );
  XNOR2_X1 U616 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U617 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n506) );
  XOR2_X1 U618 ( .A(G110), .B(G137), .Z(n508) );
  XOR2_X1 U619 ( .A(n508), .B(n507), .Z(n509) );
  NAND2_X1 U620 ( .A1(n511), .A2(G217), .ZN(n510) );
  NAND2_X1 U621 ( .A1(n511), .A2(G221), .ZN(n512) );
  INV_X1 U622 ( .A(n556), .ZN(n671) );
  NAND2_X1 U623 ( .A1(n624), .A2(n671), .ZN(n513) );
  NOR2_X1 U624 ( .A1(n560), .A2(n513), .ZN(n564) );
  XOR2_X1 U625 ( .A(KEYINPUT4), .B(G137), .Z(n515) );
  XNOR2_X1 U626 ( .A(G131), .B(KEYINPUT72), .ZN(n514) );
  XNOR2_X1 U627 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U628 ( .A(KEYINPUT79), .B(n517), .Z(n529) );
  NAND2_X1 U629 ( .A1(n529), .A2(G210), .ZN(n519) );
  NOR2_X1 U630 ( .A1(G902), .A2(n638), .ZN(n523) );
  XNOR2_X1 U631 ( .A(G472), .B(KEYINPUT77), .ZN(n522) );
  XNOR2_X1 U632 ( .A(n525), .B(n524), .ZN(n532) );
  XNOR2_X1 U633 ( .A(G131), .B(KEYINPUT99), .ZN(n526) );
  XNOR2_X1 U634 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U635 ( .A1(G214), .A2(n529), .ZN(n530) );
  XNOR2_X1 U636 ( .A(n532), .B(n531), .ZN(n716) );
  XOR2_X1 U637 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n534) );
  XNOR2_X1 U638 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n533) );
  XNOR2_X1 U639 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U640 ( .A(G475), .B(n535), .ZN(n536) );
  XOR2_X1 U641 ( .A(KEYINPUT7), .B(G122), .Z(n538) );
  XNOR2_X1 U642 ( .A(n538), .B(n537), .ZN(n542) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n540) );
  XNOR2_X1 U644 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U645 ( .A(n542), .B(n541), .ZN(n544) );
  XNOR2_X1 U646 ( .A(n543), .B(n544), .ZN(n718) );
  NOR2_X1 U647 ( .A1(G902), .A2(n718), .ZN(n545) );
  XNOR2_X1 U648 ( .A(G478), .B(n545), .ZN(n573) );
  NAND2_X1 U649 ( .A1(n568), .A2(n573), .ZN(n580) );
  AND2_X1 U650 ( .A1(n623), .A2(n660), .ZN(n546) );
  NAND2_X1 U651 ( .A1(n564), .A2(n546), .ZN(n587) );
  XNOR2_X1 U652 ( .A(KEYINPUT36), .B(n547), .ZN(n554) );
  XNOR2_X1 U653 ( .A(G101), .B(G140), .ZN(n548) );
  NAND2_X1 U654 ( .A1(n743), .A2(G227), .ZN(n550) );
  XNOR2_X1 U655 ( .A(KEYINPUT74), .B(G469), .ZN(n553) );
  INV_X1 U656 ( .A(n405), .ZN(n620) );
  NAND2_X1 U657 ( .A1(n554), .A2(n620), .ZN(n555) );
  INV_X1 U658 ( .A(n568), .ZN(n572) );
  OR2_X1 U659 ( .A1(n573), .A2(n572), .ZN(n612) );
  XOR2_X1 U660 ( .A(KEYINPUT30), .B(KEYINPUT110), .Z(n558) );
  NAND2_X1 U661 ( .A1(n563), .A2(n687), .ZN(n557) );
  NOR2_X1 U662 ( .A1(n612), .A2(n561), .ZN(n658) );
  INV_X1 U663 ( .A(n600), .ZN(n566) );
  XNOR2_X1 U664 ( .A(n567), .B(KEYINPUT84), .ZN(n661) );
  NOR2_X1 U665 ( .A1(n568), .A2(n573), .ZN(n569) );
  XOR2_X1 U666 ( .A(KEYINPUT104), .B(n569), .Z(n667) );
  NAND2_X1 U667 ( .A1(n667), .A2(n580), .ZN(n691) );
  NAND2_X1 U668 ( .A1(n661), .A2(n691), .ZN(n570) );
  XNOR2_X1 U669 ( .A(KEYINPUT47), .B(n570), .ZN(n571) );
  NOR2_X1 U670 ( .A1(n658), .A2(n571), .ZN(n584) );
  NAND2_X1 U671 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U672 ( .A1(n573), .A2(n572), .ZN(n690) );
  NOR2_X1 U673 ( .A1(n692), .A2(n690), .ZN(n575) );
  XNOR2_X1 U674 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n574) );
  XNOR2_X1 U675 ( .A(n575), .B(n574), .ZN(n704) );
  NOR2_X1 U676 ( .A1(n576), .A2(n704), .ZN(n577) );
  XNOR2_X1 U677 ( .A(n577), .B(KEYINPUT42), .ZN(n754) );
  NAND2_X1 U678 ( .A1(n688), .A2(n578), .ZN(n579) );
  XNOR2_X1 U679 ( .A(KEYINPUT40), .B(n581), .ZN(n753) );
  NOR2_X1 U680 ( .A1(n754), .A2(n753), .ZN(n582) );
  XNOR2_X1 U681 ( .A(n582), .B(KEYINPUT46), .ZN(n583) );
  XNOR2_X1 U682 ( .A(KEYINPUT48), .B(KEYINPUT73), .ZN(n585) );
  NOR2_X1 U683 ( .A1(n667), .A2(n586), .ZN(n669) );
  INV_X1 U684 ( .A(n587), .ZN(n588) );
  NAND2_X1 U685 ( .A1(n588), .A2(n687), .ZN(n589) );
  NOR2_X1 U686 ( .A1(n620), .A2(n589), .ZN(n591) );
  XNOR2_X1 U687 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n590) );
  XNOR2_X1 U688 ( .A(n591), .B(n590), .ZN(n593) );
  NAND2_X1 U689 ( .A1(n593), .A2(n592), .ZN(n670) );
  NAND2_X1 U690 ( .A1(n594), .A2(n670), .ZN(n741) );
  NOR2_X1 U691 ( .A1(G898), .A2(n724), .ZN(n732) );
  NAND2_X1 U692 ( .A1(n595), .A2(n732), .ZN(n596) );
  XOR2_X1 U693 ( .A(KEYINPUT94), .B(n596), .Z(n597) );
  NOR2_X1 U694 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U695 ( .A(KEYINPUT95), .B(n599), .ZN(n601) );
  NAND2_X1 U696 ( .A1(n603), .A2(n671), .ZN(n604) );
  NOR2_X1 U697 ( .A1(n615), .A2(n604), .ZN(n605) );
  XNOR2_X1 U698 ( .A(n605), .B(n474), .ZN(n628) );
  OR2_X1 U699 ( .A1(n620), .A2(n623), .ZN(n606) );
  NOR2_X1 U700 ( .A1(n628), .A2(n606), .ZN(n607) );
  XNOR2_X1 U701 ( .A(KEYINPUT33), .B(KEYINPUT91), .ZN(n609) );
  XNOR2_X1 U702 ( .A(KEYINPUT83), .B(KEYINPUT34), .ZN(n610) );
  INV_X1 U703 ( .A(n610), .ZN(n611) );
  NOR2_X1 U704 ( .A1(n563), .A2(n615), .ZN(n613) );
  NAND2_X1 U705 ( .A1(n614), .A2(n613), .ZN(n649) );
  NOR2_X1 U706 ( .A1(n615), .A2(n681), .ZN(n616) );
  XNOR2_X1 U707 ( .A(KEYINPUT31), .B(n616), .ZN(n666) );
  NAND2_X1 U708 ( .A1(n649), .A2(n666), .ZN(n617) );
  NAND2_X1 U709 ( .A1(n617), .A2(n691), .ZN(n618) );
  OR2_X1 U710 ( .A1(n628), .A2(n620), .ZN(n621) );
  XNOR2_X1 U711 ( .A(n621), .B(KEYINPUT105), .ZN(n622) );
  INV_X1 U712 ( .A(KEYINPUT65), .ZN(n630) );
  INV_X1 U713 ( .A(n624), .ZN(n672) );
  NOR2_X1 U714 ( .A1(n405), .A2(n672), .ZN(n625) );
  NAND2_X1 U715 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U716 ( .A1(n747), .A2(KEYINPUT44), .ZN(n633) );
  INV_X1 U717 ( .A(n634), .ZN(n635) );
  INV_X1 U718 ( .A(KEYINPUT86), .ZN(n636) );
  XNOR2_X1 U719 ( .A(n638), .B(KEYINPUT62), .ZN(n639) );
  XNOR2_X1 U720 ( .A(n640), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U721 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n643) );
  XNOR2_X1 U722 ( .A(n641), .B(KEYINPUT90), .ZN(n642) );
  XOR2_X1 U723 ( .A(G101), .B(n647), .Z(G3) );
  NOR2_X1 U724 ( .A1(n663), .A2(n649), .ZN(n648) );
  XOR2_X1 U725 ( .A(G104), .B(n648), .Z(G6) );
  NOR2_X1 U726 ( .A1(n649), .A2(n667), .ZN(n653) );
  XOR2_X1 U727 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n651) );
  XNOR2_X1 U728 ( .A(G107), .B(KEYINPUT115), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n653), .B(n652), .ZN(G9) );
  XNOR2_X1 U731 ( .A(n654), .B(G110), .ZN(G12) );
  XOR2_X1 U732 ( .A(G128), .B(KEYINPUT29), .Z(n657) );
  INV_X1 U733 ( .A(n667), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n655), .A2(n661), .ZN(n656) );
  XNOR2_X1 U735 ( .A(n657), .B(n656), .ZN(G30) );
  XOR2_X1 U736 ( .A(G143), .B(n658), .Z(n659) );
  XNOR2_X1 U737 ( .A(KEYINPUT116), .B(n659), .ZN(G45) );
  NAND2_X1 U738 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n662), .B(G146), .ZN(G48) );
  NOR2_X1 U740 ( .A1(n663), .A2(n666), .ZN(n665) );
  XNOR2_X1 U741 ( .A(G113), .B(KEYINPUT117), .ZN(n664) );
  XNOR2_X1 U742 ( .A(n665), .B(n664), .ZN(G15) );
  NOR2_X1 U743 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U744 ( .A(G116), .B(n668), .Z(G18) );
  XOR2_X1 U745 ( .A(G134), .B(n669), .Z(G36) );
  XNOR2_X1 U746 ( .A(G140), .B(n670), .ZN(G42) );
  NOR2_X1 U747 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U748 ( .A(KEYINPUT49), .B(n673), .ZN(n678) );
  XNOR2_X1 U749 ( .A(n675), .B(KEYINPUT50), .ZN(n676) );
  XNOR2_X1 U750 ( .A(KEYINPUT120), .B(n676), .ZN(n677) );
  NAND2_X1 U751 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U752 ( .A1(n563), .A2(n679), .ZN(n680) );
  XNOR2_X1 U753 ( .A(n680), .B(KEYINPUT121), .ZN(n682) );
  NAND2_X1 U754 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U755 ( .A(KEYINPUT51), .B(n683), .ZN(n684) );
  NOR2_X1 U756 ( .A1(n704), .A2(n684), .ZN(n685) );
  XNOR2_X1 U757 ( .A(n685), .B(KEYINPUT122), .ZN(n698) );
  NOR2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n695) );
  INV_X1 U760 ( .A(n691), .ZN(n693) );
  NOR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n703), .A2(n696), .ZN(n697) );
  NOR2_X1 U764 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U765 ( .A(n699), .B(KEYINPUT123), .Z(n700) );
  XNOR2_X1 U766 ( .A(KEYINPUT52), .B(n700), .ZN(n701) );
  NOR2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n706) );
  NOR2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U769 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U770 ( .A1(n707), .A2(n395), .ZN(n708) );
  XNOR2_X1 U771 ( .A(KEYINPUT53), .B(KEYINPUT124), .ZN(n709) );
  XNOR2_X1 U772 ( .A(n710), .B(n709), .ZN(G75) );
  XNOR2_X1 U773 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n713) );
  XNOR2_X1 U774 ( .A(n711), .B(KEYINPUT57), .ZN(n712) );
  XNOR2_X1 U775 ( .A(n713), .B(n712), .ZN(n715) );
  XNOR2_X1 U776 ( .A(n718), .B(KEYINPUT126), .ZN(n720) );
  NAND2_X1 U777 ( .A1(G953), .A2(G224), .ZN(n725) );
  XNOR2_X1 U778 ( .A(KEYINPUT61), .B(n725), .ZN(n726) );
  NAND2_X1 U779 ( .A1(n726), .A2(G898), .ZN(n727) );
  NAND2_X1 U780 ( .A1(n728), .A2(n727), .ZN(n734) );
  XNOR2_X1 U781 ( .A(n729), .B(n730), .ZN(n731) );
  NOR2_X1 U782 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U783 ( .A(n734), .B(n733), .ZN(G69) );
  XNOR2_X1 U784 ( .A(n735), .B(n736), .ZN(n740) );
  INV_X1 U785 ( .A(n740), .ZN(n737) );
  XNOR2_X1 U786 ( .A(G227), .B(n737), .ZN(n738) );
  NAND2_X1 U787 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n739), .A2(G953), .ZN(n746) );
  XNOR2_X1 U789 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U790 ( .A(n742), .B(KEYINPUT127), .ZN(n744) );
  NAND2_X1 U791 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U792 ( .A1(n746), .A2(n745), .ZN(G72) );
  XOR2_X1 U793 ( .A(n342), .B(G122), .Z(G24) );
  XOR2_X1 U794 ( .A(KEYINPUT118), .B(KEYINPUT37), .Z(n749) );
  XNOR2_X1 U795 ( .A(G125), .B(KEYINPUT119), .ZN(n748) );
  XNOR2_X1 U796 ( .A(n749), .B(n748), .ZN(n750) );
  XNOR2_X1 U797 ( .A(n751), .B(n750), .ZN(G27) );
  XNOR2_X1 U798 ( .A(G119), .B(n752), .ZN(G21) );
  XOR2_X1 U799 ( .A(G131), .B(n753), .Z(G33) );
  XOR2_X1 U800 ( .A(G137), .B(n754), .Z(G39) );
endmodule

