//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n595,
    new_n596, new_n597, new_n598, new_n600, new_n601, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n645, new_n646, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1236, new_n1237, new_n1238,
    new_n1239;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT65), .B(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT64), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(G137), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n462), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n467), .A2(new_n469), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n464), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n471), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n465), .A2(new_n466), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT66), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n470), .C2(G112), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n465), .A2(new_n478), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n487), .A2(new_n488), .A3(new_n491), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT3), .B(G2104), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n470), .A2(G138), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n467), .A2(new_n469), .A3(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(new_n493), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n493), .A2(new_n495), .B1(new_n497), .B2(new_n465), .ZN(new_n498));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n466), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT67), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n504), .B1(new_n500), .B2(new_n501), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n465), .A2(new_n499), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n511), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n509), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n513), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n521), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  XNOR2_X1  g101(.A(KEYINPUT69), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n514), .A2(new_n518), .A3(G89), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n533));
  AND2_X1   g108(.A1(KEYINPUT5), .A2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n516), .A2(KEYINPUT68), .A3(new_n517), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n536), .A2(new_n537), .A3(G63), .A4(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n512), .A2(G51), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n531), .A2(new_n532), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n529), .A2(new_n530), .B1(G51), .B2(new_n512), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n543), .A2(KEYINPUT70), .A3(new_n538), .A4(new_n532), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n536), .A2(new_n537), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  INV_X1    g125(.A(new_n519), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G90), .B1(G52), .B2(new_n512), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(G171));
  NAND3_X1  g129(.A1(new_n536), .A2(new_n537), .A3(G56), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT71), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  AND3_X1   g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n556), .B1(new_n555), .B2(new_n557), .ZN(new_n559));
  NOR3_X1   g134(.A1(new_n558), .A2(new_n559), .A3(new_n523), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n512), .A2(G43), .ZN(new_n562));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n519), .B2(new_n563), .ZN(new_n564));
  NOR3_X1   g139(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n555), .A2(new_n557), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT71), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n567), .A2(G651), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n564), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT72), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(G153));
  AND3_X1   g148(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G36), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT73), .ZN(G188));
  NAND2_X1  g154(.A1(new_n512), .A2(G53), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT9), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n512), .A2(new_n582), .A3(G53), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT74), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n581), .A2(new_n586), .A3(new_n583), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G78), .A2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n534), .A2(new_n535), .ZN(new_n590));
  INV_X1    g165(.A(G65), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n551), .A2(G91), .B1(new_n592), .B2(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n588), .A2(new_n593), .ZN(G299));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n550), .B2(new_n553), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n549), .A2(G651), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n597), .A2(KEYINPUT75), .A3(new_n552), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n596), .A2(new_n598), .ZN(G301));
  AND3_X1   g174(.A1(new_n542), .A2(KEYINPUT76), .A3(new_n544), .ZN(new_n600));
  AOI21_X1  g175(.A(KEYINPUT76), .B1(new_n542), .B2(new_n544), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(G286));
  INV_X1    g177(.A(G74), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n523), .B1(new_n547), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n512), .A2(G49), .ZN(new_n605));
  INV_X1    g180(.A(G87), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n519), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G288));
  NAND2_X1  g184(.A1(G73), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G61), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n590), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G651), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n612), .A2(KEYINPUT77), .A3(G651), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n512), .A2(G48), .ZN(new_n618));
  INV_X1    g193(.A(G86), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n519), .B2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(G305));
  NAND3_X1  g197(.A1(new_n536), .A2(new_n537), .A3(G60), .ZN(new_n623));
  NAND2_X1  g198(.A1(G72), .A2(G543), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n523), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n512), .A2(G47), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT78), .B(G85), .Z(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n519), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(G290));
  NAND3_X1  g205(.A1(new_n551), .A2(KEYINPUT10), .A3(G92), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT10), .ZN(new_n632));
  INV_X1    g207(.A(G92), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n519), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(G79), .A2(G543), .ZN(new_n636));
  INV_X1    g211(.A(G66), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n590), .B2(new_n637), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n638), .A2(G651), .B1(G54), .B2(new_n512), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  INV_X1    g216(.A(G301), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(G868), .ZN(G284));
  AOI21_X1  g218(.A(new_n641), .B1(new_n642), .B2(G868), .ZN(G321));
  NOR2_X1   g219(.A1(G299), .A2(G868), .ZN(new_n645));
  INV_X1    g220(.A(G286), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(G868), .ZN(G297));
  AOI21_X1  g222(.A(new_n645), .B1(new_n646), .B2(G868), .ZN(G280));
  INV_X1    g223(.A(new_n640), .ZN(new_n649));
  INV_X1    g224(.A(G559), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n649), .B1(new_n650), .B2(G860), .ZN(G148));
  NOR2_X1   g226(.A1(new_n640), .A2(G559), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT79), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G868), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT80), .Z(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(G868), .B2(new_n572), .ZN(G323));
  XNOR2_X1  g231(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g232(.A1(new_n480), .A2(new_n494), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT12), .Z(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT13), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(new_n661));
  OAI221_X1 g236(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n470), .C2(G111), .ZN(new_n662));
  INV_X1    g237(.A(G135), .ZN(new_n663));
  INV_X1    g238(.A(G123), .ZN(new_n664));
  OAI221_X1 g239(.A(new_n662), .B1(new_n484), .B2(new_n663), .C1(new_n664), .C2(new_n489), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(G2096), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n661), .A2(new_n666), .ZN(G156));
  XOR2_X1   g242(.A(KEYINPUT81), .B(KEYINPUT14), .Z(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT15), .B(G2435), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2438), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2427), .B(G2430), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n670), .B2(new_n671), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2451), .B(G2454), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT16), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1341), .B(G1348), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n673), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2443), .B(G2446), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n681), .A3(G14), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT82), .ZN(G401));
  XOR2_X1   g258(.A(G2084), .B(G2090), .Z(new_n684));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(KEYINPUT17), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  AOI21_X1  g263(.A(KEYINPUT18), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2072), .B(G2078), .Z(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n686), .B2(KEYINPUT18), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G2096), .B(G2100), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G227));
  XNOR2_X1  g269(.A(G1956), .B(G2474), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT83), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1961), .B(G1966), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(KEYINPUT84), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(KEYINPUT83), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(KEYINPUT84), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n696), .A2(new_n698), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1971), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT19), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n696), .A2(new_n699), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n698), .A2(new_n700), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n709), .A2(new_n703), .A3(new_n701), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n706), .B(new_n710), .C1(new_n703), .C2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT86), .ZN(new_n712));
  XOR2_X1   g287(.A(G1981), .B(G1986), .Z(new_n713));
  XNOR2_X1  g288(.A(G1991), .B(G1996), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n712), .B(new_n717), .ZN(G229));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G24), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n629), .B2(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(G1986), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G25), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n485), .A2(G131), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n490), .A2(G119), .ZN(new_n727));
  OAI221_X1 g302(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n725), .B1(new_n730), .B2(new_n724), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n719), .A2(G22), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G166), .B2(new_n719), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1971), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n719), .A2(G23), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n608), .B2(new_n719), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT33), .B(G1976), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G6), .A2(G16), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n620), .B1(new_n615), .B2(new_n616), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT32), .B(G1981), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n743), .B(new_n744), .Z(new_n745));
  AND3_X1   g320(.A1(new_n736), .A2(new_n740), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n723), .B(new_n733), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT88), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n747), .A2(new_n749), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT36), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n751), .A2(new_n755), .A3(new_n752), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n572), .A2(new_n719), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n719), .B2(G19), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(G1341), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(G1341), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n719), .A2(G4), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n649), .B2(new_n719), .ZN(new_n764));
  INV_X1    g339(.A(G1348), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n724), .A2(G26), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT28), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n485), .A2(G140), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n490), .A2(G128), .ZN(new_n770));
  OAI221_X1 g345(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n470), .C2(G116), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(new_n724), .ZN(new_n774));
  INV_X1    g349(.A(G2067), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n761), .A2(new_n762), .A3(new_n766), .A4(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n780), .B2(KEYINPUT24), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(KEYINPUT24), .B2(new_n780), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n482), .B2(new_n724), .ZN(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G27), .A2(G29), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G164), .B2(G29), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n785), .B1(new_n787), .B2(G2078), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n783), .A2(new_n784), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G11), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n665), .A2(new_n724), .ZN(new_n793));
  INV_X1    g368(.A(G28), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT30), .ZN(new_n795));
  AOI21_X1  g370(.A(G29), .B1(new_n794), .B2(KEYINPUT30), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n792), .B(new_n793), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n719), .A2(G5), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G171), .B2(new_n719), .ZN(new_n799));
  OAI221_X1 g374(.A(new_n797), .B1(G1961), .B2(new_n799), .C1(G2078), .C2(new_n787), .ZN(new_n800));
  AOI211_X1 g375(.A(new_n790), .B(new_n800), .C1(G1961), .C2(new_n799), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G21), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G168), .B2(G16), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT94), .B(G1966), .Z(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT93), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n719), .A2(G20), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n593), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n585), .B2(new_n587), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n809), .B1(new_n811), .B2(new_n719), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1956), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT91), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n465), .A2(G139), .A3(new_n466), .ZN(new_n816));
  NAND2_X1  g391(.A1(G103), .A2(G2104), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n470), .A2(KEYINPUT25), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(KEYINPUT25), .B1(new_n470), .B2(new_n818), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT90), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT90), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n816), .B(new_n823), .C1(new_n819), .C2(new_n820), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n494), .A2(G127), .ZN(new_n826));
  NAND2_X1  g401(.A1(G115), .A2(G2104), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n470), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n815), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  AOI211_X1 g405(.A(KEYINPUT91), .B(new_n828), .C1(new_n822), .C2(new_n824), .ZN(new_n831));
  OAI21_X1  g406(.A(G29), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G33), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(G29), .B2(new_n833), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n801), .B(new_n814), .C1(G2072), .C2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G2072), .B2(new_n834), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n777), .A2(new_n778), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n724), .A2(G35), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G162), .B2(new_n724), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT29), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G2090), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n724), .A2(G32), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n485), .A2(G141), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT92), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n490), .A2(G129), .ZN(new_n846));
  NAND3_X1  g421(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT26), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n480), .A2(G105), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n842), .B1(new_n851), .B2(new_n724), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT27), .ZN(new_n853));
  INV_X1    g428(.A(G1996), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n841), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n836), .A2(new_n837), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n757), .A2(new_n779), .A3(new_n857), .ZN(G311));
  NAND3_X1  g433(.A1(new_n757), .A2(new_n779), .A3(new_n857), .ZN(G150));
  NAND2_X1  g434(.A1(new_n512), .A2(G55), .ZN(new_n860));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n519), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(G80), .A2(G543), .ZN(new_n863));
  INV_X1    g438(.A(G67), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n547), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n862), .B1(G651), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G860), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT37), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n565), .A2(new_n571), .A3(new_n866), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n523), .B1(new_n566), .B2(KEYINPUT71), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n564), .B1(new_n871), .B2(new_n568), .ZN(new_n872));
  INV_X1    g447(.A(new_n866), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT97), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n866), .B(new_n875), .C1(new_n560), .C2(new_n564), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT98), .B1(new_n870), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n561), .B1(new_n560), .B2(new_n564), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n569), .A2(KEYINPUT72), .A3(new_n570), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n873), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n876), .A4(new_n874), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n640), .A2(new_n650), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT38), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n884), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT99), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n890), .B(new_n867), .C1(new_n888), .C2(new_n887), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n889), .A2(KEYINPUT99), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n869), .B1(new_n891), .B2(new_n892), .ZN(G145));
  XOR2_X1   g468(.A(KEYINPUT102), .B(G37), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n772), .B(new_n507), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n729), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n843), .B(KEYINPUT92), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n898), .A2(new_n846), .A3(new_n848), .A4(new_n849), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n830), .B2(new_n831), .ZN(new_n900));
  INV_X1    g475(.A(new_n830), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n825), .A2(new_n815), .A3(new_n829), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n851), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n465), .A2(G142), .A3(new_n466), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n465), .A2(G130), .A3(new_n478), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n470), .B2(G118), .ZN(new_n907));
  OAI21_X1  g482(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n470), .A2(new_n906), .A3(G118), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n904), .B(new_n905), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n912), .A2(KEYINPUT101), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(KEYINPUT101), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n659), .ZN(new_n916));
  INV_X1    g491(.A(new_n659), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n900), .A2(new_n903), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n919), .B1(new_n900), .B2(new_n903), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n897), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n900), .A2(new_n903), .ZN(new_n923));
  INV_X1    g498(.A(new_n919), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n900), .A2(new_n903), .A3(new_n919), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n896), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n665), .B(G160), .ZN(new_n928));
  XNOR2_X1  g503(.A(G162), .B(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n922), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n922), .B2(new_n927), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n894), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g509(.A(KEYINPUT103), .B(new_n894), .C1(new_n930), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g512(.A(new_n884), .B(new_n653), .ZN(new_n938));
  NAND2_X1  g513(.A1(G299), .A2(new_n649), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n811), .A2(new_n940), .A3(new_n640), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n940), .B1(new_n811), .B2(new_n640), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n942), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT104), .B1(G299), .B2(new_n649), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n946), .A2(KEYINPUT105), .A3(KEYINPUT41), .A4(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n947), .A2(KEYINPUT41), .A3(new_n941), .A4(new_n939), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT41), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n942), .B2(new_n943), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n948), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n945), .B1(new_n938), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(G290), .B(new_n742), .ZN(new_n956));
  XNOR2_X1  g531(.A(G303), .B(new_n608), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT42), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n955), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n955), .A2(new_n961), .ZN(new_n963));
  OAI21_X1  g538(.A(G868), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(G868), .B2(new_n866), .ZN(G295));
  OAI21_X1  g540(.A(new_n964), .B1(G868), .B2(new_n866), .ZN(G331));
  AOI22_X1  g541(.A1(G286), .A2(G171), .B1(G168), .B2(G301), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n878), .A2(new_n883), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n878), .B2(new_n883), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n954), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G171), .ZN(new_n971));
  INV_X1    g546(.A(G168), .ZN(new_n972));
  OAI22_X1  g547(.A1(new_n646), .A2(new_n971), .B1(new_n642), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n877), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n882), .B1(new_n974), .B2(new_n881), .ZN(new_n975));
  AND4_X1   g550(.A1(new_n882), .A2(new_n881), .A3(new_n876), .A4(new_n874), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n944), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n878), .A2(new_n883), .A3(new_n967), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n970), .A2(new_n980), .A3(new_n960), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n981), .A2(new_n894), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n960), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT106), .B1(new_n958), .B2(new_n959), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n968), .A2(new_n969), .A3(new_n944), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n953), .A2(new_n949), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n977), .B2(new_n979), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n982), .A2(new_n983), .A3(new_n984), .A4(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n984), .A3(new_n894), .A4(new_n981), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT107), .ZN(new_n995));
  AOI211_X1 g570(.A(new_n986), .B(new_n987), .C1(new_n970), .C2(new_n980), .ZN(new_n996));
  INV_X1    g571(.A(G37), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n981), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT43), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n993), .A2(new_n995), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(KEYINPUT44), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n982), .A2(KEYINPUT109), .A3(new_n992), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n1003));
  INV_X1    g578(.A(new_n992), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n981), .A2(new_n894), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1006), .A3(KEYINPUT43), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n970), .A2(new_n980), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n988), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(new_n984), .A3(new_n997), .A4(new_n981), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(KEYINPUT108), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(KEYINPUT108), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1007), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1001), .B1(KEYINPUT44), .B2(new_n1013), .ZN(G397));
  NAND4_X1  g589(.A1(new_n471), .A2(new_n479), .A3(G40), .A4(new_n481), .ZN(new_n1015));
  INV_X1    g590(.A(G1384), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n497), .A2(new_n465), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n493), .B1(new_n496), .B2(new_n475), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n503), .A2(new_n505), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(new_n462), .A3(new_n499), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1016), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1015), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT45), .B(new_n1016), .C1(new_n1019), .C2(new_n1023), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n507), .A2(KEYINPUT112), .A3(KEYINPUT45), .A4(new_n1016), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT113), .B(G1971), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1384), .B1(new_n498), .B2(new_n506), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1015), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  OAI22_X1  g613(.A1(new_n1031), .A2(new_n1032), .B1(G2090), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G8), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1040), .A2(KEYINPUT117), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1024), .A2(new_n1015), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1044), .B(new_n1046), .C1(new_n1045), .C2(G288), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G288), .A2(new_n1045), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT52), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(G305), .B2(G1981), .ZN(new_n1054));
  INV_X1    g629(.A(G1981), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n742), .A2(KEYINPUT114), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n742), .B2(new_n1055), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1054), .A2(new_n1056), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1044), .B1(new_n1060), .B2(KEYINPUT49), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1052), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G303), .A2(G8), .ZN(new_n1069));
  XOR2_X1   g644(.A(new_n1069), .B(KEYINPUT55), .Z(new_n1070));
  XNOR2_X1  g645(.A(new_n1040), .B(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1043), .A2(KEYINPUT117), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1041), .B(new_n1068), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n593), .A2(new_n584), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1076));
  INV_X1    g651(.A(G1956), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1038), .A2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT56), .B(G2072), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1076), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1038), .A2(new_n765), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1048), .A2(G2067), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n640), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1078), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1081), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1080), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1015), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1089));
  AOI21_X1  g664(.A(G1956), .B1(new_n1089), .B2(new_n1035), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n811), .A2(new_n1074), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1088), .A2(new_n1090), .B1(new_n1091), .B2(new_n1075), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(KEYINPUT61), .A3(new_n1086), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT119), .B(G1996), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .A4(new_n1094), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT58), .B(G1341), .Z(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1024), .B2(new_n1015), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1048), .A2(KEYINPUT120), .A3(new_n1096), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(new_n1102), .A3(new_n572), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1102), .B1(new_n1101), .B2(new_n572), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1093), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1078), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(new_n1081), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n649), .A2(KEYINPUT60), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n649), .A2(KEYINPUT60), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1082), .A2(new_n1084), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1348), .B1(new_n1089), .B2(new_n1035), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT60), .B(new_n649), .C1(new_n1113), .C2(new_n1083), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1087), .B1(new_n1106), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1118));
  INV_X1    g693(.A(G2078), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1037), .A4(new_n1027), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1026), .A2(KEYINPUT121), .A3(new_n1119), .A4(new_n1027), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(KEYINPUT53), .A3(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .A4(new_n1119), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n1126));
  INV_X1    g701(.A(G1961), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1125), .A2(new_n1126), .B1(new_n1038), .B2(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1124), .A2(new_n1128), .A3(G301), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT110), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT45), .B1(new_n1024), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1015), .A2(new_n1126), .A3(G2078), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1133), .A2(new_n1029), .A3(new_n1030), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n971), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT54), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n642), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1128), .A2(G301), .A3(new_n1135), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1089), .A2(new_n784), .A3(new_n1035), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1145));
  INV_X1    g720(.A(new_n804), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n972), .ZN(new_n1148));
  OAI211_X1 g723(.A(G168), .B(new_n1144), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(new_n1149), .A3(G8), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT51), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT51), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1149), .A2(new_n1152), .A3(G8), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1117), .A2(new_n1143), .A3(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1147), .A2(KEYINPUT63), .A3(G8), .A4(new_n646), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1067), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1071), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1147), .A2(G8), .A3(new_n646), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1073), .B1(new_n1155), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(G288), .A2(G1976), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1049), .B1(new_n1164), .B2(new_n1062), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1039), .A2(G8), .A3(new_n1070), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1067), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT116), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1163), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1049), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1060), .A2(KEYINPUT49), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1062), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1044), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT116), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1039), .A2(G8), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1176), .A2(new_n1177), .A3(new_n1070), .A4(new_n1052), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1174), .A2(new_n1175), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1168), .A2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1181));
  NAND2_X1  g756(.A1(new_n1158), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT122), .B1(new_n1162), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1168), .A2(new_n1179), .B1(new_n1158), .B2(new_n1181), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1159), .B1(new_n1071), .B2(new_n1157), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1101), .A2(new_n572), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1103), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1190), .A2(new_n1109), .A3(new_n1115), .A4(new_n1093), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1191), .A2(new_n1087), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1187), .B1(new_n1192), .B2(new_n1143), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1185), .B(new_n1186), .C1(new_n1193), .C2(new_n1073), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1154), .B(KEYINPUT62), .Z(new_n1195));
  NOR2_X1   g770(.A1(new_n1073), .A2(new_n1139), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1184), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1131), .A2(new_n1037), .A3(new_n1132), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1200), .A2(KEYINPUT111), .A3(new_n854), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT111), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1202), .B1(new_n1199), .B2(G1996), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n899), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1200), .A2(G1996), .A3(new_n899), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n772), .B(G2067), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1200), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n730), .A2(new_n732), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n730), .A2(new_n732), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1199), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  OR3_X1    g786(.A1(new_n1204), .A2(new_n1208), .A3(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n629), .B(new_n722), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1212), .B1(new_n1200), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1198), .A2(new_n1214), .ZN(new_n1215));
  NOR3_X1   g790(.A1(new_n1199), .A2(G1986), .A3(G290), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n1216), .B(KEYINPUT48), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1212), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1200), .B1(new_n899), .B2(new_n1206), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1219), .B(KEYINPUT124), .ZN(new_n1220));
  AND3_X1   g795(.A1(new_n1201), .A2(KEYINPUT46), .A3(new_n1203), .ZN(new_n1221));
  AOI21_X1  g796(.A(KEYINPUT46), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1220), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g798(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1224));
  OR2_X1    g799(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1218), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NOR3_X1   g802(.A1(new_n1204), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1228), .B1(new_n775), .B2(new_n773), .ZN(new_n1229));
  OR3_X1    g804(.A1(new_n1229), .A2(KEYINPUT123), .A3(new_n1199), .ZN(new_n1230));
  OAI21_X1  g805(.A(KEYINPUT123), .B1(new_n1229), .B2(new_n1199), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1227), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n1232), .B(KEYINPUT126), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1215), .A2(new_n1233), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g809(.A1(new_n459), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1236));
  AOI21_X1  g810(.A(new_n1236), .B1(new_n934), .B2(new_n935), .ZN(new_n1237));
  AND3_X1   g811(.A1(new_n1000), .A2(KEYINPUT127), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g812(.A(KEYINPUT127), .B1(new_n1000), .B2(new_n1237), .ZN(new_n1239));
  NOR2_X1   g813(.A1(new_n1238), .A2(new_n1239), .ZN(G308));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n1237), .ZN(G225));
endmodule


