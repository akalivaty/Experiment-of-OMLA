//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g0005(.A(G250), .B1(G257), .B2(G264), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(new_n207), .A2(KEYINPUT0), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n213), .B1(KEYINPUT0), .B2(new_n207), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT65), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n216), .B(new_n217), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AND2_X1   g0025(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n203), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n215), .B1(KEYINPUT1), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(G41), .ZN(new_n246));
  INV_X1    g0046(.A(G45), .ZN(new_n247));
  AOI21_X1  g0047(.A(G1), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n248), .A2(new_n250), .A3(G274), .ZN(new_n251));
  INV_X1    g0051(.A(G226), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n251), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  OAI211_X1 g0059(.A(G222), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  OAI211_X1 g0060(.A(G223), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n250), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n256), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G179), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(G169), .B2(new_n270), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G150), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n209), .A2(G33), .ZN(new_n277));
  NOR3_X1   g0077(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n275), .B1(new_n276), .B2(new_n277), .C1(new_n278), .C2(new_n209), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  AND3_X1   g0080(.A1(new_n280), .A2(KEYINPUT67), .A3(new_n208), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT67), .B1(new_n280), .B2(new_n208), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G1), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G20), .ZN(new_n287));
  INV_X1    g0087(.A(G50), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n253), .B2(G20), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n287), .B(new_n289), .C1(new_n281), .C2(new_n282), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n253), .A2(G13), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(new_n209), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n288), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n290), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n291), .B1(new_n290), .B2(new_n294), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n284), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n273), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n268), .A2(new_n269), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n246), .A2(new_n247), .ZN(new_n301));
  AND2_X1   g0101(.A1(G1), .A2(G13), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n253), .A2(new_n301), .B1(new_n302), .B2(new_n249), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G226), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n300), .A2(new_n251), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT69), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n306), .A3(G200), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT69), .B1(new_n270), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n297), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n284), .B(KEYINPUT9), .C1(new_n295), .C2(new_n296), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n270), .A2(G190), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n310), .A2(new_n312), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT10), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n307), .A2(new_n309), .B1(G190), .B2(new_n270), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(new_n313), .A4(new_n312), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n299), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT70), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G20), .A2(G77), .ZN(new_n322));
  INV_X1    g0122(.A(new_n274), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n322), .B1(new_n276), .B2(new_n323), .C1(new_n277), .C2(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(new_n283), .B1(new_n262), .B2(new_n293), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n283), .A2(new_n293), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n253), .A2(G20), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(G77), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G244), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n251), .B1(new_n331), .B2(new_n255), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n267), .A2(G232), .A3(new_n257), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n267), .A2(G238), .A3(G1698), .ZN(new_n334));
  INV_X1    g0134(.A(G107), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(new_n267), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n332), .B1(new_n336), .B2(new_n269), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n330), .B1(G190), .B2(new_n337), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n337), .A2(new_n308), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n337), .A2(new_n271), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n330), .C1(G169), .C2(new_n337), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n320), .A2(new_n321), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n321), .B1(new_n320), .B2(new_n344), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(KEYINPUT77), .A2(KEYINPUT18), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n276), .B1(new_n253), .B2(G20), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n327), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g0152(.A(KEYINPUT8), .B(G58), .Z(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n287), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n280), .A2(new_n208), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT67), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n280), .A2(KEYINPUT67), .A3(new_n208), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n258), .A2(new_n259), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT7), .B1(new_n360), .B2(new_n209), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n266), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(G68), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G159), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT75), .B1(new_n323), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT75), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n274), .A2(new_n367), .A3(G159), .ZN(new_n368));
  XNOR2_X1  g0168(.A(G58), .B(G68), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n366), .A2(new_n368), .B1(G20), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT16), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n359), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n265), .A2(new_n209), .A3(new_n266), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n376), .A2(KEYINPUT74), .A3(new_n362), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G68), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT16), .B(new_n370), .C1(new_n377), .C2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n354), .B1(new_n373), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G169), .ZN(new_n383));
  INV_X1    g0183(.A(G223), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n257), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n252), .A2(G1698), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n385), .B(new_n386), .C1(new_n258), .C2(new_n259), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G87), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n269), .ZN(new_n390));
  INV_X1    g0190(.A(G274), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n302), .B2(new_n249), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n303), .A2(G232), .B1(new_n392), .B2(new_n248), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n383), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n250), .B1(new_n387), .B2(new_n388), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n250), .A2(G232), .A3(new_n254), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n251), .A2(new_n396), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n395), .A2(new_n397), .A3(new_n271), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT76), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n390), .A2(G179), .A3(new_n393), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT76), .ZN(new_n401));
  OAI21_X1  g0201(.A(G169), .B1(new_n395), .B2(new_n397), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n350), .B1(new_n382), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n366), .A2(new_n368), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n369), .A2(G20), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G68), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n376), .B2(new_n362), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n372), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n381), .A2(new_n283), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n354), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n401), .B1(new_n400), .B2(new_n402), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(KEYINPUT77), .A2(KEYINPUT18), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n350), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n405), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G190), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n390), .A2(new_n422), .A3(new_n393), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n308), .B1(new_n395), .B2(new_n397), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT17), .B1(new_n382), .B2(new_n425), .ZN(new_n426));
  AND4_X1   g0226(.A1(KEYINPUT17), .A2(new_n412), .A3(new_n413), .A4(new_n425), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT73), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n409), .A2(G20), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n431), .B1(new_n277), .B2(new_n262), .C1(new_n323), .C2(new_n288), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n283), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT11), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n293), .A2(new_n409), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT12), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n432), .A2(new_n283), .A3(KEYINPUT11), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n359), .A2(G68), .A3(new_n287), .A4(new_n328), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n435), .A2(new_n437), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT72), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n439), .A2(new_n438), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT72), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(new_n435), .A4(new_n437), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT14), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT13), .ZN(new_n447));
  OAI211_X1 g0247(.A(G232), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT71), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT71), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n267), .A2(new_n450), .A3(G232), .A4(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G97), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n267), .A2(G226), .A3(new_n257), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n449), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n269), .ZN(new_n455));
  INV_X1    g0255(.A(G238), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n251), .B1(new_n456), .B2(new_n255), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n447), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  AOI211_X1 g0259(.A(KEYINPUT13), .B(new_n457), .C1(new_n454), .C2(new_n269), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n446), .B(G169), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n455), .A2(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT13), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n455), .A2(new_n447), .A3(new_n458), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(G179), .A3(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n459), .A2(new_n460), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT14), .B1(new_n467), .B2(new_n383), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n445), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n440), .B1(new_n467), .B2(G190), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n463), .A2(new_n464), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G200), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n430), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n445), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n446), .B1(new_n471), .B2(G169), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n461), .A2(new_n465), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(KEYINPUT73), .A3(new_n473), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n429), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n348), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(G257), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n483));
  OAI211_X1 g0283(.A(G250), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G294), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT82), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT82), .A4(new_n485), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n269), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT5), .B(G41), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n253), .A2(G45), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n491), .A2(new_n493), .B1(new_n302), .B2(new_n249), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G264), .ZN(new_n495));
  OR2_X1    g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  NAND2_X1  g0296(.A1(KEYINPUT5), .A2(G41), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n392), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n490), .A2(G179), .A3(new_n495), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT83), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n250), .B1(new_n486), .B2(new_n487), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(new_n489), .B1(G264), .B2(new_n494), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT83), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(G179), .A4(new_n499), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n490), .A2(new_n495), .A3(new_n499), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G169), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n501), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n209), .B(G87), .C1(new_n258), .C2(new_n259), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT22), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n267), .A2(new_n511), .A3(new_n209), .A4(G87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT24), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G116), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(G20), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT23), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n209), .B2(G107), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n335), .A2(KEYINPUT23), .A3(G20), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n513), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n514), .B1(new_n513), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n283), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n293), .A2(new_n335), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT25), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n253), .A2(G33), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n287), .B(new_n526), .C1(new_n281), .C2(new_n282), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(new_n335), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n508), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n506), .A2(new_n308), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n503), .A2(new_n422), .A3(new_n499), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n525), .A2(new_n528), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n513), .A2(new_n520), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT24), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n513), .A2(new_n514), .A3(new_n520), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n535), .B1(new_n539), .B2(new_n283), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n531), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n323), .A2(new_n262), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n376), .A2(new_n362), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(G107), .ZN(new_n545));
  XNOR2_X1  g0345(.A(G97), .B(G107), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g0347(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT79), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  XOR2_X1   g0350(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n551));
  OAI21_X1  g0351(.A(new_n546), .B1(new_n551), .B2(KEYINPUT79), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n221), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n550), .A2(new_n552), .A3(G20), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n545), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n283), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT80), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n293), .A2(new_n221), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n527), .B2(new_n221), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n359), .B1(new_n545), .B2(new_n554), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT80), .B1(new_n562), .B2(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n491), .A2(new_n493), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(G257), .A3(new_n250), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n499), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(KEYINPUT4), .A2(G244), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n257), .B(new_n568), .C1(new_n258), .C2(new_n259), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G283), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n331), .B1(new_n265), .B2(new_n266), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(KEYINPUT4), .ZN(new_n572));
  OAI21_X1  g0372(.A(G250), .B1(new_n258), .B2(new_n259), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n257), .B1(new_n573), .B2(KEYINPUT4), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n269), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n567), .A2(new_n575), .A3(new_n422), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n220), .B1(new_n265), .B2(new_n266), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT4), .ZN(new_n578));
  OAI21_X1  g0378(.A(G1698), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n360), .B2(new_n331), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n579), .A2(new_n569), .A3(new_n570), .A4(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n566), .B1(new_n581), .B2(new_n269), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n576), .B1(new_n582), .B2(G200), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n561), .A2(new_n563), .A3(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n567), .A2(new_n575), .A3(G179), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n383), .B1(new_n567), .B2(new_n575), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n585), .A2(new_n586), .B1(new_n562), .B2(new_n559), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G116), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n280), .A2(new_n208), .B1(G20), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n570), .B(new_n209), .C1(G33), .C2(new_n221), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT20), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(KEYINPUT20), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n589), .A2(G20), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n594), .A2(new_n595), .B1(new_n286), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n359), .A2(G116), .A3(new_n287), .A4(new_n526), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n494), .A2(G270), .B1(new_n392), .B2(new_n498), .ZN(new_n601));
  OAI211_X1 g0401(.A(G264), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n602));
  OAI211_X1 g0402(.A(G257), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n265), .A2(G303), .A3(new_n266), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n269), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n383), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n600), .A2(new_n607), .A3(KEYINPUT21), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT21), .B1(new_n600), .B2(new_n607), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n594), .A2(new_n595), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n597), .A2(new_n286), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n610), .A2(new_n599), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n601), .A2(new_n606), .A3(G179), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT81), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n601), .A2(new_n606), .A3(G190), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n599), .A3(new_n598), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n308), .B1(new_n601), .B2(new_n606), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n619), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(new_n612), .A3(KEYINPUT81), .A4(new_n617), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n220), .B1(new_n247), .B2(G1), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n253), .A2(new_n391), .A3(G45), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n250), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(G244), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n627));
  OAI211_X1 g0427(.A(G238), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(new_n515), .ZN(new_n629));
  AOI211_X1 g0429(.A(new_n422), .B(new_n626), .C1(new_n629), .C2(new_n269), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n269), .ZN(new_n632));
  INV_X1    g0432(.A(new_n626), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n359), .A2(G87), .A3(new_n287), .A4(new_n526), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT19), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n209), .B1(new_n452), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n219), .A2(new_n221), .A3(new_n335), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n209), .B(G68), .C1(new_n258), .C2(new_n259), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n637), .B1(new_n277), .B2(new_n221), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n283), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n293), .A2(new_n324), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n636), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n631), .A2(new_n635), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n634), .A2(new_n383), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n644), .B(new_n645), .C1(new_n324), .C2(new_n527), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n626), .B1(new_n629), .B2(new_n269), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n271), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n615), .A2(new_n623), .A3(new_n654), .ZN(new_n655));
  NOR4_X1   g0455(.A1(new_n482), .A2(new_n542), .A3(new_n588), .A4(new_n655), .ZN(G372));
  INV_X1    g0456(.A(new_n299), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n316), .A2(new_n319), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n426), .A2(new_n427), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n473), .A2(new_n343), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n479), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT18), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n400), .A2(new_n402), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n414), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n414), .B2(new_n663), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n658), .B1(new_n661), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n636), .A2(new_n644), .A3(new_n645), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n630), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT84), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n634), .B2(G200), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n650), .A2(KEYINPUT84), .A3(new_n308), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(new_n652), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n567), .A2(new_n575), .A3(G179), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n582), .B2(new_n383), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n561), .A2(new_n563), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n675), .A2(new_n676), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n652), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n556), .A2(new_n560), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n682), .A2(new_n678), .A3(new_n647), .A4(new_n652), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n683), .B2(KEYINPUT26), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n541), .A2(new_n584), .A3(new_n587), .A4(new_n674), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n600), .A2(new_n607), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT21), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n600), .A2(new_n607), .A3(KEYINPUT21), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n601), .A2(G179), .A3(new_n606), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n600), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n530), .B2(new_n508), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n680), .B(new_n684), .C1(new_n685), .C2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n657), .B(new_n668), .C1(new_n482), .C2(new_n695), .ZN(G369));
  OR3_X1    g0496(.A1(new_n292), .A2(KEYINPUT27), .A3(G20), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT27), .B1(new_n292), .B2(G20), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n531), .B(new_n541), .C1(new_n540), .C2(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(KEYINPUT83), .A2(new_n500), .B1(new_n506), .B2(G169), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n540), .B1(new_n704), .B2(new_n505), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n701), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n612), .A2(new_n702), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT85), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(new_n615), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n615), .A3(new_n623), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(KEYINPUT86), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT86), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n710), .B2(new_n711), .ZN(new_n715));
  OAI211_X1 g0515(.A(G330), .B(new_n707), .C1(new_n713), .C2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n530), .B1(new_n533), .B2(new_n532), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n705), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n692), .A2(new_n702), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n718), .A2(new_n720), .B1(new_n705), .B2(new_n702), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n716), .A2(new_n721), .ZN(G399));
  NOR2_X1   g0522(.A1(new_n205), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n639), .A2(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n211), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT87), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT29), .B1(new_n694), .B2(new_n702), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n653), .A2(new_n587), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n681), .B1(new_n731), .B2(new_n676), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n557), .B1(new_n556), .B2(new_n560), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n562), .A2(KEYINPUT80), .A3(new_n559), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n678), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n674), .A2(new_n652), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT26), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n732), .B(new_n737), .C1(new_n685), .C2(new_n693), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n738), .A2(new_n702), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n730), .B1(new_n739), .B2(KEYINPUT29), .ZN(new_n740));
  INV_X1    g0540(.A(G330), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n503), .A2(new_n690), .A3(new_n582), .A4(new_n650), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n613), .A2(new_n634), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n745), .A2(KEYINPUT30), .A3(new_n503), .A4(new_n582), .ZN(new_n746));
  INV_X1    g0546(.A(new_n582), .ZN(new_n747));
  AOI21_X1  g0547(.A(G179), .B1(new_n601), .B2(new_n606), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n747), .A2(new_n506), .A3(new_n634), .A4(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n744), .A2(new_n746), .A3(new_n749), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT31), .B1(new_n750), .B2(new_n701), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n655), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n584), .A2(new_n587), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n754), .A2(new_n718), .A3(new_n755), .A4(new_n702), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n741), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n740), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n729), .B1(new_n758), .B2(G1), .ZN(G364));
  OR3_X1    g0559(.A1(new_n713), .A2(G330), .A3(new_n715), .ZN(new_n760));
  OAI21_X1  g0560(.A(G330), .B1(new_n713), .B2(new_n715), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n285), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n253), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n723), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n760), .A2(new_n761), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n267), .A2(new_n204), .ZN(new_n768));
  INV_X1    g0568(.A(G355), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n768), .A2(new_n769), .B1(G116), .B2(new_n204), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n244), .A2(G45), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n205), .A2(new_n267), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n247), .B2(new_n212), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n770), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  OR3_X1    g0575(.A1(KEYINPUT88), .A2(G13), .A3(G33), .ZN(new_n776));
  OAI21_X1  g0576(.A(KEYINPUT88), .B1(G13), .B2(G33), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n209), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n208), .B1(G20), .B2(new_n383), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n765), .B1(new_n775), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(G20), .A2(G190), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n784), .A2(new_n271), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G58), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n209), .A2(G190), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(G179), .A3(new_n308), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n786), .A2(new_n787), .B1(new_n789), .B2(new_n262), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT89), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n209), .A2(new_n271), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n790), .A2(new_n791), .B1(new_n288), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n791), .B2(new_n790), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT90), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n788), .A2(new_n271), .A3(G200), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT91), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT92), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G107), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G179), .A2(G200), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n209), .B1(new_n804), .B2(G190), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G97), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n788), .A2(new_n804), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G159), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(KEYINPUT32), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n792), .A2(new_n422), .A3(G200), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n810), .A2(KEYINPUT32), .B1(new_n813), .B2(G68), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n784), .A2(new_n308), .A3(G179), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n360), .B1(G87), .B2(new_n815), .ZN(new_n816));
  AND4_X1   g0616(.A1(new_n807), .A2(new_n811), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n796), .A2(new_n803), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  INV_X1    g0619(.A(G329), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n789), .A2(new_n819), .B1(new_n808), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G317), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(KEYINPUT33), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(KEYINPUT33), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n813), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G294), .ZN(new_n826));
  INV_X1    g0626(.A(G326), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n805), .C1(new_n827), .C2(new_n793), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n821), .B(new_n828), .C1(G322), .C2(new_n785), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n267), .B1(G303), .B2(new_n815), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT93), .ZN(new_n831));
  INV_X1    g0631(.A(G283), .ZN(new_n832));
  INV_X1    g0632(.A(new_n802), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n829), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n818), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n783), .B1(new_n835), .B2(new_n780), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n712), .B2(new_n779), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n767), .A2(new_n837), .ZN(G396));
  NOR2_X1   g0638(.A1(new_n778), .A2(new_n780), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n766), .B1(new_n262), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n778), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n702), .B1(new_n329), .B2(new_n326), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n342), .B1(new_n340), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n343), .A2(new_n702), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n802), .A2(G68), .ZN(new_n847));
  INV_X1    g0647(.A(new_n815), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n288), .B2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT95), .Z(new_n850));
  AOI21_X1  g0650(.A(new_n360), .B1(new_n809), .B2(G132), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n787), .B2(new_n805), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT96), .ZN(new_n854));
  XOR2_X1   g0654(.A(KEYINPUT94), .B(G143), .Z(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n789), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n785), .A2(new_n856), .B1(new_n857), .B2(G159), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  INV_X1    g0659(.A(G150), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n858), .B1(new_n859), .B2(new_n793), .C1(new_n860), .C2(new_n812), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT34), .Z(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n853), .B2(KEYINPUT96), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n802), .A2(G87), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n809), .A2(G311), .B1(G294), .B2(new_n785), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n335), .B2(new_n848), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n807), .B(new_n360), .C1(new_n589), .C2(new_n789), .ZN(new_n867));
  INV_X1    g0667(.A(G303), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n812), .A2(new_n832), .B1(new_n793), .B2(new_n868), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n854), .A2(new_n863), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n840), .B1(new_n841), .B2(new_n846), .C1(new_n871), .C2(new_n781), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n845), .B1(new_n695), .B2(new_n701), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n846), .A2(new_n694), .A3(new_n702), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n757), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n765), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n876), .B2(new_n875), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n872), .A2(new_n878), .ZN(G384));
  NAND2_X1  g0679(.A1(new_n753), .A2(new_n756), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n441), .A2(new_n444), .A3(new_n701), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT97), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n469), .B2(new_n474), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT97), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n881), .B(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n479), .A2(new_n885), .A3(new_n473), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n845), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n412), .A2(new_n413), .A3(new_n425), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n382), .B2(new_n699), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n382), .B2(new_n404), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT98), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT37), .B1(new_n414), .B2(new_n417), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT98), .ZN(new_n894));
  INV_X1    g0694(.A(new_n699), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n414), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n893), .A2(new_n894), .A3(new_n888), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n381), .A2(new_n283), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT74), .ZN(new_n900));
  OAI211_X1 g0700(.A(G68), .B(new_n379), .C1(new_n544), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT16), .B1(new_n901), .B2(new_n370), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n413), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n895), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n663), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(new_n888), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT37), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n898), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n903), .A2(new_n895), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n429), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n892), .A2(new_n897), .B1(new_n906), .B2(KEYINPUT37), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n904), .B1(new_n421), .B2(new_n428), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n880), .B(new_n887), .C1(new_n911), .C2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n414), .A2(new_n663), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n896), .A3(new_n888), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n892), .A2(new_n897), .B1(KEYINPUT37), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n896), .B1(new_n666), .B2(new_n428), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n914), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n917), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n883), .A2(new_n886), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n925), .A2(new_n880), .A3(new_n846), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n916), .A2(new_n917), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n429), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n479), .A2(KEYINPUT73), .A3(new_n473), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT73), .B1(new_n479), .B2(new_n473), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n658), .A2(new_n657), .A3(new_n344), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT70), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n345), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n880), .ZN(new_n937));
  OAI21_X1  g0737(.A(G330), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n928), .B2(new_n937), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n918), .A2(new_n923), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n469), .A2(new_n702), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n914), .B1(new_n912), .B2(new_n913), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n918), .A2(new_n945), .A3(KEYINPUT39), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n874), .A2(new_n844), .B1(new_n886), .B2(new_n883), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n918), .A2(new_n945), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n948), .A2(new_n949), .B1(new_n667), .B2(new_n699), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n668), .A2(new_n657), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n740), .B2(new_n936), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n939), .A2(new_n954), .B1(new_n253), .B2(new_n762), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n939), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT35), .ZN(new_n958));
  OAI211_X1 g0758(.A(G116), .B(new_n210), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n958), .B2(new_n957), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT36), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n212), .B(G77), .C1(new_n787), .C2(new_n409), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n288), .A2(G68), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n253), .B(G13), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n956), .A2(new_n961), .A3(new_n964), .ZN(G367));
  XOR2_X1   g0765(.A(new_n723), .B(KEYINPUT41), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n679), .A2(new_n701), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n755), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n679), .A2(new_n678), .A3(new_n701), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n721), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n721), .A2(new_n970), .A3(KEYINPUT45), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT101), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n976), .B(KEYINPUT44), .C1(new_n721), .C2(new_n970), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(KEYINPUT44), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n970), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n721), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n976), .A2(KEYINPUT44), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n975), .A2(new_n977), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n716), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  MUX2_X1   g0785(.A(new_n542), .B(new_n707), .S(new_n719), .Z(new_n986));
  XNOR2_X1  g0786(.A(new_n761), .B(new_n986), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n975), .A2(new_n716), .A3(new_n977), .A4(new_n982), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n985), .A2(new_n987), .A3(new_n758), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n966), .B1(new_n989), .B2(new_n758), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n764), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n646), .A2(new_n702), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n681), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n736), .B2(new_n993), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT43), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT100), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n970), .A2(new_n705), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n701), .B1(new_n998), .B2(new_n587), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT42), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n588), .A2(new_n719), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(new_n707), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT99), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1002), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n531), .B1(new_n968), .B2(new_n969), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n587), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n702), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT99), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n707), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n997), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1011), .ZN(new_n1013));
  AOI211_X1 g0813(.A(KEYINPUT100), .B(new_n1013), .C1(new_n1003), .C2(new_n1009), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n996), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1009), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1008), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1011), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT100), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1010), .A2(new_n997), .A3(new_n1011), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1015), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n984), .A2(new_n970), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1015), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n992), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n805), .A2(new_n335), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n815), .A2(G116), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT46), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1029), .B(new_n1032), .C1(G294), .C2(new_n813), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n789), .A2(new_n832), .B1(new_n808), .B2(new_n822), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n267), .B(new_n1034), .C1(G303), .C2(new_n785), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n801), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(G97), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n793), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1038), .A2(G311), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1033), .A2(new_n1035), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n267), .B1(new_n801), .B2(new_n262), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n805), .A2(new_n409), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G150), .B2(new_n785), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n793), .B2(new_n855), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(KEYINPUT103), .A2(new_n1041), .B1(new_n1044), .B2(KEYINPUT102), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(KEYINPUT102), .B2(new_n1044), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n808), .A2(new_n859), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n848), .A2(new_n787), .B1(new_n789), .B2(new_n288), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G159), .C2(new_n813), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(KEYINPUT103), .B2(new_n1041), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1040), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT47), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n780), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n995), .A2(new_n779), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n324), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n782), .B1(new_n205), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n236), .A2(new_n772), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n766), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1053), .A2(new_n1054), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1028), .A2(new_n1059), .ZN(G387));
  NAND2_X1  g0860(.A1(new_n987), .A2(new_n764), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT104), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n768), .A2(new_n725), .B1(G107), .B2(new_n204), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n233), .A2(new_n247), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n725), .ZN(new_n1066));
  AOI211_X1 g0866(.A(G45), .B(new_n1066), .C1(G68), .C2(G77), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n276), .A2(G50), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT50), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n773), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1064), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n848), .A2(new_n826), .B1(new_n805), .B2(new_n832), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n857), .A2(G303), .B1(new_n785), .B2(G317), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1038), .A2(G322), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(new_n819), .C2(new_n812), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT48), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n1076), .B2(new_n1075), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT49), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n360), .B1(new_n808), .B2(new_n827), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n1036), .B2(G116), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n802), .A2(G97), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n806), .A2(new_n1055), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1083), .B(new_n267), .C1(new_n860), .C2(new_n808), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G50), .A2(new_n785), .B1(new_n815), .B2(G77), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n409), .B2(new_n789), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n365), .A2(new_n793), .B1(new_n812), .B2(new_n276), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1079), .A2(new_n1081), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n765), .B1(new_n782), .B2(new_n1071), .C1(new_n1089), .C2(new_n781), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT105), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n707), .B2(new_n779), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1063), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n987), .A2(new_n758), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n987), .A2(new_n758), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n723), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1094), .A2(new_n1097), .ZN(G393));
  INV_X1    g0898(.A(new_n988), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n982), .A2(new_n977), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n716), .B1(new_n1100), .B2(new_n975), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1096), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n723), .A3(new_n989), .ZN(new_n1103));
  OAI21_X1  g0903(.A(KEYINPUT106), .B1(new_n1101), .B2(new_n1099), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT106), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n985), .A2(new_n1105), .A3(new_n988), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n764), .A3(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n970), .A2(new_n779), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1109), .A2(KEYINPUT107), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(KEYINPUT107), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n786), .A2(new_n819), .B1(new_n793), .B2(new_n822), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT52), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n360), .B1(new_n789), .B2(new_n826), .C1(new_n812), .C2(new_n868), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G116), .B2(new_n806), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n809), .A2(G322), .B1(G283), .B2(new_n815), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT108), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n803), .A2(new_n1113), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n786), .A2(new_n365), .B1(new_n793), .B2(new_n860), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT51), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n848), .A2(new_n409), .B1(new_n789), .B2(new_n276), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n812), .A2(new_n288), .B1(new_n805), .B2(new_n262), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n267), .B1(new_n855), .B2(new_n808), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n864), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n781), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n241), .A2(new_n773), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n782), .B1(G97), .B2(new_n205), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n766), .B(new_n1126), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT109), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1110), .A2(new_n1111), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1103), .A2(new_n1107), .A3(new_n1131), .ZN(G390));
  INV_X1    g0932(.A(new_n946), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT39), .B1(new_n918), .B2(new_n923), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1133), .A2(new_n1134), .B1(new_n948), .B2(new_n944), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n738), .A2(new_n702), .A3(new_n843), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n844), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n925), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n944), .B1(new_n918), .B2(new_n923), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1138), .A2(new_n1139), .A3(KEYINPUT110), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT110), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1135), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n757), .A2(new_n887), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NOR4_X1   g0945(.A1(new_n542), .A2(new_n655), .A3(new_n588), .A4(new_n701), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n750), .A2(new_n701), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT31), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(G330), .B(new_n846), .C1(new_n1146), .C2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n925), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1137), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1154), .A2(new_n1155), .A3(new_n1143), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n874), .A2(new_n844), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1154), .B2(new_n1143), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT111), .B1(new_n936), .B2(new_n757), .ZN(new_n1160));
  AND4_X1   g0960(.A1(KEYINPUT111), .A2(new_n348), .A3(new_n481), .A4(new_n757), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n953), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1135), .B(new_n1143), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1145), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(KEYINPUT112), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT112), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1145), .A2(new_n1164), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n723), .B(new_n1165), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n267), .B1(new_n801), .B2(new_n288), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1172), .A2(KEYINPUT113), .B1(G125), .B2(new_n809), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(KEYINPUT113), .B2(new_n1172), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT114), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n785), .A2(G132), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT54), .B(G143), .ZN(new_n1177));
  XOR2_X1   g0977(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n815), .A2(G150), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1176), .B1(new_n789), .B2(new_n1177), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G137), .A2(new_n813), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1182));
  INV_X1    g0982(.A(G128), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1182), .B1(new_n1183), .B2(new_n793), .C1(new_n365), .C2(new_n805), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1175), .A2(new_n1181), .A3(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n809), .A2(G294), .B1(G116), .B2(new_n785), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n221), .B2(new_n789), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n360), .B1(new_n805), .B2(new_n262), .C1(new_n848), .C2(new_n219), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n812), .A2(new_n335), .B1(new_n793), .B2(new_n832), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n847), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n780), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n839), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(new_n765), .C1(new_n353), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n942), .A2(new_n946), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n778), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1170), .B2(new_n764), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1171), .A2(new_n1197), .ZN(G378));
  INV_X1    g0998(.A(KEYINPUT57), .ZN(new_n1199));
  XOR2_X1   g0999(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT117), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n298), .A2(new_n699), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n320), .A2(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n299), .B(new_n1203), .C1(new_n316), .C2(new_n319), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1202), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n320), .A2(new_n1204), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1209), .A2(new_n1206), .A3(KEYINPUT117), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1201), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1205), .A2(new_n1207), .A3(new_n1202), .ZN(new_n1212));
  OAI21_X1  g1012(.A(KEYINPUT117), .B1(new_n1209), .B2(new_n1206), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n1200), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n911), .A2(new_n915), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n887), .A2(new_n880), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n917), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n924), .A2(new_n926), .ZN(new_n1219));
  AND4_X1   g1019(.A1(G330), .A2(new_n1215), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1215), .B1(new_n927), .B2(G330), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n951), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1218), .A2(G330), .A3(new_n1219), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1215), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n951), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n927), .A2(G330), .A3(new_n1215), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1199), .B1(new_n1222), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1162), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1165), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1165), .A2(new_n1230), .B1(new_n1222), .B2(new_n1228), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n723), .C1(KEYINPUT57), .C2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n763), .B1(new_n1222), .B2(new_n1228), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1224), .A2(new_n778), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1036), .A2(G58), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n360), .A2(new_n246), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1238), .B(new_n1042), .C1(G77), .C2(new_n815), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n813), .A2(G97), .B1(new_n1038), .B2(G116), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n789), .A2(new_n324), .B1(new_n808), .B2(new_n832), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G107), .B2(new_n785), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1237), .A2(new_n1239), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT58), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G50), .B1(new_n264), .B2(new_n246), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1243), .A2(new_n1244), .B1(new_n1238), .B2(new_n1245), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n786), .A2(new_n1183), .B1(new_n789), .B2(new_n859), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n848), .A2(new_n1177), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(KEYINPUT116), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G150), .B2(new_n806), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n813), .A2(G132), .B1(new_n1038), .B2(G125), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1247), .B(new_n1252), .C1(KEYINPUT116), .C2(new_n1248), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT59), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1036), .A2(G159), .ZN(new_n1256));
  AOI211_X1 g1056(.A(G33), .B(G41), .C1(new_n809), .C2(G124), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1254), .A2(KEYINPUT59), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1246), .B1(new_n1244), .B2(new_n1243), .C1(new_n1258), .C2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n780), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n839), .A2(new_n288), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1236), .A2(new_n765), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT118), .B1(new_n1235), .B2(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1226), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n764), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT118), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1263), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1265), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1234), .A2(new_n1271), .ZN(G375));
  AND2_X1   g1072(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1273));
  OR3_X1    g1073(.A1(new_n1169), .A2(new_n966), .A3(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n765), .B1(new_n1193), .B2(G68), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n786), .A2(new_n859), .B1(new_n789), .B2(new_n860), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(G159), .B2(new_n815), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n267), .B1(new_n808), .B2(new_n1183), .C1(new_n812), .C2(new_n1177), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1038), .A2(G132), .B1(new_n806), .B2(G50), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1237), .A2(new_n1277), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n833), .A2(new_n262), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n786), .A2(new_n832), .B1(new_n808), .B2(new_n868), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(G97), .B2(new_n815), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n813), .A2(G116), .B1(new_n1038), .B2(G294), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n267), .B1(new_n857), .B2(G107), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1083), .A4(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1281), .B1(new_n1282), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1275), .B1(new_n1288), .B2(new_n780), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(new_n925), .B2(new_n841), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1159), .A2(new_n763), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1291), .B2(KEYINPUT119), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(KEYINPUT119), .B2(new_n1291), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1274), .A2(new_n1293), .ZN(G381));
  XOR2_X1   g1094(.A(G375), .B(KEYINPUT120), .Z(new_n1295));
  INV_X1    g1095(.A(G390), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1027), .B1(new_n764), .B2(new_n990), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1024), .B1(new_n1015), .B2(new_n1022), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1059), .B(new_n1296), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1097), .ZN(new_n1300));
  OR3_X1    g1100(.A1(new_n1093), .A2(G396), .A3(new_n1300), .ZN(new_n1301));
  OR3_X1    g1101(.A1(G381), .A2(G384), .A3(new_n1301), .ZN(new_n1302));
  OR4_X1    g1102(.A1(G378), .A2(new_n1295), .A3(new_n1299), .A4(new_n1302), .ZN(G407));
  INV_X1    g1103(.A(G378), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n700), .A2(G213), .ZN(new_n1305));
  XOR2_X1   g1105(.A(new_n1305), .B(KEYINPUT121), .Z(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G407), .B(G213), .C1(new_n1295), .C2(new_n1307), .ZN(G409));
  INV_X1    g1108(.A(new_n1163), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1273), .B1(new_n1309), .B2(KEYINPUT60), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1159), .A2(new_n1162), .A3(KEYINPUT60), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n723), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1293), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(G384), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1293), .B(G384), .C1(new_n1310), .C2(new_n1312), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1317), .A2(G213), .A3(new_n700), .A4(G2897), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1306), .ZN(new_n1319));
  INV_X1    g1119(.A(G2897), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1318), .B1(new_n1317), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1233), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1268), .B(new_n1263), .C1(new_n1323), .C2(new_n966), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1304), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1234), .A2(new_n1271), .A3(G378), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1305), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1322), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1327), .A2(new_n1305), .A3(new_n1317), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1327), .A2(new_n1319), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1317), .ZN(new_n1335));
  OAI21_X1  g1135(.A(G396), .B1(new_n1093), .B2(new_n1300), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1301), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT122), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1299), .A2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1296), .B1(new_n1028), .B2(new_n1059), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1338), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1027), .ZN(new_n1343));
  NOR3_X1   g1143(.A1(new_n1343), .A2(new_n991), .A3(new_n1298), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1059), .ZN(new_n1345));
  OAI21_X1  g1145(.A(G390), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1346), .A2(new_n1339), .A3(new_n1299), .A4(new_n1337), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1342), .A2(new_n1347), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1348), .A2(KEYINPUT61), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1329), .A2(new_n1332), .A3(new_n1335), .A4(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1334), .A2(KEYINPUT62), .A3(new_n1317), .ZN(new_n1351));
  XOR2_X1   g1151(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n1352));
  NAND2_X1  g1152(.A1(new_n1330), .A2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1351), .A2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(KEYINPUT61), .B1(new_n1322), .B2(new_n1333), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1348), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1350), .B1(new_n1356), .B2(new_n1357), .ZN(G405));
  INV_X1    g1158(.A(KEYINPUT126), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1234), .A2(new_n1271), .A3(G378), .ZN(new_n1360));
  AOI21_X1  g1160(.A(G378), .B1(new_n1234), .B2(new_n1271), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1317), .B1(new_n1360), .B2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(G375), .A2(new_n1304), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1363), .A2(new_n1364), .A3(new_n1326), .ZN(new_n1365));
  AOI211_X1 g1165(.A(KEYINPUT125), .B(new_n1348), .C1(new_n1362), .C2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT125), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1362), .A2(new_n1365), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1367), .B1(new_n1368), .B2(new_n1357), .ZN(new_n1369));
  NOR2_X1   g1169(.A1(new_n1366), .A2(new_n1369), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1362), .A2(new_n1365), .A3(new_n1348), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT124), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1373));
  NAND4_X1  g1173(.A1(new_n1362), .A2(new_n1365), .A3(new_n1348), .A4(KEYINPUT124), .ZN(new_n1374));
  AND2_X1   g1174(.A1(new_n1373), .A2(new_n1374), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1359), .B1(new_n1370), .B2(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1373), .A2(new_n1374), .ZN(new_n1377));
  OAI211_X1 g1177(.A(new_n1377), .B(KEYINPUT126), .C1(new_n1369), .C2(new_n1366), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1376), .A2(new_n1378), .ZN(G402));
endmodule


