//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n588, new_n591, new_n592, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n637,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT64), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  XOR2_X1   g032(.A(G325), .B(KEYINPUT65), .Z(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(KEYINPUT66), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(KEYINPUT66), .B2(new_n460), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND3_X1   g038(.A1(KEYINPUT67), .A2(G113), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT67), .B1(G113), .B2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n463), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n463), .C1(new_n467), .C2(new_n468), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n463), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT68), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(G124), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n480), .A2(new_n485), .ZN(G162));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n467), .B2(new_n468), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(KEYINPUT69), .A3(new_n488), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(KEYINPUT4), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n489), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n498));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n494), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  OR2_X1    g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT70), .ZN(new_n507));
  AOI21_X1  g082(.A(KEYINPUT70), .B1(new_n505), .B2(new_n506), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G88), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n505), .A2(G62), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(KEYINPUT71), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n505), .A2(new_n520), .A3(G62), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n517), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n510), .B(new_n516), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n518), .A2(KEYINPUT71), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n521), .ZN(new_n528));
  OAI21_X1  g103(.A(G651), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(KEYINPUT72), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n524), .A2(new_n530), .ZN(G166));
  AND2_X1   g106(.A1(new_n505), .A2(G63), .ZN(new_n532));
  AND3_X1   g107(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n533));
  OAI21_X1  g108(.A(G651), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT73), .B(G51), .Z(new_n535));
  INV_X1    g110(.A(KEYINPUT7), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n515), .A2(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n509), .A2(G89), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(new_n509), .A2(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AND2_X1   g118(.A1(KEYINPUT5), .A2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(KEYINPUT5), .A2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G651), .B1(new_n515), .B2(G52), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n517), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n553), .A2(new_n554), .B1(G43), .B2(new_n515), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT74), .B1(new_n552), .B2(new_n517), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n509), .A2(G81), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n555), .A2(KEYINPUT75), .A3(new_n556), .A4(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g140(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n566));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(new_n515), .A2(G53), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT77), .B1(new_n507), .B2(new_n508), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n573), .B1(new_n546), .B2(new_n513), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT70), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n572), .A2(G91), .A3(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(new_n517), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n571), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT78), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G299));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n550), .B(new_n588), .ZN(G301));
  INV_X1    g164(.A(G168), .ZN(G286));
  NAND2_X1  g165(.A1(new_n529), .A2(KEYINPUT72), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n522), .A2(new_n523), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n591), .A2(new_n592), .A3(new_n510), .A4(new_n516), .ZN(G303));
  NAND3_X1  g168(.A1(new_n572), .A2(G87), .A3(new_n577), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n505), .A2(G74), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(new_n515), .B2(G49), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(G288));
  NAND2_X1  g172(.A1(new_n515), .A2(G48), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(G61), .B1(new_n544), .B2(new_n545), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g179(.A(KEYINPUT80), .B(G61), .C1(new_n544), .C2(new_n545), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n517), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(KEYINPUT81), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n572), .A2(G86), .A3(new_n577), .ZN(new_n608));
  INV_X1    g183(.A(G61), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n503), .B2(new_n504), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n600), .B1(new_n610), .B2(KEYINPUT80), .ZN(new_n611));
  INV_X1    g186(.A(new_n605), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT81), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n607), .A2(new_n608), .A3(new_n615), .ZN(G305));
  XNOR2_X1  g191(.A(KEYINPUT82), .B(G85), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n509), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(G72), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G60), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n546), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n621), .A2(G651), .B1(new_n515), .B2(G47), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(G290));
  INV_X1    g198(.A(new_n515), .ZN(new_n624));
  INV_X1    g199(.A(G54), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n626));
  OAI22_X1  g201(.A1(new_n624), .A2(new_n625), .B1(new_n626), .B2(new_n517), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n572), .A2(G92), .A3(new_n577), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n572), .A2(KEYINPUT10), .A3(G92), .A4(new_n577), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  MUX2_X1   g208(.A(new_n633), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g209(.A(new_n633), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g210(.A1(G286), .A2(G868), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT83), .Z(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n586), .ZN(G297));
  OAI21_X1  g213(.A(new_n637), .B1(G868), .B2(new_n586), .ZN(G280));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n632), .B1(new_n640), .B2(G860), .ZN(G148));
  OAI21_X1  g216(.A(KEYINPUT84), .B1(new_n563), .B2(G868), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n633), .A2(G559), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G868), .ZN(new_n645));
  MUX2_X1   g220(.A(KEYINPUT84), .B(new_n642), .S(new_n645), .Z(G323));
  XNOR2_X1  g221(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g222(.A1(new_n492), .A2(new_n472), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n651), .A2(G2100), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT85), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n478), .A2(G135), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n484), .A2(G123), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n463), .A2(G111), .ZN(new_n656));
  OAI21_X1  g231(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n654), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2096), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n651), .B2(G2100), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n653), .A2(new_n660), .ZN(G156));
  INV_X1    g236(.A(KEYINPUT14), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2427), .B(G2438), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2430), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2451), .B(G2454), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1341), .B(G1348), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n667), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2443), .B(G2446), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  AND3_X1   g250(.A1(new_n674), .A2(G14), .A3(new_n675), .ZN(G401));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  XNOR2_X1  g252(.A(G2067), .B(G2678), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  NOR2_X1   g254(.A1(G2072), .A2(G2078), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n444), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n677), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(KEYINPUT17), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n679), .B2(new_n683), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n677), .B(new_n678), .C1(new_n444), .C2(new_n680), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT18), .Z(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n679), .A3(new_n677), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2096), .B(G2100), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1956), .B(G2474), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT87), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1961), .B(G1966), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n695), .A2(new_n697), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n693), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n701), .A2(new_n698), .A3(new_n693), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n699), .B1(new_n698), .B2(new_n693), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(G1981), .B(G1986), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(G229));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G35), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G162), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(KEYINPUT29), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n717), .B(new_n714), .C1(G162), .C2(new_n713), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G2090), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT103), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT26), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n484), .A2(G129), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n478), .A2(G141), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n472), .A2(G105), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(new_n713), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n713), .B2(G32), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT27), .B(G1996), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G2084), .ZN(new_n734));
  INV_X1    g309(.A(G34), .ZN(new_n735));
  AOI21_X1  g310(.A(G29), .B1(new_n735), .B2(KEYINPUT24), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(KEYINPUT24), .B2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(G160), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n713), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n733), .B1(new_n734), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G16), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G5), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G171), .B2(new_n741), .ZN(new_n743));
  INV_X1    g318(.A(G1961), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n713), .A2(G33), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n492), .A2(G127), .ZN(new_n747));
  NAND2_X1  g322(.A1(G115), .A2(G2104), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n463), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n478), .A2(G139), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT25), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n749), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n746), .B1(new_n754), .B2(new_n713), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(new_n442), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n739), .A2(new_n734), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n731), .A2(new_n732), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n756), .A2(KEYINPUT100), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT30), .B(G28), .ZN(new_n760));
  OR2_X1    g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  NAND2_X1  g336(.A1(KEYINPUT31), .A2(G11), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n760), .A2(new_n713), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n658), .B2(new_n713), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT102), .Z(new_n765));
  NAND4_X1  g340(.A1(new_n740), .A2(new_n745), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  AND3_X1   g341(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n767));
  OAI22_X1  g342(.A1(new_n767), .A2(KEYINPUT100), .B1(new_n719), .B2(G2090), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n721), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(G168), .A2(G16), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n770), .B(KEYINPUT101), .C1(G16), .C2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(KEYINPUT101), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G1966), .ZN(new_n773));
  NOR2_X1   g348(.A1(G27), .A2(G29), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G164), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(new_n443), .ZN(new_n776));
  INV_X1    g351(.A(G1966), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n771), .B(new_n777), .C1(KEYINPUT101), .C2(new_n770), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n773), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT91), .B(G16), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G19), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n563), .B2(new_n780), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT94), .B(G1341), .Z(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n782), .A2(new_n784), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n779), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n780), .A2(G20), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT23), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n586), .B2(new_n741), .ZN(new_n790));
  INV_X1    g365(.A(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n632), .A2(G16), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G4), .B2(G16), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT93), .B(G1348), .Z(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n794), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n478), .A2(G140), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT95), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n484), .A2(G128), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT96), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n463), .A2(G116), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n800), .B(new_n802), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G29), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT97), .B(KEYINPUT28), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT98), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n713), .A2(G26), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n808), .B(new_n809), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT99), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(KEYINPUT99), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G2067), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n812), .A2(G2067), .A3(new_n813), .ZN(new_n817));
  AOI211_X1 g392(.A(new_n797), .B(new_n798), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n769), .A2(new_n787), .A3(new_n792), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G6), .A2(G16), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n607), .A2(new_n608), .A3(new_n615), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(G16), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT32), .B(G1981), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(G1971), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n780), .A2(G22), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G166), .B2(new_n780), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n824), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(G1971), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n741), .A2(G23), .ZN(new_n832));
  INV_X1    g407(.A(G288), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n741), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT33), .B(G1976), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n822), .A2(new_n823), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OR3_X1    g413(.A1(new_n831), .A2(KEYINPUT34), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n713), .A2(G25), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n478), .A2(G131), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT89), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n484), .A2(G119), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n463), .A2(G107), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT90), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n840), .B1(new_n847), .B2(new_n713), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G1991), .Z(new_n849));
  XOR2_X1   g424(.A(new_n848), .B(new_n849), .Z(new_n850));
  INV_X1    g425(.A(new_n780), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(G24), .ZN(new_n852));
  INV_X1    g427(.A(G290), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(new_n851), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT92), .B(G1986), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT34), .B1(new_n831), .B2(new_n838), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n839), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT36), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT36), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n839), .A2(new_n857), .A3(new_n861), .A4(new_n858), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n819), .B1(new_n860), .B2(new_n862), .ZN(G311));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n862), .ZN(new_n864));
  INV_X1    g439(.A(new_n819), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT104), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n867));
  AOI211_X1 g442(.A(new_n867), .B(new_n819), .C1(new_n860), .C2(new_n862), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n866), .A2(new_n868), .ZN(G150));
  AOI22_X1  g444(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(new_n517), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT105), .B(G55), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n515), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n574), .A2(new_n576), .ZN(new_n874));
  INV_X1    g449(.A(G93), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n871), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(new_n560), .B2(new_n561), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n558), .A2(new_n876), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT38), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n633), .A2(new_n640), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n884));
  AOI21_X1  g459(.A(G860), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n884), .B2(new_n883), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n876), .A2(G860), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(KEYINPUT37), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(G145));
  XOR2_X1   g464(.A(KEYINPUT107), .B(G37), .Z(new_n890));
  OR2_X1    g465(.A1(new_n805), .A2(new_n501), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n805), .A2(new_n501), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n728), .B2(new_n725), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n754), .A2(KEYINPUT106), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n729), .A3(new_n892), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(KEYINPUT106), .A3(new_n754), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n754), .A2(KEYINPUT106), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n894), .A2(new_n899), .A3(new_n895), .A4(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n846), .B(new_n649), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n478), .A2(G142), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n484), .A2(G130), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n463), .A2(G118), .ZN(new_n905));
  OAI21_X1  g480(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n903), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n902), .B(new_n907), .Z(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n901), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n658), .B(G160), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(G162), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n898), .A2(new_n908), .A3(new_n900), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n910), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n910), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n890), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT42), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n920), .A2(KEYINPUT42), .ZN(new_n922));
  NAND2_X1  g497(.A1(G166), .A2(G305), .ZN(new_n923));
  NAND2_X1  g498(.A1(G303), .A2(new_n821), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n833), .A2(G290), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n853), .A2(G288), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n923), .A2(new_n924), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n923), .A2(new_n924), .B1(new_n926), .B2(new_n925), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n921), .B(new_n922), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n923), .A2(new_n924), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n925), .A2(new_n926), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(new_n927), .A3(new_n920), .A4(KEYINPUT42), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n919), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n632), .B1(new_n583), .B2(new_n585), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n583), .A2(new_n585), .A3(new_n632), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n644), .A2(new_n880), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n643), .B1(new_n878), .B2(new_n879), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT41), .ZN(new_n944));
  INV_X1    g519(.A(new_n938), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(new_n936), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n937), .A2(KEYINPUT41), .A3(new_n938), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n946), .A2(new_n947), .B1(new_n940), .B2(new_n941), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n935), .B1(new_n943), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n930), .A2(new_n919), .A3(new_n934), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n935), .A2(new_n948), .A3(new_n943), .ZN(new_n952));
  OAI21_X1  g527(.A(G868), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n877), .A2(G868), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(G295));
  NOR2_X1   g531(.A1(new_n948), .A2(new_n943), .ZN(new_n957));
  INV_X1    g532(.A(new_n935), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(new_n950), .A3(new_n949), .ZN(new_n960));
  AOI211_X1 g535(.A(KEYINPUT110), .B(new_n954), .C1(new_n960), .C2(G868), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n953), .B2(new_n955), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(G331));
  NAND2_X1  g539(.A1(new_n946), .A2(new_n947), .ZN(new_n965));
  NAND2_X1  g540(.A1(G286), .A2(new_n550), .ZN(new_n966));
  OAI221_X1 g541(.A(new_n966), .B1(G301), .B2(G286), .C1(new_n878), .C2(new_n879), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n966), .B1(G301), .B2(G286), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n880), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n965), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n939), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(new_n971), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n933), .A2(new_n927), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT111), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n972), .B(new_n975), .C1(new_n973), .C2(new_n971), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT43), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n971), .A2(new_n973), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n970), .B1(new_n946), .B2(new_n947), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n976), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AND4_X1   g557(.A1(KEYINPUT43), .A2(new_n978), .A3(new_n982), .A4(new_n890), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT44), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n977), .B2(new_n978), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n986), .A2(new_n978), .A3(new_n982), .A4(new_n890), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n989), .ZN(G397));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n491), .A2(KEYINPUT4), .A3(new_n493), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n465), .ZN(new_n997));
  NAND3_X1  g572(.A1(KEYINPUT67), .A2(G113), .A3(G2104), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G125), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n476), .B2(new_n477), .ZN(new_n1001));
  OAI21_X1  g576(.A(G2105), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n471), .A2(new_n473), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(G40), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(G160), .A2(KEYINPUT112), .A3(G40), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n996), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n805), .B(new_n815), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n846), .B(new_n849), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n729), .B(G1996), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(G1986), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n995), .A2(G1384), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n992), .B2(new_n993), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT45), .B1(new_n501), .B2(new_n991), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT113), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT112), .B1(G160), .B2(G40), .ZN(new_n1023));
  AND4_X1   g598(.A1(KEYINPUT112), .A2(new_n1002), .A3(new_n1003), .A4(G40), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(new_n996), .A3(new_n1026), .A4(new_n1019), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT124), .B(new_n1017), .C1(new_n1028), .C2(G2078), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT124), .ZN(new_n1030));
  AOI21_X1  g605(.A(G2078), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(KEYINPUT53), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n1034), .B2(new_n494), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n994), .A2(KEYINPUT50), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1037), .A2(new_n1025), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1019), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n996), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n501), .A2(KEYINPUT118), .A3(new_n1018), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1017), .A2(G2078), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n744), .A2(new_n1040), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(G301), .B1(new_n1033), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G301), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT125), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1004), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n996), .B2(new_n1052), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1021), .A2(KEYINPUT125), .A3(new_n1004), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1019), .A2(new_n1047), .ZN(new_n1056));
  OAI22_X1  g631(.A1(new_n1055), .A2(new_n1056), .B1(G1961), .B2(new_n1039), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n1050), .B(new_n1057), .C1(new_n1029), .C2(new_n1032), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1016), .B1(new_n1049), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1022), .A2(new_n1027), .A3(new_n825), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1008), .B1(KEYINPUT50), .B2(new_n994), .ZN(new_n1061));
  INV_X1    g636(.A(G2090), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n1037), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(G8), .ZN(new_n1065));
  OAI211_X1 g640(.A(KEYINPUT55), .B(G8), .C1(new_n524), .C2(new_n530), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT114), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n1068));
  INV_X1    g643(.A(G8), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(G166), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n1071));
  NAND4_X1  g646(.A1(G303), .A2(new_n1071), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1067), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1065), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1981), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n607), .A2(new_n608), .A3(new_n615), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G86), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n598), .B1(new_n874), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(G1981), .B1(new_n1078), .B2(new_n606), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(KEYINPUT49), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1076), .A2(KEYINPUT116), .A3(KEYINPUT49), .A4(new_n1079), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT49), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1035), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G8), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n594), .A2(G1976), .A3(new_n596), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1086), .A2(G8), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT52), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1090), .A2(new_n1092), .B1(G288), .B2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1084), .A2(new_n1088), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1069), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1067), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1074), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n777), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n734), .A2(new_n1037), .A3(new_n1025), .A4(new_n1038), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(KEYINPUT119), .B(new_n777), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1103), .A2(G168), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G8), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1044), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1041), .A2(new_n1019), .B1(new_n994), .B2(new_n995), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1966), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1104), .B1(new_n1111), .B2(KEYINPUT119), .ZN(new_n1112));
  AOI21_X1  g687(.A(G168), .B1(new_n1112), .B2(new_n1103), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT51), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1107), .A2(new_n1115), .A3(G8), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1100), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1033), .A2(G301), .A3(new_n1048), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1057), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1118), .B(KEYINPUT54), .C1(new_n550), .C2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1059), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n578), .A2(KEYINPUT120), .A3(new_n580), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n582), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n581), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1956), .B1(new_n1061), .B2(new_n1037), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1025), .A2(new_n996), .A3(new_n1019), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1125), .B(new_n1126), .C1(new_n1127), .C2(new_n1131), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1039), .A2(G1348), .B1(G2067), .B2(new_n1086), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT121), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n1135));
  OAI221_X1 g710(.A(new_n1135), .B1(G2067), .B2(new_n1086), .C1(new_n1039), .C2(G1348), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1132), .B1(new_n1137), .B2(new_n633), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1128), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1129), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1025), .A2(new_n1038), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1037), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n791), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1138), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1132), .A2(new_n1147), .A3(new_n1145), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1147), .B1(new_n1132), .B2(new_n1145), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n1150));
  INV_X1    g725(.A(G1996), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1025), .A2(new_n996), .A3(new_n1151), .A4(new_n1019), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT58), .B(G1341), .Z(new_n1155));
  AOI22_X1  g730(.A1(new_n1152), .A2(new_n1153), .B1(new_n1086), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1150), .B1(new_n1157), .B2(new_n563), .ZN(new_n1158));
  AOI211_X1 g733(.A(KEYINPUT59), .B(new_n562), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1148), .A2(new_n1149), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT123), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n1162));
  OAI221_X1 g737(.A(new_n1162), .B1(new_n1158), .B2(new_n1159), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n633), .B1(new_n1137), .B2(KEYINPUT60), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT60), .ZN(new_n1165));
  AOI211_X1 g740(.A(new_n1165), .B(new_n632), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1164), .A2(new_n1166), .B1(KEYINPUT60), .B2(new_n1137), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1161), .A2(new_n1163), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1121), .B1(new_n1146), .B2(new_n1168), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1087), .B(new_n1085), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1170));
  OR2_X1    g745(.A1(G288), .A2(G1976), .ZN(new_n1171));
  OAI211_X1 g746(.A(KEYINPUT117), .B(new_n1076), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT117), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1171), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1076), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1087), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1172), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1181));
  AOI211_X1 g756(.A(new_n1069), .B(G286), .C1(new_n1112), .C2(new_n1103), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1181), .A2(new_n1074), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1181), .A2(KEYINPUT63), .A3(new_n1074), .A4(new_n1182), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1180), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT62), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1114), .A2(new_n1190), .A3(new_n1116), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1049), .A2(new_n1074), .A3(new_n1181), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1189), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1187), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1015), .B1(new_n1169), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1009), .A2(new_n1151), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT46), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1010), .A2(new_n729), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n1009), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  XOR2_X1   g775(.A(new_n1200), .B(KEYINPUT126), .Z(new_n1201));
  OR2_X1    g776(.A1(new_n1201), .A2(KEYINPUT47), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(KEYINPUT47), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n847), .A2(new_n849), .ZN(new_n1205));
  OAI22_X1  g780(.A1(new_n1204), .A2(new_n1205), .B1(G2067), .B2(new_n805), .ZN(new_n1206));
  NOR4_X1   g781(.A1(new_n996), .A2(new_n1008), .A3(G1986), .A4(G290), .ZN(new_n1207));
  XNOR2_X1  g782(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1207), .B(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1013), .A2(new_n1009), .ZN(new_n1210));
  AOI22_X1  g785(.A1(new_n1206), .A2(new_n1009), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AND3_X1   g786(.A1(new_n1202), .A2(new_n1203), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1195), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g788(.A1(G319), .A2(new_n690), .ZN(new_n1215));
  NOR3_X1   g789(.A1(G229), .A2(G401), .A3(new_n1215), .ZN(new_n1216));
  OAI211_X1 g790(.A(new_n917), .B(new_n1216), .C1(new_n987), .C2(new_n988), .ZN(G225));
  INV_X1    g791(.A(G225), .ZN(G308));
endmodule


