//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955;
  AOI21_X1  g000(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT98), .ZN(new_n203));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT8), .ZN(new_n206));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT99), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT99), .A2(G99gat), .A3(G106gat), .ZN(new_n210));
  INV_X1    g009(.A(G85gat), .ZN(new_n211));
  INV_X1    g010(.A(G92gat), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT100), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT7), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G99gat), .B(G106gat), .Z(new_n219));
  OR2_X1    g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT101), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n219), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n218), .A2(KEYINPUT101), .A3(new_n219), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G36gat), .ZN(new_n226));
  AND2_X1   g025(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G29gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT15), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(KEYINPUT15), .ZN(new_n234));
  XNOR2_X1  g033(.A(G43gat), .B(G50gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n234), .B2(new_n235), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n225), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(KEYINPUT17), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(new_n224), .A3(new_n223), .ZN(new_n240));
  NAND3_X1  g039(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(G190gat), .B(G218gat), .Z(new_n243));
  OR2_X1    g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n243), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n205), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(new_n205), .A3(new_n245), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G15gat), .B(G22gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT16), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n251), .B1(new_n252), .B2(G1gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(G1gat), .B2(new_n251), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G8gat), .ZN(new_n255));
  AND2_X1   g054(.A1(G71gat), .A2(G78gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(G71gat), .A2(G78gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(G57gat), .B(G64gat), .Z(new_n259));
  INV_X1    g058(.A(KEYINPUT94), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(KEYINPUT9), .B2(new_n256), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n262), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT97), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n255), .B1(new_n267), .B2(KEYINPUT21), .ZN(new_n268));
  INV_X1    g067(.A(new_n265), .ZN(new_n269));
  XOR2_X1   g068(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G127gat), .B(G155gat), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n268), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G231gat), .A2(G233gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT96), .ZN(new_n276));
  XOR2_X1   g075(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G183gat), .B(G211gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n274), .B(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT102), .B1(new_n250), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G113gat), .B(G141gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G197gat), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT11), .B(G169gat), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n286), .B(KEYINPUT12), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n255), .B(KEYINPUT91), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n239), .A2(new_n289), .B1(new_n255), .B2(new_n237), .ZN(new_n290));
  NAND2_X1  g089(.A1(G229gat), .A2(G233gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(KEYINPUT18), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n237), .B(new_n255), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n291), .B(KEYINPUT13), .Z(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT92), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n290), .A2(new_n291), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT18), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n296), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(KEYINPUT92), .A3(new_n299), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n288), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT93), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n300), .A2(new_n288), .A3(new_n295), .A4(new_n292), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT93), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT102), .ZN(new_n310));
  INV_X1    g109(.A(new_n281), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n249), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n223), .A2(new_n269), .A3(new_n224), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT10), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n220), .A2(new_n265), .A3(new_n222), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n225), .A2(KEYINPUT10), .A3(new_n267), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G230gat), .A2(G233gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(new_n313), .B2(new_n315), .ZN(new_n321));
  XOR2_X1   g120(.A(G120gat), .B(G148gat), .Z(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT103), .ZN(new_n323));
  XNOR2_X1  g122(.A(G176gat), .B(G204gat), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  NOR2_X1   g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n319), .B(KEYINPUT104), .Z(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(new_n316), .B2(new_n317), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n325), .B1(new_n329), .B2(new_n321), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n282), .A2(new_n309), .A3(new_n312), .A4(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G78gat), .B(G106gat), .ZN(new_n334));
  INV_X1    g133(.A(G50gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n341));
  INV_X1    g140(.A(G141gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT79), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G141gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n345), .A3(G148gat), .ZN(new_n346));
  INV_X1    g145(.A(G148gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G141gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT2), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n342), .A2(G148gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n348), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n351), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n353), .A2(new_n350), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n349), .A2(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n341), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n346), .A2(new_n348), .B1(new_n354), .B2(new_n352), .ZN(new_n363));
  XNOR2_X1  g162(.A(G155gat), .B(G162gat), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n351), .B2(new_n357), .ZN(new_n365));
  NOR4_X1   g164(.A1(new_n363), .A2(new_n365), .A3(KEYINPUT80), .A4(KEYINPUT3), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n340), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G211gat), .A2(G218gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT22), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G197gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT74), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT74), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G197gat), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n372), .A2(new_n374), .A3(G204gat), .ZN(new_n375));
  AOI21_X1  g174(.A(G204gat), .B1(new_n372), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n370), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G211gat), .ZN(new_n378));
  INV_X1    g177(.A(G218gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n368), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(KEYINPUT75), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  OAI221_X1 g182(.A(new_n370), .B1(KEYINPUT75), .B2(new_n381), .C1(new_n375), .C2(new_n376), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n377), .B2(new_n381), .ZN(new_n388));
  INV_X1    g187(.A(new_n381), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n389), .B(new_n370), .C1(new_n375), .C2(new_n376), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT3), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT84), .B1(new_n391), .B2(new_n360), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n381), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(new_n340), .A3(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n361), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n396));
  XNOR2_X1  g195(.A(G141gat), .B(G148gat), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n359), .B1(new_n397), .B2(KEYINPUT2), .ZN(new_n398));
  INV_X1    g197(.A(new_n348), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT79), .B(G141gat), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(G148gat), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n353), .B1(new_n351), .B2(new_n350), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n398), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n396), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n387), .A2(new_n392), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G22gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n385), .A2(new_n340), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n361), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n410), .B2(new_n403), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n361), .B(new_n398), .C1(new_n401), .C2(new_n402), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT80), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n349), .A2(new_n355), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n414), .A2(new_n341), .A3(new_n361), .A4(new_n398), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT85), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n386), .B1(new_n416), .B2(KEYINPUT85), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n411), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n407), .A2(new_n408), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n408), .B1(new_n407), .B2(new_n420), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n339), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n360), .B1(new_n394), .B2(new_n361), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n386), .A2(new_n367), .B1(new_n424), .B2(new_n396), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n425), .A2(new_n392), .B1(G228gat), .B2(G233gat), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT3), .B1(new_n385), .B2(new_n340), .ZN(new_n427));
  OAI211_X1 g226(.A(G228gat), .B(G233gat), .C1(new_n427), .C2(new_n360), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n385), .B1(new_n367), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n417), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(G22gat), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n407), .A2(new_n420), .A3(new_n408), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n338), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n423), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT35), .ZN(new_n436));
  INV_X1    g235(.A(G134gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G127gat), .ZN(new_n438));
  INV_X1    g237(.A(G127gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G134gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT1), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT70), .ZN(new_n443));
  INV_X1    g242(.A(G120gat), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(G113gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(G113gat), .ZN(new_n446));
  INV_X1    g245(.A(G113gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n442), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n438), .A2(new_n440), .ZN(new_n451));
  XNOR2_X1  g250(.A(G113gat), .B(G120gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(KEYINPUT1), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n360), .B(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(G225gat), .A2(G233gat), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT5), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n413), .A2(new_n415), .ZN(new_n458));
  INV_X1    g257(.A(new_n446), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n444), .A2(G113gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n441), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n461), .A2(new_n451), .B1(new_n442), .B2(new_n449), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(KEYINPUT3), .B2(new_n403), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n465));
  NAND3_X1  g264(.A1(new_n360), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n403), .A2(new_n454), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n466), .B(KEYINPUT82), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n360), .A2(new_n462), .A3(new_n465), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT82), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n464), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n456), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n457), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n465), .B1(new_n403), .B2(new_n454), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(KEYINPUT5), .A3(new_n456), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(KEYINPUT4), .B2(new_n467), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n464), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G1gat), .B(G29gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(KEYINPUT0), .ZN(new_n482));
  XNOR2_X1  g281(.A(G57gat), .B(G85gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n458), .A2(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n487), .A2(new_n456), .A3(new_n469), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n488), .A2(new_n457), .B1(new_n464), .B2(new_n478), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n484), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(KEYINPUT6), .A3(new_n484), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n495));
  AND2_X1   g294(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT23), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(G169gat), .ZN(new_n500));
  INV_X1    g299(.A(G169gat), .ZN(new_n501));
  INV_X1    g300(.A(G176gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G169gat), .A2(G176gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT23), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n498), .A2(new_n500), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(G183gat), .A2(G190gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT64), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n510), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT64), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT25), .B1(new_n506), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(new_n512), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT25), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n505), .B2(new_n503), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT66), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(new_n501), .A3(new_n502), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(KEYINPUT23), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT67), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n509), .A2(new_n511), .A3(new_n513), .ZN(new_n526));
  OR2_X1    g325(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n500), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n505), .A2(new_n503), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n517), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT67), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n523), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT26), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT68), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT68), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT26), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n536), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n504), .A2(new_n535), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n503), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n539), .A2(new_n541), .B1(G183gat), .B2(G190gat), .ZN(new_n542));
  INV_X1    g341(.A(G183gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT27), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT27), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G183gat), .ZN(new_n546));
  INV_X1    g345(.A(G190gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT28), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G183gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(KEYINPUT28), .A3(new_n547), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT69), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n542), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n542), .B2(new_n553), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n525), .B(new_n534), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G226gat), .A2(G233gat), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(KEYINPUT76), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n532), .A2(new_n523), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n542), .A2(new_n553), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT29), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT77), .B1(new_n564), .B2(new_n560), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT77), .ZN(new_n566));
  INV_X1    g365(.A(new_n560), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n532), .A2(new_n523), .B1(new_n553), .B2(new_n542), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(KEYINPUT29), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n561), .A2(new_n565), .A3(new_n385), .A4(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n560), .A2(KEYINPUT29), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n558), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n560), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n386), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G8gat), .B(G36gat), .Z(new_n576));
  XOR2_X1   g375(.A(G64gat), .B(G92gat), .Z(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n495), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n570), .A2(new_n574), .A3(KEYINPUT30), .A4(new_n578), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n578), .B(KEYINPUT78), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n435), .A2(new_n436), .A3(new_n494), .A4(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n525), .A2(new_n534), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT71), .ZN(new_n587));
  INV_X1    g386(.A(new_n557), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n555), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n586), .A2(new_n587), .A3(new_n454), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n454), .A2(new_n587), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n462), .A2(KEYINPUT71), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n558), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G227gat), .ZN(new_n594));
  INV_X1    g393(.A(G233gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT32), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT33), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G15gat), .B(G43gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT72), .ZN(new_n602));
  XNOR2_X1  g401(.A(G71gat), .B(G99gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  NAND3_X1  g403(.A1(new_n598), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n597), .B(KEYINPUT32), .C1(new_n599), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n596), .B1(new_n590), .B2(new_n593), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT34), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI211_X1 g410(.A(KEYINPUT34), .B(new_n596), .C1(new_n590), .C2(new_n593), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT73), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n608), .A2(new_n613), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n611), .A2(new_n612), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(new_n605), .A3(new_n607), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(KEYINPUT73), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n585), .B1(new_n615), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n618), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n421), .A2(new_n422), .A3(new_n339), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n338), .B1(new_n432), .B2(new_n433), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT90), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n494), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT90), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n435), .A2(new_n616), .A3(new_n629), .A4(new_n618), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n620), .B1(new_n631), .B2(KEYINPUT35), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT86), .B(KEYINPUT40), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n456), .B1(new_n487), .B2(new_n469), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n484), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n473), .A2(new_n474), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n635), .B1(new_n455), .B2(new_n456), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n633), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT87), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n473), .A2(new_n635), .A3(new_n474), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n639), .A2(KEYINPUT40), .A3(new_n485), .A4(new_n642), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n640), .A2(new_n641), .B1(new_n643), .B2(KEYINPUT88), .ZN(new_n644));
  INV_X1    g443(.A(new_n633), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n485), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n455), .A2(new_n456), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT39), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n473), .B2(new_n474), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n645), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n650), .A2(KEYINPUT87), .B1(new_n484), .B2(new_n489), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT88), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n636), .A2(new_n652), .A3(KEYINPUT40), .A4(new_n639), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n644), .A2(new_n651), .A3(new_n627), .A4(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n655));
  NAND3_X1  g454(.A1(new_n570), .A2(new_n574), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n579), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT37), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n570), .B2(new_n574), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT38), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n582), .A2(new_n661), .ZN(new_n662));
  AOI22_X1  g461(.A1(new_n558), .A2(new_n571), .B1(new_n560), .B2(new_n568), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n658), .B1(new_n663), .B2(new_n385), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n561), .A2(new_n565), .A3(new_n386), .A4(new_n569), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n570), .A2(new_n574), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n666), .A2(new_n656), .B1(new_n667), .B2(new_n578), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n660), .A2(new_n668), .A3(new_n493), .A4(new_n492), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n435), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n621), .A2(KEYINPUT36), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT36), .B1(new_n619), .B2(new_n615), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n632), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n333), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n626), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT105), .B(G1gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1324gat));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n627), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n681), .A2(G8gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT16), .B(G8gat), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT42), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(KEYINPUT42), .B2(new_n684), .ZN(G1325gat));
  NAND2_X1  g485(.A1(new_n619), .A2(new_n615), .ZN(new_n687));
  AOI21_X1  g486(.A(G15gat), .B1(new_n677), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n674), .A2(new_n673), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G15gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT106), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n688), .B1(new_n677), .B2(new_n692), .ZN(G1326gat));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n624), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT43), .B(G22gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  OAI21_X1  g495(.A(new_n250), .B1(new_n632), .B2(new_n675), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n308), .A2(new_n311), .A3(new_n331), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(G29gat), .A3(new_n494), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT45), .Z(new_n702));
  AND2_X1   g501(.A1(new_n697), .A2(KEYINPUT44), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n249), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n247), .A2(KEYINPUT107), .A3(new_n248), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n704), .B(new_n708), .C1(new_n632), .C2(new_n675), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n699), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n711), .A2(new_n494), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n713), .A2(KEYINPUT108), .ZN(new_n714));
  OAI21_X1  g513(.A(G29gat), .B1(new_n713), .B2(KEYINPUT108), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n702), .B1(new_n714), .B2(new_n715), .ZN(G1328gat));
  NOR3_X1   g515(.A1(new_n700), .A2(G36gat), .A3(new_n584), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT46), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n711), .A2(new_n584), .A3(new_n712), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n226), .B2(new_n719), .ZN(G1329gat));
  NOR2_X1   g519(.A1(new_n711), .A2(new_n712), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(G43gat), .A3(new_n690), .ZN(new_n722));
  INV_X1    g521(.A(new_n687), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n700), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(G43gat), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1330gat));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n435), .B1(new_n700), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n728), .B2(new_n700), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n435), .A2(new_n335), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n730), .A2(new_n335), .B1(new_n721), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g532(.A1(new_n282), .A2(new_n312), .A3(new_n308), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n676), .A2(new_n734), .A3(new_n332), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n626), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n627), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT49), .B(G64gat), .Z(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n738), .B2(new_n740), .ZN(G1333gat));
  INV_X1    g540(.A(new_n735), .ZN(new_n742));
  OAI21_X1  g541(.A(G71gat), .B1(new_n742), .B2(new_n689), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n723), .A2(G71gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1334gat));
  NAND2_X1  g546(.A1(new_n735), .A2(new_n624), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT112), .B(G78gat), .Z(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1335gat));
  NAND3_X1  g549(.A1(new_n308), .A2(new_n281), .A3(new_n331), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n703), .B2(new_n710), .ZN(new_n753));
  OAI21_X1  g552(.A(G85gat), .B1(new_n753), .B2(new_n494), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n309), .A2(new_n311), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n698), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT51), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n698), .A2(new_n758), .A3(new_n755), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n331), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n626), .A2(new_n211), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n754), .B1(new_n760), .B2(new_n761), .ZN(G1336gat));
  NOR2_X1   g561(.A1(new_n584), .A2(G92gat), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n757), .A2(new_n331), .A3(new_n759), .A4(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n697), .A2(KEYINPUT44), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n584), .B(new_n751), .C1(new_n766), .C2(new_n709), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n764), .B(new_n765), .C1(new_n212), .C2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n767), .B2(new_n212), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n627), .B(new_n752), .C1(new_n703), .C2(new_n710), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(KEYINPUT113), .A3(G92gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n772), .A3(new_n764), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n773), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT114), .B1(new_n773), .B2(KEYINPUT52), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n768), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT115), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n778), .B(new_n768), .C1(new_n774), .C2(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1337gat));
  INV_X1    g579(.A(G99gat), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n753), .A2(new_n781), .A3(new_n689), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n760), .A2(new_n723), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n781), .ZN(G1338gat));
  INV_X1    g583(.A(G106gat), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n753), .A2(new_n435), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787));
  OAI221_X1 g586(.A(new_n785), .B1(new_n760), .B2(new_n435), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(G106gat), .B1(new_n786), .B2(KEYINPUT116), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT53), .Z(G1339gat));
  NOR2_X1   g590(.A1(new_n734), .A2(new_n331), .ZN(new_n792));
  INV_X1    g591(.A(new_n328), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n320), .B(KEYINPUT54), .C1(new_n793), .C2(new_n318), .ZN(new_n794));
  INV_X1    g593(.A(new_n325), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n329), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n798), .A2(new_n799), .B1(new_n320), .B2(new_n326), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n290), .A2(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n286), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n306), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n794), .A2(KEYINPUT55), .A3(new_n797), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n708), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n303), .A2(new_n307), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n800), .A3(new_n305), .A4(new_n804), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n803), .A2(new_n331), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n708), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n809), .B1(new_n808), .B2(new_n810), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n806), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n792), .B1(new_n815), .B2(new_n281), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n625), .A2(new_n630), .ZN(new_n817));
  NOR4_X1   g616(.A1(new_n816), .A2(new_n494), .A3(new_n627), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n447), .A3(new_n309), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n816), .A2(new_n723), .A3(new_n624), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n494), .A2(new_n627), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n309), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(KEYINPUT118), .A3(G113gat), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT118), .B1(new_n822), .B2(G113gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n819), .B1(new_n824), .B2(new_n825), .ZN(G1340gat));
  NAND3_X1  g625(.A1(new_n818), .A2(new_n444), .A3(new_n331), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n820), .A2(new_n331), .A3(new_n821), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(KEYINPUT119), .A3(G120gat), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT119), .B1(new_n828), .B2(G120gat), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(G1341gat));
  NAND2_X1  g631(.A1(new_n820), .A2(new_n821), .ZN(new_n833));
  OAI21_X1  g632(.A(G127gat), .B1(new_n833), .B2(new_n281), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n439), .A3(new_n311), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1342gat));
  NAND3_X1  g635(.A1(new_n818), .A2(new_n437), .A3(new_n250), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n838));
  OAI21_X1  g637(.A(G134gat), .B1(new_n833), .B2(new_n249), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G1343gat));
  NAND2_X1  g640(.A1(new_n689), .A2(new_n821), .ZN(new_n842));
  INV_X1    g641(.A(new_n792), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n808), .A2(new_n810), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n844), .A2(new_n249), .B1(new_n805), .B2(new_n708), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n845), .B2(new_n311), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n435), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n847), .B1(new_n846), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n848), .B1(new_n816), .B2(new_n435), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n842), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n400), .B1(new_n854), .B2(new_n309), .ZN(new_n855));
  INV_X1    g654(.A(new_n816), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n690), .A2(new_n627), .A3(new_n435), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n856), .A2(new_n626), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n342), .A3(new_n309), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT58), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n308), .B(new_n842), .C1(new_n852), .C2(new_n853), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n859), .B(new_n862), .C1(new_n863), .C2(new_n400), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(G1344gat));
  AND4_X1   g664(.A1(new_n626), .A2(new_n856), .A3(new_n331), .A4(new_n857), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n347), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n851), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n842), .A2(new_n332), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n867), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n849), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n816), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n250), .B1(new_n808), .B2(new_n810), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n876), .B1(new_n250), .B2(new_n805), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n843), .B1(new_n877), .B2(new_n311), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n878), .B2(new_n624), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n872), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n868), .A2(new_n873), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT121), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n873), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1345gat));
  INV_X1    g685(.A(G155gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n858), .A2(new_n887), .A3(new_n311), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n854), .A2(new_n311), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n887), .ZN(G1346gat));
  INV_X1    g689(.A(G162gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n858), .A2(new_n891), .A3(new_n250), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n854), .A2(new_n708), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n891), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n816), .A2(new_n626), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n895), .A2(new_n627), .A3(new_n625), .A4(new_n630), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n501), .B1(new_n896), .B2(new_n308), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n723), .A2(new_n624), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n626), .A2(new_n584), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n844), .A2(KEYINPUT117), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n812), .A3(new_n811), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n311), .B1(new_n901), .B2(new_n806), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n898), .B(new_n899), .C1(new_n902), .C2(new_n792), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n856), .A2(KEYINPUT122), .A3(new_n898), .A4(new_n899), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n905), .A2(new_n906), .A3(G169gat), .A4(new_n309), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n897), .A2(new_n907), .ZN(G1348gat));
  OAI21_X1  g707(.A(new_n502), .B1(new_n896), .B2(new_n332), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n332), .A2(new_n498), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n905), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n909), .A2(new_n911), .ZN(G1349gat));
  NAND3_X1  g711(.A1(new_n905), .A2(new_n906), .A3(new_n311), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G183gat), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n311), .A2(new_n551), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n896), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT60), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n914), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1350gat));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n250), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n922), .A2(new_n923), .A3(G190gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n922), .B2(G190gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n708), .A2(new_n547), .ZN(new_n926));
  OAI22_X1  g725(.A1(new_n924), .A2(new_n925), .B1(new_n896), .B2(new_n926), .ZN(G1351gat));
  NAND4_X1  g726(.A1(new_n895), .A2(new_n689), .A3(new_n627), .A4(new_n624), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n928), .A2(KEYINPUT123), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(KEYINPUT123), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g730(.A(KEYINPUT124), .B(G197gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n309), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n689), .A2(new_n899), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n934), .B1(new_n875), .B2(new_n879), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(new_n308), .ZN(new_n936));
  OAI22_X1  g735(.A1(new_n931), .A2(new_n933), .B1(new_n936), .B2(new_n932), .ZN(G1352gat));
  OR2_X1    g736(.A1(new_n332), .A2(G204gat), .ZN(new_n938));
  XOR2_X1   g737(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  OR3_X1    g739(.A1(new_n928), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(G204gat), .B1(new_n935), .B2(new_n332), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n940), .B1(new_n928), .B2(new_n938), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G1353gat));
  NAND2_X1  g743(.A1(new_n311), .A2(new_n378), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n311), .B(new_n934), .C1(new_n875), .C2(new_n879), .ZN(new_n946));
  AND4_X1   g745(.A1(KEYINPUT126), .A2(new_n946), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n947));
  OAI21_X1  g746(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AOI22_X1  g748(.A1(new_n946), .A2(new_n949), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n950));
  OAI22_X1  g749(.A1(new_n931), .A2(new_n945), .B1(new_n947), .B2(new_n950), .ZN(G1354gat));
  NOR2_X1   g750(.A1(new_n249), .A2(new_n379), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT127), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n935), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n929), .A2(new_n708), .A3(new_n930), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n379), .ZN(G1355gat));
endmodule


