//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT0), .B(G128), .Z(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(KEYINPUT64), .A3(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G143), .B(G146), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  OAI211_X1 g011(.A(KEYINPUT0), .B(G128), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n200), .B(KEYINPUT89), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT92), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT90), .B(G224), .Z(new_n203));
  OR2_X1    g017(.A1(new_n203), .A2(G953), .ZN(new_n204));
  AOI22_X1  g018(.A1(new_n201), .A2(new_n202), .B1(KEYINPUT7), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n194), .A2(new_n206), .A3(G128), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n191), .B(new_n193), .C1(KEYINPUT1), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n201), .B1(G125), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n205), .B(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G104), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G107), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT3), .B1(new_n217), .B2(G107), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT78), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n215), .A3(G104), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT79), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n225), .A2(new_n215), .A3(KEYINPUT79), .A4(G104), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(G101), .B1(new_n217), .B2(G107), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n224), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT81), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n222), .A2(new_n223), .B1(new_n228), .B2(new_n229), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(new_n231), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n219), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT2), .B(G113), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G116), .B(G119), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(KEYINPUT66), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n242));
  INV_X1    g056(.A(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G116), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n242), .B1(new_n247), .B2(new_n238), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n240), .A2(KEYINPUT5), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n250), .B(G113), .C1(KEYINPUT5), .C2(new_n244), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n237), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(G110), .B(G122), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n254), .B(KEYINPUT8), .Z(new_n255));
  OR2_X1    g069(.A1(new_n251), .A2(KEYINPUT86), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n251), .A2(KEYINPUT86), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n256), .A2(new_n249), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n219), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n235), .B1(new_n234), .B2(new_n231), .ZN(new_n260));
  AND4_X1   g074(.A1(new_n235), .A2(new_n224), .A3(new_n230), .A4(new_n231), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n255), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n213), .B1(new_n253), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n249), .B1(new_n240), .B2(new_n239), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n224), .A2(new_n230), .A3(new_n218), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G101), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(G101), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT80), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT80), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(new_n272), .A3(G101), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT4), .B1(new_n260), .B2(new_n261), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT85), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n258), .A2(new_n237), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n267), .B1(new_n233), .B2(new_n236), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n271), .A3(new_n273), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT85), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n269), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n277), .A2(new_n254), .A3(new_n278), .A4(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(G902), .B1(new_n264), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(KEYINPUT6), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n265), .A2(new_n268), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n266), .A2(new_n272), .A3(G101), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n272), .B1(new_n266), .B2(G101), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n286), .B1(new_n289), .B2(new_n279), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n290), .A2(new_n281), .B1(new_n237), .B2(new_n258), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n254), .B1(new_n291), .B2(new_n277), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT87), .B1(new_n285), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n254), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n282), .A2(new_n278), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n290), .A2(new_n281), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT87), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT6), .A4(new_n283), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT88), .B(KEYINPUT6), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n294), .B(new_n301), .C1(new_n295), .C2(new_n296), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n212), .B(new_n204), .Z(new_n303));
  AND4_X1   g117(.A1(KEYINPUT91), .A2(new_n300), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n302), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n305), .B1(new_n293), .B2(new_n299), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT91), .B1(new_n306), .B2(new_n303), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n284), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G210), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n309), .B(new_n284), .C1(new_n304), .C2(new_n307), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n188), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  XOR2_X1   g128(.A(new_n314), .B(KEYINPUT69), .Z(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT11), .ZN(new_n317));
  INV_X1    g131(.A(G134), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(G137), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT11), .A3(G134), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(G137), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G131), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT65), .B(G131), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n325), .A2(new_n319), .A3(new_n321), .A4(new_n322), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n198), .A3(new_n195), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT30), .ZN(new_n329));
  INV_X1    g143(.A(new_n322), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n318), .A2(G137), .ZN(new_n331));
  OAI21_X1  g145(.A(G131), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n326), .A2(new_n207), .A3(new_n332), .A4(new_n209), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n328), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n329), .B1(new_n328), .B2(new_n333), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n265), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G237), .ZN(new_n337));
  INV_X1    g151(.A(G953), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(G210), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT27), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G101), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n324), .A2(new_n326), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n333), .B1(new_n343), .B2(new_n199), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(new_n265), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT31), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT67), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n336), .A2(KEYINPUT67), .A3(new_n342), .A4(new_n346), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n350), .B1(new_n354), .B2(KEYINPUT31), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n344), .A2(new_n265), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(KEYINPUT68), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT68), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n344), .B2(new_n265), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n346), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT28), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n346), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n342), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(KEYINPUT32), .B(new_n316), .C1(new_n355), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT73), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n363), .ZN(new_n367));
  INV_X1    g181(.A(new_n342), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(new_n350), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT73), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT32), .A4(new_n316), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n366), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n346), .A2(new_n356), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(new_n362), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT72), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT72), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n363), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n377), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n342), .A2(KEYINPUT29), .ZN(new_n381));
  AOI21_X1  g195(.A(G902), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT71), .B1(new_n367), .B2(new_n368), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT71), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n361), .A2(new_n384), .A3(new_n342), .A4(new_n363), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n344), .A2(KEYINPUT30), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n328), .A2(new_n329), .A3(new_n333), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n345), .B1(new_n388), .B2(new_n265), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT29), .B1(new_n390), .B2(new_n368), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n383), .A2(new_n385), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n382), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G472), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT70), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT67), .B1(new_n389), .B2(new_n342), .ZN(new_n396));
  INV_X1    g210(.A(new_n353), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT31), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n364), .B1(new_n398), .B2(new_n349), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n395), .B1(new_n399), .B2(new_n315), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n371), .A2(KEYINPUT70), .A3(new_n316), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT32), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n374), .A2(new_n394), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G217), .ZN(new_n405));
  INV_X1    g219(.A(G902), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n405), .B1(G234), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G125), .B(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT16), .ZN(new_n410));
  INV_X1    g224(.A(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G125), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(KEYINPUT16), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n190), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT75), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n410), .B(G146), .C1(KEYINPUT16), .C2(new_n412), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n413), .A2(KEYINPUT75), .A3(new_n190), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n208), .A2(G119), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n243), .A2(G128), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(KEYINPUT24), .B(G110), .Z(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT74), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT74), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .ZN(new_n427));
  INV_X1    g241(.A(new_n419), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n427), .B(new_n420), .C1(new_n428), .C2(KEYINPUT23), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n424), .A2(new_n426), .B1(G110), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n417), .A2(new_n418), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n409), .B(KEYINPUT76), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n190), .ZN(new_n433));
  OAI22_X1  g247(.A1(new_n429), .A2(G110), .B1(new_n421), .B2(new_n422), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n416), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT22), .B(G137), .ZN(new_n437));
  INV_X1    g251(.A(G221), .ZN(new_n438));
  INV_X1    g252(.A(G234), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n438), .A2(new_n439), .A3(G953), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n437), .B(new_n440), .Z(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n431), .A2(new_n435), .A3(new_n441), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n406), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT25), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n446), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n408), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n443), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n451));
  INV_X1    g265(.A(new_n444), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n451), .B1(new_n450), .B2(new_n452), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n407), .A2(G902), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n449), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n404), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT9), .B(G234), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n438), .B1(new_n462), .B2(new_n406), .ZN(new_n463));
  INV_X1    g277(.A(G469), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT10), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n262), .B2(new_n210), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n237), .A2(KEYINPUT10), .A3(new_n211), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n268), .A2(new_n198), .A3(new_n195), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n289), .B2(new_n279), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT83), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n469), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n280), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT83), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n473), .A2(new_n474), .A3(new_n466), .A4(new_n467), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n327), .A3(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n473), .A2(new_n343), .A3(new_n466), .A4(new_n467), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G140), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n338), .A2(G227), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(KEYINPUT82), .A2(KEYINPUT12), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n237), .A2(new_n211), .ZN(new_n485));
  AOI211_X1 g299(.A(new_n210), .B(new_n219), .C1(new_n233), .C2(new_n236), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n327), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n262), .A2(new_n210), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n237), .A2(new_n211), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n343), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  XOR2_X1   g304(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n491));
  OAI21_X1  g305(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n477), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n480), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n483), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n464), .B1(new_n495), .B2(new_n406), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT84), .B(G469), .Z(new_n498));
  AND2_X1   g312(.A1(new_n482), .A2(new_n492), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n481), .B1(new_n476), .B2(new_n477), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n406), .B(new_n498), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n463), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G478), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n245), .A2(G122), .ZN(new_n507));
  INV_X1    g321(.A(G122), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(G116), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n215), .ZN(new_n511));
  XNOR2_X1  g325(.A(G128), .B(G143), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(new_n318), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n508), .A2(KEYINPUT14), .A3(G116), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(new_n508), .B2(G116), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n515), .A2(KEYINPUT97), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(KEYINPUT97), .ZN(new_n517));
  AOI211_X1 g331(.A(new_n507), .B(new_n514), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n511), .B(new_n513), .C1(new_n518), .C2(new_n215), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n510), .B(new_n215), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n192), .A2(G128), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(G134), .C1(new_n523), .C2(new_n521), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n512), .A2(new_n318), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n461), .A2(new_n405), .A3(G953), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n519), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n527), .B1(new_n519), .B2(new_n526), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n406), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT98), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n519), .A2(new_n526), .ZN(new_n534));
  INV_X1    g348(.A(new_n527), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(G902), .B1(new_n536), .B2(new_n528), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT98), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n506), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n505), .B1(new_n531), .B2(new_n532), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n539), .A2(KEYINPUT99), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT99), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n537), .A2(KEYINPUT98), .ZN(new_n543));
  AOI211_X1 g357(.A(new_n532), .B(G902), .C1(new_n536), .C2(new_n528), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n505), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n540), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(G113), .B(G122), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(new_n217), .ZN(new_n551));
  INV_X1    g365(.A(new_n409), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G146), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n433), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n337), .A2(new_n338), .A3(G214), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n192), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n337), .A2(new_n338), .A3(G143), .A4(G214), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(KEYINPUT18), .A2(G131), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n417), .A2(new_n418), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n325), .B1(new_n556), .B2(new_n557), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n556), .A2(new_n325), .A3(new_n557), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n565), .B2(new_n564), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n551), .B(new_n561), .C1(new_n562), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n552), .A2(KEYINPUT19), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT76), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n409), .B(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n190), .B(new_n570), .C1(new_n572), .C2(KEYINPUT19), .ZN(new_n573));
  INV_X1    g387(.A(new_n566), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT93), .B1(new_n574), .B2(new_n563), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n564), .A2(new_n576), .A3(new_n566), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n573), .A2(new_n575), .A3(new_n416), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(KEYINPUT94), .A3(new_n561), .ZN(new_n579));
  INV_X1    g393(.A(new_n551), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT94), .B1(new_n578), .B2(new_n561), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n569), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(G475), .A2(G902), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n569), .B(KEYINPUT95), .C1(new_n581), .C2(new_n582), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n588), .A2(KEYINPUT20), .B1(new_n583), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G475), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n561), .B1(new_n562), .B2(new_n568), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n580), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n569), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n591), .B1(new_n594), .B2(new_n406), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n406), .B(new_n338), .C1(G234), .C2(G237), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT21), .B(G898), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n338), .A2(G952), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n439), .B2(new_n337), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n549), .A2(new_n596), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n503), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n313), .A2(new_n460), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  AND2_X1   g421(.A1(new_n313), .A2(new_n603), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n504), .A2(new_n406), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n537), .B2(new_n504), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT33), .B1(new_n529), .B2(new_n530), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n536), .A2(new_n612), .A3(new_n528), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(G478), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n596), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n400), .A2(new_n401), .ZN(new_n617));
  OAI21_X1  g431(.A(G472), .B1(new_n399), .B2(G902), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n458), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n503), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n608), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  XNOR2_X1  g437(.A(new_n588), .B(KEYINPUT20), .ZN(new_n624));
  INV_X1    g438(.A(new_n595), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n549), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n608), .A2(new_n620), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G107), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT100), .B(KEYINPUT35), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NAND2_X1  g445(.A1(new_n617), .A2(new_n618), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n436), .B(KEYINPUT101), .Z(new_n633));
  OR2_X1    g447(.A1(new_n442), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n449), .B1(new_n635), .B2(new_n457), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n313), .A2(new_n605), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT102), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT37), .B(G110), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n597), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n601), .ZN(new_n644));
  AND4_X1   g458(.A1(new_n625), .A2(new_n548), .A3(new_n624), .A4(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n636), .ZN(new_n646));
  AND4_X1   g460(.A1(new_n404), .A2(new_n502), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n311), .A2(new_n312), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n648), .A3(new_n187), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XNOR2_X1  g464(.A(new_n648), .B(KEYINPUT38), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n644), .B(KEYINPUT39), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n502), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  INV_X1    g470(.A(new_n375), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n354), .B1(new_n368), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(G472), .B1(new_n658), .B2(G902), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n374), .A2(new_n659), .A3(new_n403), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n549), .A2(new_n596), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n187), .A3(new_n636), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n656), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n651), .A2(new_n655), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  INV_X1    g480(.A(new_n615), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n667), .B(new_n644), .C1(new_n590), .C2(new_n595), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n404), .A2(new_n502), .A3(new_n646), .A4(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n648), .A3(new_n187), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G146), .ZN(G48));
  OAI21_X1  g486(.A(new_n406), .B1(new_n499), .B2(new_n500), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G469), .ZN(new_n674));
  INV_X1    g488(.A(new_n463), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n675), .A3(new_n501), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT103), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n674), .A2(new_n678), .A3(new_n675), .A4(new_n501), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n459), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n313), .A3(new_n603), .A4(new_n616), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NAND4_X1  g498(.A1(new_n681), .A2(new_n313), .A3(new_n603), .A4(new_n627), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NAND2_X1  g500(.A1(new_n404), .A2(new_n646), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n604), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n677), .A2(new_n679), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n313), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  XNOR2_X1  g505(.A(new_n458), .B(KEYINPUT104), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n377), .B(new_n368), .C1(new_n376), .C2(new_n379), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n316), .B1(new_n694), .B2(new_n355), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n692), .A2(new_n618), .A3(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n680), .A2(new_n696), .A3(new_n602), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n313), .A3(new_n662), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  OR2_X1    g513(.A1(new_n590), .A2(new_n595), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(KEYINPUT105), .A3(new_n667), .A4(new_n644), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n646), .A2(new_n618), .A3(new_n695), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n668), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n648), .A2(new_n689), .A3(new_n187), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  NAND3_X1  g521(.A1(new_n406), .A2(KEYINPUT106), .A3(G469), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n495), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n496), .B2(KEYINPUT106), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n463), .B1(new_n710), .B2(new_n501), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n311), .A2(new_n187), .A3(new_n312), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n701), .A2(new_n704), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(KEYINPUT42), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n713), .A2(new_n460), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n458), .B(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n394), .A2(new_n365), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n402), .B1(new_n399), .B2(new_n315), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n704), .A3(new_n701), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT42), .B1(new_n722), .B2(new_n712), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(G131), .Z(G33));
  NAND3_X1  g539(.A1(new_n713), .A2(new_n460), .A3(new_n645), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G134), .ZN(G36));
  NAND3_X1  g541(.A1(new_n311), .A2(new_n187), .A3(new_n312), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n700), .A2(KEYINPUT43), .A3(new_n615), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n615), .B1(new_n700), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n731), .B2(new_n700), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n730), .B1(new_n733), .B2(KEYINPUT43), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n632), .A3(new_n646), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n729), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n737), .A2(KEYINPUT108), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(KEYINPUT108), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n464), .B1(new_n495), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n740), .B2(new_n495), .ZN(new_n742));
  NAND2_X1  g556(.A1(G469), .A2(G902), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT46), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n501), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n742), .A2(KEYINPUT46), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n675), .A3(new_n652), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n749), .B1(new_n735), .B2(new_n736), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n738), .A2(new_n739), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT109), .B(G137), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT110), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n751), .B(new_n753), .ZN(G39));
  AOI21_X1  g568(.A(new_n463), .B1(new_n746), .B2(new_n747), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT47), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n404), .A2(new_n458), .A3(new_n668), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n756), .A2(new_n729), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT111), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G140), .ZN(G42));
  NOR2_X1   g574(.A1(new_n696), .A2(new_n601), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n734), .A2(new_n761), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n651), .A2(new_n762), .A3(new_n187), .A4(new_n680), .ZN(new_n763));
  NOR2_X1   g577(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n765), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n674), .A2(new_n501), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n756), .B1(new_n463), .B2(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n770), .A2(new_n728), .A3(new_n762), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n729), .A2(new_n689), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT119), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n601), .B1(new_n772), .B2(KEYINPUT119), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n702), .A2(new_n773), .A3(new_n734), .A4(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n767), .A2(new_n771), .A3(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n773), .A2(new_n774), .A3(new_n458), .A4(new_n661), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT120), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n596), .A2(new_n615), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT51), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n773), .A2(new_n774), .A3(new_n721), .A4(new_n734), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(KEYINPUT121), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(KEYINPUT121), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(KEYINPUT48), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n313), .A2(new_n689), .ZN(new_n786));
  OAI221_X1 g600(.A(new_n600), .B1(new_n786), .B2(new_n762), .C1(new_n784), .C2(KEYINPUT48), .ZN(new_n787));
  INV_X1    g601(.A(new_n778), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n787), .B1(new_n616), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n781), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n713), .A2(new_n705), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n313), .B(new_n605), .C1(new_n460), .C2(new_n637), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n595), .B(new_n590), .C1(new_n545), .C2(new_n546), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n616), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n313), .A2(new_n603), .A3(new_n620), .A4(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n726), .A2(new_n791), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n687), .A2(new_n503), .ZN(new_n798));
  INV_X1    g612(.A(new_n644), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n626), .A2(new_n539), .A3(new_n540), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n311), .A2(new_n187), .A3(new_n312), .A4(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n798), .B1(new_n801), .B2(KEYINPUT113), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(KEYINPUT113), .B2(new_n801), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT116), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n792), .A2(new_n796), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n801), .A2(KEYINPUT113), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n801), .A2(KEYINPUT113), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n798), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n712), .A2(new_n459), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n810), .A2(new_n645), .B1(new_n713), .B2(new_n705), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n805), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n804), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n706), .A2(new_n649), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n646), .A2(new_n799), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n711), .A2(new_n660), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n648), .A3(new_n187), .A4(new_n662), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n313), .B2(new_n670), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n814), .A2(new_n815), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n818), .A2(KEYINPUT52), .A3(new_n671), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n706), .A2(new_n649), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT114), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n818), .A2(new_n706), .A3(new_n649), .A4(new_n671), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n819), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n821), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n682), .A2(new_n698), .A3(new_n685), .A4(new_n690), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n828), .A2(new_n724), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT117), .B1(new_n813), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n804), .A2(new_n812), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n834), .A3(new_n827), .A4(new_n830), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n828), .A2(new_n797), .A3(new_n803), .A4(new_n724), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n826), .B1(new_n823), .B2(new_n822), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n832), .A2(new_n835), .B1(new_n829), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT53), .B1(new_n836), .B2(new_n827), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT115), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n829), .B2(new_n838), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n842), .A2(KEYINPUT115), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n841), .B1(new_n846), .B2(new_n840), .ZN(new_n847));
  OAI22_X1  g661(.A1(new_n790), .A2(new_n847), .B1(G952), .B2(G953), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n692), .A2(new_n187), .A3(new_n675), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n849), .B(new_n733), .C1(KEYINPUT49), .C2(new_n768), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n768), .A2(KEYINPUT49), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT112), .Z(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n661), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n848), .B1(new_n651), .B2(new_n853), .ZN(G75));
  XNOR2_X1  g668(.A(new_n306), .B(new_n303), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT55), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n839), .A2(new_n406), .ZN(new_n857));
  INV_X1    g671(.A(G210), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n856), .B1(new_n859), .B2(KEYINPUT56), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n338), .A2(G952), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n859), .A2(KEYINPUT56), .A3(new_n856), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(G51));
  XOR2_X1   g679(.A(new_n743), .B(KEYINPUT57), .Z(new_n866));
  INV_X1    g680(.A(new_n841), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n839), .A2(new_n840), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n500), .B2(new_n499), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n857), .A2(new_n742), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n861), .B1(new_n870), .B2(new_n871), .ZN(G54));
  INV_X1    g686(.A(new_n857), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n585), .A2(new_n587), .ZN(new_n874));
  NAND2_X1  g688(.A1(KEYINPUT58), .A2(G475), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n874), .B1(new_n873), .B2(new_n876), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n877), .A2(new_n878), .A3(new_n861), .ZN(G60));
  NAND2_X1  g693(.A1(new_n611), .A2(new_n613), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n609), .B(KEYINPUT59), .Z(new_n881));
  AND2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n867), .B2(new_n868), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n883), .A2(new_n884), .A3(new_n862), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n884), .B1(new_n883), .B2(new_n862), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n880), .B1(new_n847), .B2(new_n881), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(G63));
  INV_X1    g702(.A(new_n456), .ZN(new_n889));
  NAND2_X1  g703(.A1(G217), .A2(G902), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT60), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n839), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n862), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n832), .A2(new_n835), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n838), .A2(new_n829), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT123), .B1(new_n896), .B2(new_n635), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n900));
  INV_X1    g714(.A(new_n635), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n839), .A2(new_n901), .A3(new_n891), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT123), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n898), .A2(new_n899), .A3(new_n900), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n899), .A2(new_n900), .ZN(new_n905));
  NAND2_X1  g719(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n862), .B(new_n892), .C1(new_n902), .C2(KEYINPUT123), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n896), .A2(KEYINPUT123), .A3(new_n635), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n905), .B(new_n906), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n904), .A2(new_n909), .ZN(G66));
  OAI21_X1  g724(.A(G953), .B1(new_n203), .B2(new_n598), .ZN(new_n911));
  INV_X1    g725(.A(new_n805), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n828), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n913), .B2(G953), .ZN(new_n914));
  INV_X1    g728(.A(new_n306), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(G898), .B2(new_n338), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n914), .B(new_n916), .ZN(G69));
  AOI21_X1  g731(.A(new_n823), .B1(new_n313), .B2(new_n670), .ZN(new_n918));
  INV_X1    g732(.A(new_n749), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n919), .A2(new_n313), .A3(new_n662), .A4(new_n721), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n759), .A2(new_n751), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n716), .A2(new_n726), .A3(new_n723), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT126), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n338), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n338), .A2(G900), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT127), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n924), .A2(new_n929), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n570), .B1(new_n572), .B2(KEYINPUT19), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n388), .B(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n338), .B1(G227), .B2(G900), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n729), .A2(new_n460), .A3(new_n653), .A4(new_n795), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n759), .A2(new_n751), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n918), .A2(new_n665), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT62), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT125), .Z(new_n942));
  OAI211_X1 g756(.A(new_n939), .B(new_n942), .C1(KEYINPUT62), .C2(new_n940), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n934), .B1(new_n943), .B2(new_n338), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n935), .A2(new_n937), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n933), .B1(new_n928), .B2(new_n930), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n936), .B1(new_n947), .B2(new_n944), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(G72));
  NOR3_X1   g763(.A1(new_n943), .A2(new_n828), .A3(new_n912), .ZN(new_n950));
  NAND2_X1  g764(.A1(G472), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT63), .Z(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n342), .B(new_n390), .C1(new_n950), .C2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n354), .B1(new_n368), .B2(new_n390), .ZN(new_n955));
  OR3_X1    g769(.A1(new_n846), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n921), .A2(new_n923), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n913), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n952), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n390), .A2(new_n342), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n861), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n954), .A2(new_n956), .A3(new_n961), .ZN(G57));
endmodule


