

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(n638), .A2(G1996), .ZN(n616) );
  NOR2_X1 U552 ( .A1(n965), .A2(n619), .ZN(n634) );
  AND2_X1 U553 ( .A1(n600), .A2(n599), .ZN(n638) );
  XOR2_X1 U554 ( .A(n649), .B(KEYINPUT29), .Z(n666) );
  XNOR2_X1 U555 ( .A(n679), .B(KEYINPUT32), .ZN(n680) );
  INV_X1 U556 ( .A(KEYINPUT23), .ZN(n578) );
  XNOR2_X1 U557 ( .A(n579), .B(n578), .ZN(n581) );
  AND2_X1 U558 ( .A1(G2104), .A2(n530), .ZN(n527) );
  NOR2_X1 U559 ( .A1(G651), .A2(n564), .ZN(n798) );
  XOR2_X1 U560 ( .A(KEYINPUT0), .B(G543), .Z(n564) );
  INV_X1 U561 ( .A(G651), .ZN(n517) );
  NOR2_X1 U562 ( .A1(n564), .A2(n517), .ZN(n805) );
  NAND2_X1 U563 ( .A1(G75), .A2(n805), .ZN(n520) );
  NOR2_X1 U564 ( .A1(G543), .A2(n517), .ZN(n518) );
  XOR2_X1 U565 ( .A(KEYINPUT1), .B(n518), .Z(n797) );
  NAND2_X1 U566 ( .A1(G62), .A2(n797), .ZN(n519) );
  NAND2_X1 U567 ( .A1(n520), .A2(n519), .ZN(n523) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n801) );
  NAND2_X1 U569 ( .A1(n801), .A2(G88), .ZN(n521) );
  XOR2_X1 U570 ( .A(KEYINPUT86), .B(n521), .Z(n522) );
  NOR2_X1 U571 ( .A1(n523), .A2(n522), .ZN(n525) );
  NAND2_X1 U572 ( .A1(n798), .A2(G50), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(G303) );
  INV_X1 U574 ( .A(G303), .ZN(G166) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  XOR2_X1 U576 ( .A(KEYINPUT17), .B(n526), .Z(n575) );
  NAND2_X1 U577 ( .A1(G138), .A2(n575), .ZN(n529) );
  INV_X1 U578 ( .A(G2105), .ZN(n530) );
  XNOR2_X1 U579 ( .A(n527), .B(KEYINPUT66), .ZN(n708) );
  NAND2_X1 U580 ( .A1(G102), .A2(n708), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n534) );
  NOR2_X2 U582 ( .A1(G2104), .A2(n530), .ZN(n870) );
  NAND2_X1 U583 ( .A1(G126), .A2(n870), .ZN(n532) );
  AND2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n871) );
  NAND2_X1 U585 ( .A1(G114), .A2(n871), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U587 ( .A1(n534), .A2(n533), .ZN(G164) );
  NAND2_X1 U588 ( .A1(G64), .A2(n797), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G52), .A2(n798), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n541) );
  NAND2_X1 U591 ( .A1(G90), .A2(n801), .ZN(n538) );
  NAND2_X1 U592 ( .A1(G77), .A2(n805), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U594 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NOR2_X1 U595 ( .A1(n541), .A2(n540), .ZN(G171) );
  NAND2_X1 U596 ( .A1(G91), .A2(n801), .ZN(n543) );
  NAND2_X1 U597 ( .A1(G78), .A2(n805), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U599 ( .A1(G65), .A2(n797), .ZN(n545) );
  NAND2_X1 U600 ( .A1(G53), .A2(n798), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U602 ( .A(KEYINPUT70), .B(n546), .ZN(n547) );
  NOR2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U604 ( .A(n549), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U605 ( .A1(n805), .A2(G76), .ZN(n550) );
  XNOR2_X1 U606 ( .A(KEYINPUT78), .B(n550), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n801), .A2(G89), .ZN(n551) );
  XNOR2_X1 U608 ( .A(KEYINPUT4), .B(n551), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U610 ( .A(n554), .B(KEYINPUT5), .ZN(n559) );
  NAND2_X1 U611 ( .A1(G63), .A2(n797), .ZN(n556) );
  NAND2_X1 U612 ( .A1(G51), .A2(n798), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U614 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U616 ( .A(n560), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U618 ( .A1(G49), .A2(n798), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G74), .A2(G651), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U621 ( .A1(n797), .A2(n563), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n564), .A2(G87), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n566), .A2(n565), .ZN(G288) );
  NAND2_X1 U624 ( .A1(G73), .A2(n805), .ZN(n567) );
  XOR2_X1 U625 ( .A(KEYINPUT2), .B(n567), .Z(n572) );
  NAND2_X1 U626 ( .A1(G86), .A2(n801), .ZN(n569) );
  NAND2_X1 U627 ( .A1(G61), .A2(n797), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U629 ( .A(KEYINPUT85), .B(n570), .Z(n571) );
  NOR2_X1 U630 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n798), .A2(G48), .ZN(n573) );
  NAND2_X1 U632 ( .A1(n574), .A2(n573), .ZN(G305) );
  INV_X1 U633 ( .A(KEYINPUT65), .ZN(n587) );
  BUF_X1 U634 ( .A(n575), .Z(n874) );
  NAND2_X1 U635 ( .A1(G137), .A2(n874), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G113), .A2(n871), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n585) );
  NAND2_X1 U638 ( .A1(n708), .A2(G101), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n870), .A2(G125), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n581), .A2(n580), .ZN(n583) );
  INV_X1 U641 ( .A(KEYINPUT67), .ZN(n582) );
  XNOR2_X1 U642 ( .A(n583), .B(n582), .ZN(n584) );
  NOR2_X1 U643 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U644 ( .A(n587), .B(n586), .ZN(n600) );
  BUF_X1 U645 ( .A(n600), .Z(G160) );
  NAND2_X1 U646 ( .A1(G60), .A2(n797), .ZN(n589) );
  NAND2_X1 U647 ( .A1(G47), .A2(n798), .ZN(n588) );
  NAND2_X1 U648 ( .A1(n589), .A2(n588), .ZN(n594) );
  NAND2_X1 U649 ( .A1(G85), .A2(n801), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G72), .A2(n805), .ZN(n590) );
  NAND2_X1 U651 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U652 ( .A(KEYINPUT68), .B(n592), .ZN(n593) );
  NOR2_X1 U653 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U654 ( .A(n595), .B(KEYINPUT69), .ZN(G290) );
  NAND2_X1 U655 ( .A1(G8), .A2(G166), .ZN(n596) );
  NOR2_X1 U656 ( .A1(G2090), .A2(n596), .ZN(n597) );
  XNOR2_X1 U657 ( .A(n597), .B(KEYINPUT105), .ZN(n682) );
  XOR2_X1 U658 ( .A(G2078), .B(KEYINPUT25), .Z(n980) );
  NOR2_X1 U659 ( .A1(G1384), .A2(G164), .ZN(n598) );
  XNOR2_X1 U660 ( .A(n598), .B(KEYINPUT64), .ZN(n721) );
  AND2_X1 U661 ( .A1(G40), .A2(n721), .ZN(n599) );
  NAND2_X1 U662 ( .A1(n600), .A2(n599), .ZN(n669) );
  NOR2_X1 U663 ( .A1(n980), .A2(n669), .ZN(n602) );
  NOR2_X1 U664 ( .A1(n638), .A2(G1961), .ZN(n601) );
  NOR2_X1 U665 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U666 ( .A(KEYINPUT97), .B(n603), .ZN(n654) );
  NAND2_X1 U667 ( .A1(n654), .A2(G171), .ZN(n664) );
  XOR2_X1 U668 ( .A(KEYINPUT14), .B(KEYINPUT73), .Z(n605) );
  NAND2_X1 U669 ( .A1(G56), .A2(n797), .ZN(n604) );
  XNOR2_X1 U670 ( .A(n605), .B(n604), .ZN(n612) );
  XNOR2_X1 U671 ( .A(KEYINPUT74), .B(KEYINPUT13), .ZN(n610) );
  NAND2_X1 U672 ( .A1(n801), .A2(G81), .ZN(n606) );
  XNOR2_X1 U673 ( .A(n606), .B(KEYINPUT12), .ZN(n608) );
  NAND2_X1 U674 ( .A1(G68), .A2(n805), .ZN(n607) );
  NAND2_X1 U675 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U676 ( .A(n610), .B(n609), .ZN(n611) );
  NAND2_X1 U677 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U678 ( .A(n613), .B(KEYINPUT75), .ZN(n615) );
  NAND2_X1 U679 ( .A1(G43), .A2(n798), .ZN(n614) );
  NAND2_X1 U680 ( .A1(n615), .A2(n614), .ZN(n965) );
  XOR2_X1 U681 ( .A(KEYINPUT26), .B(n616), .Z(n618) );
  NAND2_X1 U682 ( .A1(n669), .A2(G1341), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U684 ( .A1(G54), .A2(n798), .ZN(n626) );
  NAND2_X1 U685 ( .A1(G79), .A2(n805), .ZN(n621) );
  NAND2_X1 U686 ( .A1(G66), .A2(n797), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U688 ( .A1(n801), .A2(G92), .ZN(n622) );
  XOR2_X1 U689 ( .A(KEYINPUT76), .B(n622), .Z(n623) );
  NOR2_X1 U690 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U691 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U692 ( .A(n627), .B(KEYINPUT15), .ZN(n949) );
  NAND2_X1 U693 ( .A1(n634), .A2(n949), .ZN(n632) );
  AND2_X1 U694 ( .A1(n638), .A2(G2067), .ZN(n628) );
  XNOR2_X1 U695 ( .A(n628), .B(KEYINPUT99), .ZN(n630) );
  NAND2_X1 U696 ( .A1(n669), .A2(G1348), .ZN(n629) );
  NAND2_X1 U697 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U698 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U699 ( .A(KEYINPUT100), .B(n633), .Z(n636) );
  NOR2_X1 U700 ( .A1(n949), .A2(n634), .ZN(n635) );
  NOR2_X1 U701 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U702 ( .A(n637), .B(KEYINPUT101), .ZN(n643) );
  NAND2_X1 U703 ( .A1(n638), .A2(G2072), .ZN(n639) );
  XNOR2_X1 U704 ( .A(n639), .B(KEYINPUT27), .ZN(n641) );
  AND2_X1 U705 ( .A1(G1956), .A2(n669), .ZN(n640) );
  NOR2_X1 U706 ( .A1(n641), .A2(n640), .ZN(n644) );
  INV_X1 U707 ( .A(G299), .ZN(n814) );
  NAND2_X1 U708 ( .A1(n644), .A2(n814), .ZN(n642) );
  NAND2_X1 U709 ( .A1(n643), .A2(n642), .ZN(n648) );
  NOR2_X1 U710 ( .A1(n644), .A2(n814), .ZN(n646) );
  XOR2_X1 U711 ( .A(KEYINPUT98), .B(KEYINPUT28), .Z(n645) );
  XNOR2_X1 U712 ( .A(n646), .B(n645), .ZN(n647) );
  NAND2_X1 U713 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U714 ( .A1(n664), .A2(n666), .ZN(n658) );
  NAND2_X1 U715 ( .A1(G8), .A2(n669), .ZN(n704) );
  NOR2_X1 U716 ( .A1(G1966), .A2(n704), .ZN(n660) );
  NOR2_X1 U717 ( .A1(G2084), .A2(n669), .ZN(n659) );
  NOR2_X1 U718 ( .A1(n660), .A2(n659), .ZN(n650) );
  NAND2_X1 U719 ( .A1(G8), .A2(n650), .ZN(n651) );
  XNOR2_X1 U720 ( .A(KEYINPUT30), .B(n651), .ZN(n652) );
  XNOR2_X1 U721 ( .A(n652), .B(KEYINPUT102), .ZN(n653) );
  NOR2_X1 U722 ( .A1(G168), .A2(n653), .ZN(n656) );
  NOR2_X1 U723 ( .A1(G171), .A2(n654), .ZN(n655) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U725 ( .A(KEYINPUT31), .B(n657), .Z(n667) );
  AND2_X1 U726 ( .A1(n658), .A2(n667), .ZN(n663) );
  AND2_X1 U727 ( .A1(G8), .A2(n659), .ZN(n661) );
  OR2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  OR2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n681) );
  AND2_X1 U730 ( .A1(n664), .A2(G286), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n677) );
  INV_X1 U732 ( .A(G286), .ZN(n668) );
  OR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n675) );
  NOR2_X1 U734 ( .A1(G1971), .A2(n704), .ZN(n671) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n669), .ZN(n670) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U737 ( .A1(n672), .A2(G303), .ZN(n673) );
  XOR2_X1 U738 ( .A(KEYINPUT103), .B(n673), .Z(n674) );
  AND2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U741 ( .A1(n678), .A2(G8), .ZN(n679) );
  NAND2_X1 U742 ( .A1(n681), .A2(n680), .ZN(n688) );
  NAND2_X1 U743 ( .A1(n682), .A2(n688), .ZN(n683) );
  NAND2_X1 U744 ( .A1(n683), .A2(n704), .ZN(n700) );
  NOR2_X1 U745 ( .A1(G1971), .A2(G303), .ZN(n685) );
  NOR2_X1 U746 ( .A1(G288), .A2(G1976), .ZN(n684) );
  XNOR2_X1 U747 ( .A(n684), .B(KEYINPUT104), .ZN(n692) );
  NOR2_X1 U748 ( .A1(n685), .A2(n692), .ZN(n946) );
  INV_X1 U749 ( .A(KEYINPUT33), .ZN(n686) );
  AND2_X1 U750 ( .A1(n946), .A2(n686), .ZN(n687) );
  NAND2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n698) );
  INV_X1 U752 ( .A(n704), .ZN(n689) );
  NAND2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n945) );
  AND2_X1 U754 ( .A1(n689), .A2(n945), .ZN(n690) );
  NOR2_X1 U755 ( .A1(KEYINPUT33), .A2(n690), .ZN(n691) );
  XNOR2_X1 U756 ( .A(G1981), .B(G305), .ZN(n961) );
  NOR2_X1 U757 ( .A1(n691), .A2(n961), .ZN(n696) );
  INV_X1 U758 ( .A(n692), .ZN(n693) );
  NOR2_X1 U759 ( .A1(n704), .A2(n693), .ZN(n694) );
  NAND2_X1 U760 ( .A1(KEYINPUT33), .A2(n694), .ZN(n695) );
  AND2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U764 ( .A(n701), .B(KEYINPUT106), .ZN(n707) );
  NOR2_X1 U765 ( .A1(G1981), .A2(G305), .ZN(n702) );
  XOR2_X1 U766 ( .A(n702), .B(KEYINPUT24), .Z(n703) );
  NOR2_X1 U767 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U768 ( .A(n705), .B(KEYINPUT96), .ZN(n706) );
  NOR2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n743) );
  NAND2_X1 U770 ( .A1(G140), .A2(n874), .ZN(n711) );
  INV_X1 U771 ( .A(n708), .ZN(n709) );
  INV_X1 U772 ( .A(n709), .ZN(n875) );
  NAND2_X1 U773 ( .A1(G104), .A2(n875), .ZN(n710) );
  NAND2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U775 ( .A(KEYINPUT34), .B(n712), .ZN(n718) );
  NAND2_X1 U776 ( .A1(G128), .A2(n870), .ZN(n714) );
  NAND2_X1 U777 ( .A1(G116), .A2(n871), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U779 ( .A(KEYINPUT35), .B(n715), .ZN(n716) );
  XNOR2_X1 U780 ( .A(KEYINPUT91), .B(n716), .ZN(n717) );
  NOR2_X1 U781 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U782 ( .A(KEYINPUT36), .B(n719), .ZN(n869) );
  XNOR2_X1 U783 ( .A(G2067), .B(KEYINPUT37), .ZN(n746) );
  NOR2_X1 U784 ( .A1(n869), .A2(n746), .ZN(n996) );
  NAND2_X1 U785 ( .A1(G160), .A2(G40), .ZN(n720) );
  NOR2_X1 U786 ( .A1(n721), .A2(n720), .ZN(n756) );
  NAND2_X1 U787 ( .A1(n996), .A2(n756), .ZN(n753) );
  NAND2_X1 U788 ( .A1(G131), .A2(n874), .ZN(n723) );
  NAND2_X1 U789 ( .A1(G119), .A2(n870), .ZN(n722) );
  NAND2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n727) );
  NAND2_X1 U791 ( .A1(n871), .A2(G107), .ZN(n725) );
  NAND2_X1 U792 ( .A1(G95), .A2(n875), .ZN(n724) );
  NAND2_X1 U793 ( .A1(n725), .A2(n724), .ZN(n726) );
  OR2_X1 U794 ( .A1(n727), .A2(n726), .ZN(n883) );
  NAND2_X1 U795 ( .A1(G1991), .A2(n883), .ZN(n728) );
  XNOR2_X1 U796 ( .A(n728), .B(KEYINPUT92), .ZN(n739) );
  XOR2_X1 U797 ( .A(KEYINPUT38), .B(KEYINPUT94), .Z(n730) );
  NAND2_X1 U798 ( .A1(G105), .A2(n875), .ZN(n729) );
  XNOR2_X1 U799 ( .A(n730), .B(n729), .ZN(n735) );
  NAND2_X1 U800 ( .A1(G129), .A2(n870), .ZN(n732) );
  NAND2_X1 U801 ( .A1(G117), .A2(n871), .ZN(n731) );
  NAND2_X1 U802 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U803 ( .A(KEYINPUT93), .B(n733), .Z(n734) );
  NOR2_X1 U804 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U805 ( .A1(n874), .A2(G141), .ZN(n736) );
  NAND2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n863) );
  NAND2_X1 U807 ( .A1(G1996), .A2(n863), .ZN(n738) );
  NAND2_X1 U808 ( .A1(n739), .A2(n738), .ZN(n1007) );
  NAND2_X1 U809 ( .A1(n1007), .A2(n756), .ZN(n740) );
  XOR2_X1 U810 ( .A(KEYINPUT95), .B(n740), .Z(n741) );
  NAND2_X1 U811 ( .A1(n753), .A2(n741), .ZN(n742) );
  NOR2_X1 U812 ( .A1(n743), .A2(n742), .ZN(n745) );
  XNOR2_X1 U813 ( .A(G1986), .B(G290), .ZN(n953) );
  NAND2_X1 U814 ( .A1(n953), .A2(n756), .ZN(n744) );
  NAND2_X1 U815 ( .A1(n745), .A2(n744), .ZN(n759) );
  NAND2_X1 U816 ( .A1(n869), .A2(n746), .ZN(n994) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n863), .ZN(n1011) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n748) );
  NOR2_X1 U819 ( .A1(G1991), .A2(n883), .ZN(n747) );
  XOR2_X1 U820 ( .A(KEYINPUT107), .B(n747), .Z(n1003) );
  NOR2_X1 U821 ( .A1(n748), .A2(n1003), .ZN(n749) );
  NOR2_X1 U822 ( .A1(n1007), .A2(n749), .ZN(n750) );
  NOR2_X1 U823 ( .A1(n1011), .A2(n750), .ZN(n751) );
  XNOR2_X1 U824 ( .A(KEYINPUT39), .B(n751), .ZN(n752) );
  XNOR2_X1 U825 ( .A(n752), .B(KEYINPUT108), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U827 ( .A1(n994), .A2(n755), .ZN(n757) );
  NAND2_X1 U828 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U829 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U830 ( .A(n760), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U831 ( .A(G2443), .B(G2446), .Z(n762) );
  XNOR2_X1 U832 ( .A(G2427), .B(G2451), .ZN(n761) );
  XNOR2_X1 U833 ( .A(n762), .B(n761), .ZN(n768) );
  XOR2_X1 U834 ( .A(G2430), .B(G2454), .Z(n764) );
  XNOR2_X1 U835 ( .A(G1341), .B(G1348), .ZN(n763) );
  XNOR2_X1 U836 ( .A(n764), .B(n763), .ZN(n766) );
  XOR2_X1 U837 ( .A(G2435), .B(G2438), .Z(n765) );
  XNOR2_X1 U838 ( .A(n766), .B(n765), .ZN(n767) );
  XOR2_X1 U839 ( .A(n768), .B(n767), .Z(n769) );
  AND2_X1 U840 ( .A1(G14), .A2(n769), .ZN(G401) );
  AND2_X1 U841 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U842 ( .A1(G123), .A2(n870), .ZN(n770) );
  XNOR2_X1 U843 ( .A(n770), .B(KEYINPUT18), .ZN(n777) );
  NAND2_X1 U844 ( .A1(G135), .A2(n874), .ZN(n772) );
  NAND2_X1 U845 ( .A1(G99), .A2(n875), .ZN(n771) );
  NAND2_X1 U846 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U847 ( .A1(G111), .A2(n871), .ZN(n773) );
  XNOR2_X1 U848 ( .A(KEYINPUT81), .B(n773), .ZN(n774) );
  NOR2_X1 U849 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U850 ( .A1(n777), .A2(n776), .ZN(n1004) );
  XNOR2_X1 U851 ( .A(G2096), .B(n1004), .ZN(n778) );
  OR2_X1 U852 ( .A1(G2100), .A2(n778), .ZN(G156) );
  INV_X1 U853 ( .A(G57), .ZN(G237) );
  INV_X1 U854 ( .A(G82), .ZN(G220) );
  NAND2_X1 U855 ( .A1(G7), .A2(G661), .ZN(n779) );
  XNOR2_X1 U856 ( .A(n779), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U857 ( .A(G223), .ZN(n838) );
  NAND2_X1 U858 ( .A1(n838), .A2(G567), .ZN(n780) );
  XOR2_X1 U859 ( .A(KEYINPUT11), .B(n780), .Z(G234) );
  INV_X1 U860 ( .A(n965), .ZN(n781) );
  NAND2_X1 U861 ( .A1(n781), .A2(G860), .ZN(G153) );
  INV_X1 U862 ( .A(G171), .ZN(G301) );
  NOR2_X1 U863 ( .A1(n949), .A2(G868), .ZN(n782) );
  XNOR2_X1 U864 ( .A(n782), .B(KEYINPUT77), .ZN(n784) );
  NAND2_X1 U865 ( .A1(G868), .A2(G301), .ZN(n783) );
  NAND2_X1 U866 ( .A1(n784), .A2(n783), .ZN(G284) );
  NAND2_X1 U867 ( .A1(G286), .A2(G868), .ZN(n786) );
  OR2_X1 U868 ( .A1(n814), .A2(G868), .ZN(n785) );
  NAND2_X1 U869 ( .A1(n786), .A2(n785), .ZN(G297) );
  INV_X1 U870 ( .A(G559), .ZN(n787) );
  NOR2_X1 U871 ( .A1(G860), .A2(n787), .ZN(n788) );
  XNOR2_X1 U872 ( .A(KEYINPUT79), .B(n788), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n789), .A2(n949), .ZN(n790) );
  XNOR2_X1 U874 ( .A(n790), .B(KEYINPUT16), .ZN(n791) );
  XNOR2_X1 U875 ( .A(KEYINPUT80), .B(n791), .ZN(G148) );
  NOR2_X1 U876 ( .A1(G868), .A2(n965), .ZN(n794) );
  NAND2_X1 U877 ( .A1(n949), .A2(G868), .ZN(n792) );
  NOR2_X1 U878 ( .A1(G559), .A2(n792), .ZN(n793) );
  NOR2_X1 U879 ( .A1(n794), .A2(n793), .ZN(G282) );
  XNOR2_X1 U880 ( .A(n965), .B(KEYINPUT82), .ZN(n796) );
  NAND2_X1 U881 ( .A1(n949), .A2(G559), .ZN(n795) );
  XNOR2_X1 U882 ( .A(n796), .B(n795), .ZN(n818) );
  NOR2_X1 U883 ( .A1(n818), .A2(G860), .ZN(n809) );
  NAND2_X1 U884 ( .A1(G67), .A2(n797), .ZN(n800) );
  NAND2_X1 U885 ( .A1(G55), .A2(n798), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G93), .A2(n801), .ZN(n802) );
  XNOR2_X1 U888 ( .A(KEYINPUT83), .B(n802), .ZN(n803) );
  NOR2_X1 U889 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U890 ( .A1(n805), .A2(G80), .ZN(n806) );
  AND2_X1 U891 ( .A1(n807), .A2(n806), .ZN(n811) );
  XNOR2_X1 U892 ( .A(n811), .B(KEYINPUT84), .ZN(n808) );
  XNOR2_X1 U893 ( .A(n809), .B(n808), .ZN(G145) );
  NOR2_X1 U894 ( .A1(G868), .A2(n811), .ZN(n810) );
  XNOR2_X1 U895 ( .A(n810), .B(KEYINPUT87), .ZN(n821) );
  XNOR2_X1 U896 ( .A(KEYINPUT19), .B(G288), .ZN(n812) );
  XOR2_X1 U897 ( .A(n812), .B(n811), .Z(n813) );
  XNOR2_X1 U898 ( .A(G290), .B(n813), .ZN(n816) );
  XNOR2_X1 U899 ( .A(n814), .B(G166), .ZN(n815) );
  XNOR2_X1 U900 ( .A(n816), .B(n815), .ZN(n817) );
  XNOR2_X1 U901 ( .A(n817), .B(G305), .ZN(n889) );
  XOR2_X1 U902 ( .A(n889), .B(n818), .Z(n819) );
  NAND2_X1 U903 ( .A1(G868), .A2(n819), .ZN(n820) );
  NAND2_X1 U904 ( .A1(n821), .A2(n820), .ZN(G295) );
  NAND2_X1 U905 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U906 ( .A(KEYINPUT20), .B(n822), .Z(n823) );
  NAND2_X1 U907 ( .A1(G2090), .A2(n823), .ZN(n824) );
  XNOR2_X1 U908 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U909 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U910 ( .A(KEYINPUT88), .B(G44), .ZN(n826) );
  XNOR2_X1 U911 ( .A(n826), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U912 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  NOR2_X1 U913 ( .A1(G219), .A2(G220), .ZN(n827) );
  XOR2_X1 U914 ( .A(KEYINPUT22), .B(n827), .Z(n828) );
  NOR2_X1 U915 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U916 ( .A1(G96), .A2(n829), .ZN(n844) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n844), .ZN(n833) );
  NAND2_X1 U918 ( .A1(G69), .A2(G120), .ZN(n830) );
  NOR2_X1 U919 ( .A1(G237), .A2(n830), .ZN(n831) );
  NAND2_X1 U920 ( .A1(G108), .A2(n831), .ZN(n845) );
  NAND2_X1 U921 ( .A1(G567), .A2(n845), .ZN(n832) );
  NAND2_X1 U922 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U923 ( .A(KEYINPUT89), .B(n834), .ZN(G319) );
  NAND2_X1 U924 ( .A1(G661), .A2(G483), .ZN(n836) );
  INV_X1 U925 ( .A(G319), .ZN(n835) );
  NOR2_X1 U926 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U927 ( .A(n837), .B(KEYINPUT90), .ZN(n843) );
  NAND2_X1 U928 ( .A1(G36), .A2(n843), .ZN(G176) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n838), .ZN(G217) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n840) );
  INV_X1 U931 ( .A(G661), .ZN(n839) );
  NOR2_X1 U932 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U933 ( .A(n841), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U935 ( .A1(n843), .A2(n842), .ZN(G188) );
  XOR2_X1 U936 ( .A(G96), .B(KEYINPUT110), .Z(G221) );
  INV_X1 U938 ( .A(G120), .ZN(G236) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n845), .A2(n844), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  NAND2_X1 U942 ( .A1(G136), .A2(n874), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n846), .B(KEYINPUT112), .ZN(n850) );
  XOR2_X1 U944 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n848) );
  NAND2_X1 U945 ( .A1(G124), .A2(n870), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  NAND2_X1 U947 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U948 ( .A1(n871), .A2(G112), .ZN(n852) );
  NAND2_X1 U949 ( .A1(G100), .A2(n875), .ZN(n851) );
  NAND2_X1 U950 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U951 ( .A1(n854), .A2(n853), .ZN(G162) );
  NAND2_X1 U952 ( .A1(G139), .A2(n874), .ZN(n856) );
  NAND2_X1 U953 ( .A1(G103), .A2(n875), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n856), .A2(n855), .ZN(n861) );
  NAND2_X1 U955 ( .A1(G127), .A2(n870), .ZN(n858) );
  NAND2_X1 U956 ( .A1(G115), .A2(n871), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U958 ( .A(KEYINPUT47), .B(n859), .Z(n860) );
  NOR2_X1 U959 ( .A1(n861), .A2(n860), .ZN(n997) );
  XOR2_X1 U960 ( .A(G162), .B(n997), .Z(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U962 ( .A(n864), .B(KEYINPUT48), .Z(n866) );
  XNOR2_X1 U963 ( .A(G164), .B(KEYINPUT46), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U965 ( .A(G160), .B(n867), .Z(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n885) );
  NAND2_X1 U967 ( .A1(G130), .A2(n870), .ZN(n873) );
  NAND2_X1 U968 ( .A1(G118), .A2(n871), .ZN(n872) );
  NAND2_X1 U969 ( .A1(n873), .A2(n872), .ZN(n880) );
  NAND2_X1 U970 ( .A1(G142), .A2(n874), .ZN(n877) );
  NAND2_X1 U971 ( .A1(G106), .A2(n875), .ZN(n876) );
  NAND2_X1 U972 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U973 ( .A(n878), .B(KEYINPUT45), .Z(n879) );
  NOR2_X1 U974 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U975 ( .A(n881), .B(n1004), .ZN(n882) );
  XNOR2_X1 U976 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U977 ( .A(n885), .B(n884), .ZN(n886) );
  NOR2_X1 U978 ( .A1(G37), .A2(n886), .ZN(G395) );
  XNOR2_X1 U979 ( .A(n965), .B(G286), .ZN(n888) );
  XNOR2_X1 U980 ( .A(G171), .B(n949), .ZN(n887) );
  XNOR2_X1 U981 ( .A(n888), .B(n887), .ZN(n890) );
  XNOR2_X1 U982 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U983 ( .A1(G37), .A2(n891), .ZN(G397) );
  XOR2_X1 U984 ( .A(G2100), .B(G2096), .Z(n893) );
  XNOR2_X1 U985 ( .A(KEYINPUT42), .B(G2678), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n893), .B(n892), .ZN(n897) );
  XOR2_X1 U987 ( .A(KEYINPUT43), .B(G2090), .Z(n895) );
  XNOR2_X1 U988 ( .A(G2072), .B(G2067), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U990 ( .A(n897), .B(n896), .Z(n899) );
  XNOR2_X1 U991 ( .A(G2078), .B(G2084), .ZN(n898) );
  XNOR2_X1 U992 ( .A(n899), .B(n898), .ZN(G227) );
  XOR2_X1 U993 ( .A(G1986), .B(G1956), .Z(n901) );
  XNOR2_X1 U994 ( .A(G1966), .B(G1961), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U996 ( .A(n902), .B(G2474), .Z(n904) );
  XNOR2_X1 U997 ( .A(G1971), .B(G1976), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U999 ( .A(KEYINPUT41), .B(G1991), .Z(n906) );
  XNOR2_X1 U1000 ( .A(G1996), .B(G1981), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(G229) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n909) );
  XOR2_X1 U1004 ( .A(KEYINPUT115), .B(n909), .Z(n916) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n912), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(KEYINPUT114), .B(n914), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1014 ( .A(G1986), .B(G24), .Z(n920) );
  XNOR2_X1 U1015 ( .A(G1971), .B(G22), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(G23), .B(G1976), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n922), .B(n921), .ZN(n935) );
  XNOR2_X1 U1021 ( .A(G1348), .B(KEYINPUT59), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(n923), .B(G4), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(G1341), .B(G19), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(G6), .B(G1981), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n930) );
  XOR2_X1 U1027 ( .A(G20), .B(G1956), .Z(n928) );
  XNOR2_X1 U1028 ( .A(KEYINPUT123), .B(n928), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1030 ( .A(KEYINPUT60), .B(n931), .Z(n933) );
  XNOR2_X1 U1031 ( .A(G1961), .B(G5), .ZN(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(G21), .B(G1966), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(KEYINPUT124), .B(n936), .ZN(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(KEYINPUT61), .B(n939), .ZN(n940) );
  XNOR2_X1 U1038 ( .A(n940), .B(KEYINPUT126), .ZN(n942) );
  INV_X1 U1039 ( .A(G16), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(G11), .A2(n943), .ZN(n1024) );
  XOR2_X1 U1042 ( .A(G16), .B(KEYINPUT56), .Z(n970) );
  INV_X1 U1043 ( .A(G1971), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(G166), .A2(n944), .ZN(n948) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(n949), .B(G1348), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(G171), .B(G1961), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1052 ( .A(G1956), .B(G299), .Z(n956) );
  XNOR2_X1 U1053 ( .A(KEYINPUT119), .B(n956), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT120), .B(n959), .ZN(n964) );
  XOR2_X1 U1056 ( .A(G168), .B(G1966), .Z(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1058 ( .A(KEYINPUT57), .B(n962), .Z(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G1341), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1062 ( .A(KEYINPUT121), .B(n968), .Z(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(KEYINPUT122), .B(n971), .ZN(n993) );
  XNOR2_X1 U1065 ( .A(G1996), .B(G32), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(G1991), .B(G25), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n979) );
  XOR2_X1 U1068 ( .A(G2072), .B(G33), .Z(n974) );
  NAND2_X1 U1069 ( .A1(n974), .A2(G28), .ZN(n977) );
  XOR2_X1 U1070 ( .A(KEYINPUT117), .B(G2067), .Z(n975) );
  XNOR2_X1 U1071 ( .A(G26), .B(n975), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(G27), .B(n980), .ZN(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1076 ( .A(KEYINPUT53), .B(n983), .Z(n986) );
  XOR2_X1 U1077 ( .A(KEYINPUT54), .B(G34), .Z(n984) );
  XNOR2_X1 U1078 ( .A(G2084), .B(n984), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(G35), .B(G2090), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1082 ( .A(KEYINPUT55), .B(n989), .Z(n990) );
  NOR2_X1 U1083 ( .A1(G29), .A2(n990), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT118), .B(n991), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n1022) );
  INV_X1 U1086 ( .A(n994), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n1009) );
  XOR2_X1 U1088 ( .A(G2072), .B(n997), .Z(n999) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1091 ( .A(n1000), .B(KEYINPUT116), .Z(n1001) );
  XNOR2_X1 U1092 ( .A(KEYINPUT50), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1016) );
  XNOR2_X1 U1097 ( .A(G160), .B(G2084), .ZN(n1014) );
  XOR2_X1 U1098 ( .A(G2090), .B(G162), .Z(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(KEYINPUT51), .B(n1012), .Z(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(KEYINPUT52), .B(n1017), .ZN(n1019) );
  INV_X1 U1104 ( .A(KEYINPUT55), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(G29), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1109 ( .A(KEYINPUT127), .B(n1025), .Z(n1026) );
  XNOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1026), .ZN(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

