//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT65), .Z(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n462), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n462), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(new_n472), .ZN(G160));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n463), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n463), .A2(new_n474), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(new_n462), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n462), .A2(G114), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n490), .A2(new_n492), .A3(KEYINPUT67), .A4(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n463), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n498), .B(new_n499), .C1(new_n468), .C2(new_n467), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n463), .B2(new_n498), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n494), .B(new_n496), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n507), .A2(new_n509), .B1(new_n506), .B2(G543), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(G543), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n513), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n514), .A2(G51), .A3(G543), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n510), .A2(new_n514), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT69), .B(G89), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n512), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n515), .A2(new_n532), .B1(new_n533), .B2(new_n518), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  AOI22_X1  g110(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n512), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n514), .A2(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G43), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n540), .B2(new_n515), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n514), .A2(G53), .A3(G543), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n514), .A2(KEYINPUT70), .A3(G53), .A4(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n549), .ZN(new_n554));
  AOI21_X1  g129(.A(KEYINPUT71), .B1(new_n554), .B2(new_n548), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT72), .B(G65), .Z(new_n557));
  AOI22_X1  g132(.A1(new_n510), .A2(new_n557), .B1(G78), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n512), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n551), .A2(KEYINPUT71), .A3(new_n552), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n526), .A2(G91), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n556), .A2(new_n559), .A3(new_n560), .A4(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  NAND2_X1  g138(.A1(new_n525), .A2(new_n528), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n538), .A2(G49), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n510), .A2(G87), .A3(new_n514), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n566), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n570), .A2(new_n567), .A3(KEYINPUT73), .A4(new_n568), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G288));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  INV_X1    g151(.A(G48), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n515), .A2(new_n576), .B1(new_n577), .B2(new_n518), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n510), .A2(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n512), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n512), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n515), .A2(new_n586), .B1(new_n587), .B2(new_n518), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n507), .A2(new_n509), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n506), .A2(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(G54), .B2(new_n538), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n510), .A2(G92), .A3(new_n514), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT74), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT74), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n510), .A2(new_n602), .A3(G92), .A4(new_n514), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n601), .B1(new_n600), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n591), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n591), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  XOR2_X1   g187(.A(G280), .B(KEYINPUT75), .Z(G297));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n480), .A2(G123), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  INV_X1    g198(.A(G111), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G2105), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(new_n478), .B2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n463), .A2(new_n470), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n628), .A2(new_n629), .A3(new_n633), .ZN(G156));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT77), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n642), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n639), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  OAI21_X1  g222(.A(G14), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(G401));
  XOR2_X1   g224(.A(G2067), .B(G2678), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT78), .ZN(new_n651));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n652), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n652), .B(KEYINPUT17), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n656), .B(new_n653), .C1(new_n651), .C2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n653), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n651), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n655), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1991), .B(G1996), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n668), .B2(new_n674), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1981), .ZN(new_n678));
  INV_X1    g253(.A(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT79), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n682), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n665), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n680), .A2(new_n682), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n682), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n686), .A2(new_n664), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(G229));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G25), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n478), .A2(G131), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n480), .A2(G119), .ZN(new_n693));
  OR2_X1    g268(.A1(G95), .A2(G2105), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n694), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(KEYINPUT80), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT80), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n692), .A2(new_n693), .A3(new_n698), .A4(new_n695), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n691), .B1(new_n701), .B2(new_n690), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT81), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(KEYINPUT81), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT35), .B(G1991), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n706), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n703), .A2(new_n708), .A3(new_n704), .ZN(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G24), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n589), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT82), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1986), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(KEYINPUT86), .B2(KEYINPUT36), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n707), .A2(new_n709), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G6), .A2(G16), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n582), .B2(G16), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT32), .B(G1981), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G16), .A2(G23), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT83), .ZN(new_n721));
  INV_X1    g296(.A(new_n569), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(new_n570), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT84), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT33), .B(G1976), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n724), .A2(G22), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G166), .B2(new_n724), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1971), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT85), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n726), .A2(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n726), .A2(new_n728), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n731), .A2(new_n732), .ZN(new_n735));
  AND4_X1   g310(.A1(new_n719), .A2(new_n733), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT34), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n715), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n741), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n715), .A2(new_n743), .A3(new_n738), .A4(new_n739), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n690), .A2(G35), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G162), .B2(new_n690), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT29), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G2090), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n724), .A2(G20), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT23), .Z(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G299), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1956), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT94), .Z(new_n754));
  OR2_X1    g329(.A1(new_n747), .A2(G2090), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n724), .A2(G21), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G168), .B2(new_n724), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT91), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1966), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n724), .A2(G5), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G171), .B2(new_n724), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n761), .A2(G1961), .ZN(new_n762));
  NOR2_X1   g337(.A1(G16), .A2(G19), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n542), .B2(G16), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT88), .B(G1341), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n690), .A2(G32), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n478), .A2(G141), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n480), .A2(G129), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT26), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n772), .A2(new_n773), .B1(G105), .B2(new_n470), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n768), .A2(new_n769), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n767), .B1(new_n775), .B2(G29), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT27), .B(G1996), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n762), .B(new_n766), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  AND3_X1   g353(.A1(new_n755), .A2(new_n759), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT24), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n690), .B1(new_n780), .B2(G34), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n780), .B2(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G160), .B2(G29), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G2084), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n786), .B1(G1961), .B2(new_n761), .C1(new_n776), .C2(new_n777), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT93), .Z(new_n788));
  NOR2_X1   g363(.A1(G4), .A2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT87), .Z(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n606), .B2(new_n724), .ZN(new_n791));
  INV_X1    g366(.A(G1348), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n690), .A2(G26), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT28), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n478), .A2(G140), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n480), .A2(G128), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n462), .A2(G116), .ZN(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n796), .B1(new_n801), .B2(G29), .ZN(new_n802));
  INV_X1    g377(.A(G2067), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT31), .B(G11), .Z(new_n805));
  NOR2_X1   g380(.A1(new_n784), .A2(new_n785), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT92), .B(G28), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT30), .ZN(new_n808));
  AOI21_X1  g383(.A(G29), .B1(new_n807), .B2(KEYINPUT30), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n805), .B(new_n806), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(G164), .A2(G29), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G27), .B2(G29), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(new_n443), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n622), .A2(G29), .A3(new_n626), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n443), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n810), .A2(new_n813), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(G29), .A2(G33), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n462), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT25), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g397(.A(G139), .B(new_n462), .C1(new_n475), .C2(new_n476), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT89), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT89), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n822), .A2(new_n826), .A3(new_n823), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n817), .B1(new_n828), .B2(new_n690), .ZN(new_n829));
  AOI211_X1 g404(.A(new_n804), .B(new_n816), .C1(new_n442), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n442), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT90), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n779), .A2(new_n794), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n754), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n742), .A2(new_n744), .A3(new_n834), .ZN(G311));
  NAND3_X1  g410(.A1(new_n742), .A2(new_n744), .A3(new_n834), .ZN(G150));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  INV_X1    g412(.A(G67), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n595), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G651), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n538), .A2(G55), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n526), .A2(G93), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n607), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n840), .A2(new_n849), .A3(new_n842), .A4(new_n841), .ZN(new_n850));
  INV_X1    g425(.A(G93), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n841), .B1(new_n851), .B2(new_n515), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n510), .A2(G67), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n512), .B1(new_n853), .B2(new_n837), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT96), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n850), .A2(new_n855), .A3(new_n542), .ZN(new_n856));
  OAI221_X1 g431(.A(KEYINPUT96), .B1(new_n852), .B2(new_n854), .C1(new_n537), .C2(new_n541), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n848), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  INV_X1    g437(.A(G860), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n861), .B2(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n845), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(G145));
  XOR2_X1   g442(.A(new_n484), .B(G160), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n627), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n801), .B(G164), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n828), .A2(KEYINPUT98), .ZN(new_n873));
  INV_X1    g448(.A(new_n775), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n828), .A2(KEYINPUT98), .A3(new_n775), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n875), .A2(new_n876), .A3(new_n700), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n700), .B1(new_n875), .B2(new_n876), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n876), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n775), .B1(new_n828), .B2(KEYINPUT98), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n701), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n875), .A2(new_n876), .A3(new_n700), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n871), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n478), .A2(G142), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n480), .A2(G130), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n462), .A2(G118), .ZN(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n885), .B(new_n886), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n631), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n879), .A2(new_n884), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n890), .B1(new_n879), .B2(new_n884), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n870), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n879), .A2(new_n884), .ZN(new_n896));
  INV_X1    g471(.A(new_n890), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n898), .A2(new_n892), .A3(new_n869), .A4(new_n891), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(KEYINPUT99), .B(G37), .Z(new_n901));
  AND3_X1   g476(.A1(new_n900), .A2(KEYINPUT40), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT40), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(G395));
  XNOR2_X1  g479(.A(new_n859), .B(new_n616), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n606), .A2(G299), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n606), .A2(G299), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n607), .A2(new_n611), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n606), .A2(G299), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(KEYINPUT41), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n905), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n907), .A2(new_n908), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n915), .B2(new_n905), .ZN(new_n916));
  NAND3_X1  g491(.A1(G305), .A2(new_n570), .A3(new_n722), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n723), .A2(new_n582), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n513), .B2(new_n519), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n513), .A2(new_n519), .A3(new_n920), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n922), .A2(new_n923), .A3(new_n589), .ZN(new_n924));
  NAND2_X1  g499(.A1(G166), .A2(KEYINPUT101), .ZN(new_n925));
  AOI21_X1  g500(.A(G290), .B1(new_n925), .B2(new_n921), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n919), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n589), .B1(new_n922), .B2(new_n923), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(G290), .A3(new_n921), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n917), .A4(new_n918), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT42), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n916), .B(new_n932), .Z(new_n933));
  MUX2_X1   g508(.A(new_n843), .B(new_n933), .S(G868), .Z(G295));
  MUX2_X1   g509(.A(new_n843), .B(new_n933), .S(G868), .Z(G331));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  NAND2_X1  g511(.A1(G168), .A2(G171), .ZN(new_n937));
  OAI21_X1  g512(.A(G286), .B1(new_n531), .B2(new_n534), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n858), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n857), .A2(new_n856), .A3(new_n937), .A4(new_n938), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n940), .A2(new_n911), .A3(new_n910), .A4(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n941), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(new_n909), .A3(new_n912), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n915), .A2(KEYINPUT104), .A3(new_n941), .A4(new_n940), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n927), .A2(new_n930), .A3(KEYINPUT105), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT105), .B1(new_n927), .B2(new_n930), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n936), .B1(new_n952), .B2(G37), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n948), .A2(new_n931), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n948), .B2(new_n951), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(KEYINPUT106), .ZN(new_n956));
  XOR2_X1   g531(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n953), .A2(new_n956), .A3(new_n960), .A4(new_n957), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n946), .A2(new_n942), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n951), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n964), .B(new_n901), .C1(new_n931), .C2(new_n948), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n962), .B1(new_n965), .B2(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n959), .A2(new_n961), .A3(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n968));
  AOI21_X1  g543(.A(new_n957), .B1(new_n953), .B2(new_n956), .ZN(new_n969));
  INV_X1    g544(.A(new_n957), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n968), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(G397));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n503), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT45), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n976), .B2(new_n975), .ZN(new_n978));
  INV_X1    g553(.A(new_n472), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n464), .A2(new_n465), .ZN(new_n980));
  OAI211_X1 g555(.A(G40), .B(new_n979), .C1(new_n980), .C2(new_n462), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1996), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(KEYINPUT46), .A3(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT124), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT46), .B1(new_n982), .B2(new_n983), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n801), .B(new_n803), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n874), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n988), .B2(new_n982), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT125), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n985), .A2(KEYINPUT47), .A3(new_n989), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n982), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n700), .A2(new_n708), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n775), .B(new_n983), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n987), .A3(new_n998), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n801), .A2(G2067), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n996), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n701), .A2(new_n706), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n987), .A2(new_n998), .ZN(new_n1003));
  OR3_X1    g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n997), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n982), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n982), .A2(new_n679), .A3(new_n589), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1007));
  XNOR2_X1  g582(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1001), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n995), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n993), .B1(new_n992), .B2(new_n994), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n526), .A2(G86), .B1(G48), .B2(new_n538), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n579), .A2(new_n580), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G651), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT113), .B(G1981), .Z(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n498), .B1(new_n467), .B2(new_n468), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT4), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1020), .A2(new_n500), .B1(new_n463), .B2(new_n495), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n1021), .B2(new_n494), .ZN(new_n1022));
  INV_X1    g597(.A(G40), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n466), .A2(new_n472), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1018), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(G1981), .B1(new_n578), .B2(new_n581), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1017), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT49), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AOI211_X1 g607(.A(KEYINPUT114), .B(KEYINPUT49), .C1(new_n1017), .C2(new_n1026), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1029), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n574), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1017), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1025), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n975), .A2(KEYINPUT50), .ZN(new_n1040));
  INV_X1    g615(.A(G2090), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n503), .A2(new_n1042), .A3(new_n974), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1024), .A4(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT45), .B1(new_n503), .B2(new_n974), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1024), .B(new_n1046), .C1(new_n1047), .C2(KEYINPUT109), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1022), .A2(new_n1049), .A3(KEYINPUT45), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT110), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1971), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n975), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1049), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n981), .B1(new_n1022), .B2(KEYINPUT45), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT110), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1047), .A2(KEYINPUT109), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1051), .A2(new_n1052), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1018), .B1(new_n1045), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G166), .A2(new_n1018), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(KEYINPUT55), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n722), .A2(G1976), .A3(new_n570), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1025), .B2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1025), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G288), .A2(new_n1036), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(new_n1029), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1039), .B1(new_n1070), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1966), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1046), .A2(new_n1024), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1047), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1040), .A2(new_n785), .A3(new_n1024), .A4(new_n1043), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(G168), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(G8), .ZN(new_n1085));
  AOI21_X1  g660(.A(G168), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT51), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(new_n1089), .A3(G8), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1087), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1088), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n981), .B1(new_n975), .B2(KEYINPUT50), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1043), .ZN(new_n1094));
  INV_X1    g669(.A(G1961), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1056), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1054), .ZN(new_n1097));
  AOI21_X1  g672(.A(G2078), .B1(new_n1051), .B2(new_n1059), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1096), .B(new_n1097), .C1(new_n1098), .C2(KEYINPUT53), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1091), .A2(new_n1092), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1078), .B1(new_n1061), .B2(new_n1069), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1060), .A2(new_n1044), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1068), .B1(new_n1103), .B2(new_n1018), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1079), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(G8), .A3(G168), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1102), .A2(new_n1104), .A3(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT115), .B(KEYINPUT63), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1109), .A2(KEYINPUT63), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1102), .B(new_n1113), .C1(new_n1069), .C2(new_n1061), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1106), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1099), .A2(G171), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT122), .B(G2078), .Z(new_n1119));
  NAND4_X1  g694(.A1(new_n978), .A2(KEYINPUT53), .A3(new_n1056), .A4(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1096), .B(new_n1120), .C1(new_n1098), .C2(KEYINPUT53), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(G171), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1117), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1102), .A2(new_n1104), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1055), .A2(new_n1058), .A3(new_n1056), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT56), .B(G2072), .Z(new_n1128));
  OR2_X1    g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT116), .B(G1956), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1094), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n1133));
  NAND2_X1  g708(.A1(G299), .A2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n1134), .B(KEYINPUT57), .Z(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1134), .B(KEYINPUT57), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1138), .A2(new_n1131), .A3(new_n1129), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1132), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(KEYINPUT61), .A3(new_n1138), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT58), .B(G1341), .Z(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n975), .B2(new_n981), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1127), .B2(G1996), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n542), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1146), .A2(KEYINPUT59), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(KEYINPUT59), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1140), .A2(new_n1142), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1024), .A2(new_n974), .A3(new_n803), .A4(new_n503), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1022), .A2(KEYINPUT118), .A3(new_n803), .A4(new_n1024), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n1155));
  AOI21_X1  g730(.A(G1348), .B1(new_n1093), .B2(new_n1043), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1094), .A2(new_n792), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT119), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT60), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1161), .A2(KEYINPUT121), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1155), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1158), .A2(KEYINPUT119), .A3(new_n1159), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n607), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1161), .A2(KEYINPUT121), .A3(new_n606), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1162), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1171), .A2(KEYINPUT60), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1149), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1141), .A2(KEYINPUT120), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1135), .B1(new_n1141), .B2(KEYINPUT120), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1171), .A2(new_n606), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1139), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1126), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1117), .B1(new_n1121), .B2(G171), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1180), .B1(G171), .B2(new_n1099), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1116), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1004), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n589), .B(G1986), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n996), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1012), .B1(new_n1184), .B2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g763(.A1(new_n900), .A2(new_n901), .ZN(new_n1190));
  INV_X1    g764(.A(G319), .ZN(new_n1191));
  OR2_X1    g765(.A1(G227), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n1193));
  OR2_X1    g767(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1195));
  AOI21_X1  g769(.A(G401), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AND3_X1   g770(.A1(new_n1196), .A2(new_n685), .A3(new_n688), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1190), .A2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n969), .A2(new_n971), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n1199), .ZN(G308));
  OAI211_X1 g774(.A(new_n1190), .B(new_n1197), .C1(new_n969), .C2(new_n971), .ZN(G225));
endmodule


