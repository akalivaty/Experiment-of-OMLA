//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G71gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G99gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT72), .Z(new_n206));
  XOR2_X1   g005(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT27), .B(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT28), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213));
  INV_X1    g012(.A(G169gat), .ZN(new_n214));
  INV_X1    g013(.A(G176gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(KEYINPUT66), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT28), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n224), .A3(new_n210), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n212), .A2(new_n222), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n227), .A2(new_n228), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n210), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(KEYINPUT24), .A3(new_n223), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n233), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT23), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n229), .A2(new_n232), .A3(new_n234), .A4(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n237), .A2(KEYINPUT64), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n237), .B2(KEYINPUT64), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n226), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G127gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G134gat), .ZN(new_n243));
  INV_X1    g042(.A(G134gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G127gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n245), .A3(KEYINPUT67), .ZN(new_n246));
  OR3_X1    g045(.A1(new_n244), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n246), .B(new_n247), .C1(KEYINPUT1), .C2(new_n248), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n243), .A2(new_n245), .ZN(new_n250));
  XOR2_X1   g049(.A(G113gat), .B(G120gat), .Z(new_n251));
  XOR2_X1   g050(.A(KEYINPUT68), .B(KEYINPUT1), .Z(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n241), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g054(.A1(G227gat), .A2(G233gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n254), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n257), .B(new_n226), .C1(new_n239), .C2(new_n240), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n208), .A2(KEYINPUT32), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263));
  INV_X1    g062(.A(new_n207), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n259), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n259), .B2(new_n264), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n205), .B1(new_n259), .B2(KEYINPUT32), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n259), .A2(new_n264), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT70), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n259), .A2(new_n263), .A3(new_n264), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n271), .A2(new_n262), .A3(new_n268), .A4(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n261), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT74), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n271), .A2(new_n268), .A3(new_n272), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n260), .B1(new_n279), .B2(new_n273), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT74), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n256), .B1(new_n255), .B2(new_n258), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT34), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(KEYINPUT73), .B2(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n283), .A2(KEYINPUT73), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n277), .A2(new_n281), .A3(new_n287), .ZN(new_n288));
  AOI211_X1 g087(.A(new_n276), .B(new_n260), .C1(new_n279), .C2(new_n273), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n286), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n288), .A2(KEYINPUT90), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT90), .B1(new_n288), .B2(new_n290), .ZN(new_n292));
  XNOR2_X1  g091(.A(G8gat), .B(G36gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT76), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(G64gat), .ZN(new_n295));
  INV_X1    g094(.A(G92gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G197gat), .ZN(new_n298));
  INV_X1    g097(.A(G204gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G197gat), .A2(G204gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT22), .ZN(new_n302));
  NAND2_X1  g101(.A1(G211gat), .A2(G218gat), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n300), .A2(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G211gat), .ZN(new_n305));
  INV_X1    g104(.A(G218gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n303), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n304), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n311));
  INV_X1    g110(.A(G226gat), .ZN(new_n312));
  INV_X1    g111(.A(G233gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n241), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n314), .B(new_n226), .C1(new_n239), .C2(new_n240), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n310), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n310), .A3(new_n317), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n297), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n297), .A3(new_n320), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT30), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(KEYINPUT30), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n321), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G141gat), .ZN(new_n329));
  INV_X1    g128(.A(G148gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT80), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G148gat), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n329), .A2(G148gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT81), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT82), .B(G155gat), .ZN(new_n341));
  INV_X1    g140(.A(G162gat), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT2), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT80), .B(G148gat), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n344), .B(new_n335), .C1(new_n345), .C2(new_n329), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n337), .A2(new_n340), .A3(new_n343), .A4(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT2), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT78), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n330), .A2(G141gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n339), .A2(new_n353), .A3(KEYINPUT2), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n338), .A2(KEYINPUT77), .A3(new_n339), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n357));
  NOR2_X1   g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n357), .B1(new_n348), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n355), .A2(new_n360), .A3(KEYINPUT79), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT79), .B1(new_n355), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n347), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n257), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n254), .B(new_n347), .C1(new_n361), .C2(new_n362), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(KEYINPUT83), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n347), .B(new_n372), .C1(new_n361), .C2(new_n362), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n254), .B1(new_n363), .B2(KEYINPUT3), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n365), .A2(KEYINPUT4), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n355), .A2(new_n360), .A3(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n347), .A4(new_n254), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n373), .A2(new_n374), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n371), .B1(new_n383), .B2(new_n367), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n375), .A2(new_n382), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n363), .A2(KEYINPUT3), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n257), .A3(new_n373), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n385), .A2(new_n387), .A3(new_n367), .A4(new_n371), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n370), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G1gat), .B(G29gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT0), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(G57gat), .ZN(new_n393));
  INV_X1    g192(.A(G85gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397));
  INV_X1    g196(.A(new_n370), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n385), .A2(new_n387), .A3(new_n367), .ZN(new_n399));
  INV_X1    g198(.A(new_n371), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n398), .B1(new_n401), .B2(new_n388), .ZN(new_n402));
  INV_X1    g201(.A(new_n395), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n396), .A2(new_n397), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(KEYINPUT6), .A3(new_n403), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n328), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT85), .B(G50gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT31), .ZN(new_n409));
  XNOR2_X1  g208(.A(G78gat), .B(G106gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n310), .B1(new_n373), .B2(new_n311), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT3), .B1(new_n310), .B2(new_n311), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n380), .B2(new_n347), .ZN(new_n414));
  OAI211_X1 g213(.A(G228gat), .B(G233gat), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n307), .A2(new_n303), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n416), .A2(KEYINPUT87), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(KEYINPUT87), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n304), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n304), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(KEYINPUT87), .A3(new_n416), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n421), .A3(new_n311), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n372), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n423), .A2(new_n363), .B1(G228gat), .B2(G233gat), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n373), .A2(new_n311), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(new_n310), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n415), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G22gat), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT86), .ZN(new_n429));
  INV_X1    g228(.A(G22gat), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n411), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(KEYINPUT88), .A3(new_n431), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n415), .A2(new_n426), .A3(new_n430), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n430), .B1(new_n415), .B2(new_n426), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT86), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n435), .B1(new_n438), .B2(KEYINPUT88), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n439), .B2(new_n411), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT35), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n407), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n291), .A2(new_n292), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT91), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n397), .B1(new_n402), .B2(new_n403), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n395), .B(new_n398), .C1(new_n401), .C2(new_n388), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n406), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n327), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n440), .B(new_n450), .C1(new_n288), .C2(new_n290), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n445), .B1(new_n451), .B2(new_n442), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n280), .A2(KEYINPUT74), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n453), .A2(new_n289), .A3(new_n286), .ZN(new_n454));
  INV_X1    g253(.A(new_n290), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n441), .B(new_n407), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(KEYINPUT91), .A3(KEYINPUT35), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n444), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT36), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n454), .B2(new_n455), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n450), .A2(new_n440), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n288), .A2(new_n290), .A3(KEYINPUT36), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n297), .ZN(new_n464));
  INV_X1    g263(.A(new_n320), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT37), .B1(new_n465), .B2(new_n318), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT37), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n319), .A2(new_n467), .A3(new_n320), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n464), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT38), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n321), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n405), .A2(new_n471), .A3(new_n406), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n469), .A2(new_n470), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n405), .A2(new_n471), .A3(KEYINPUT89), .A4(new_n406), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n385), .A2(new_n387), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n368), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(KEYINPUT39), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(new_n403), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n479), .B(KEYINPUT39), .C1(new_n368), .C2(new_n366), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT40), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n327), .A2(new_n483), .A3(new_n447), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(KEYINPUT40), .A3(new_n482), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n440), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n477), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n463), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n202), .B1(new_n458), .B2(new_n488), .ZN(new_n489));
  OR3_X1    g288(.A1(new_n291), .A2(new_n292), .A3(new_n443), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n440), .B1(new_n288), .B2(new_n290), .ZN(new_n491));
  AOI211_X1 g290(.A(new_n445), .B(new_n442), .C1(new_n491), .C2(new_n407), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT91), .B1(new_n456), .B2(KEYINPUT35), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n488), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(KEYINPUT92), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G29gat), .ZN(new_n497));
  INV_X1    g296(.A(G36gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT14), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(G29gat), .B2(G36gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G43gat), .A2(G50gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(G43gat), .A2(G50gat), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT15), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT93), .B(G50gat), .Z(new_n510));
  OAI211_X1 g309(.A(new_n509), .B(new_n505), .C1(new_n510), .C2(G43gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(G29gat), .A2(G36gat), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n512), .B(KEYINPUT95), .Z(new_n513));
  NAND4_X1  g312(.A1(new_n504), .A2(new_n508), .A3(new_n511), .A4(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n502), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(new_n508), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT17), .ZN(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT16), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(G1gat), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(G1gat), .B2(new_n518), .ZN(new_n521));
  INV_X1    g320(.A(G8gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n523), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n516), .ZN(new_n526));
  NAND2_X1  g325(.A1(G229gat), .A2(G233gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT96), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(KEYINPUT18), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n525), .B(new_n516), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n527), .B(KEYINPUT13), .Z(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n530), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(G197gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT11), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(new_n214), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT12), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n531), .A2(new_n541), .A3(new_n534), .A4(new_n535), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT97), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n544), .A2(new_n545), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G120gat), .B(G148gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(new_n215), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(new_n299), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT106), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT104), .ZN(new_n554));
  XOR2_X1   g353(.A(G99gat), .B(G106gat), .Z(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n555), .A2(KEYINPUT102), .B1(KEYINPUT8), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n394), .A2(new_n296), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n394), .A2(new_n296), .ZN(new_n559));
  NAND2_X1  g358(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT101), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT101), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(KEYINPUT100), .A3(KEYINPUT7), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n559), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n559), .B1(new_n561), .B2(new_n563), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n557), .B(new_n558), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n555), .A2(KEYINPUT102), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n564), .A2(new_n565), .ZN(new_n569));
  INV_X1    g368(.A(new_n567), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n558), .A4(new_n557), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT98), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G78gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT103), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n568), .A2(new_n577), .A3(new_n571), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n572), .A2(KEYINPUT103), .A3(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT10), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n554), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI211_X1 g385(.A(KEYINPUT104), .B(KEYINPUT10), .C1(new_n582), .C2(new_n583), .ZN(new_n587));
  INV_X1    g386(.A(new_n579), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT10), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR3_X1   g389(.A1(new_n586), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT105), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n553), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n584), .A2(new_n585), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT104), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n584), .A2(new_n554), .A3(new_n585), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n589), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n593), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(KEYINPUT106), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n584), .A2(new_n599), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n552), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n599), .ZN(new_n604));
  INV_X1    g403(.A(new_n552), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n604), .B(new_n605), .C1(new_n599), .C2(new_n584), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n489), .A2(new_n496), .A3(new_n549), .A4(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G162gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n572), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n517), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n516), .A2(new_n572), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n617), .A2(G134gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(G134gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n618), .B2(new_n619), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n612), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(new_n611), .A3(new_n622), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT21), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n577), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n242), .ZN(new_n630));
  NAND2_X1  g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n523), .B1(new_n628), .B2(new_n577), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT99), .B(G155gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n637));
  XNOR2_X1  g436(.A(G183gat), .B(G211gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n636), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n627), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n609), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n448), .A2(new_n449), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n328), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n646), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(G8gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  MUX2_X1   g449(.A(new_n648), .B(new_n650), .S(KEYINPUT42), .Z(G1325gat));
  NOR2_X1   g450(.A1(new_n291), .A2(new_n292), .ZN(new_n652));
  AOI21_X1  g451(.A(G15gat), .B1(new_n642), .B2(new_n652), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n288), .A2(KEYINPUT36), .A3(new_n290), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT36), .B1(new_n288), .B2(new_n290), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n657), .A2(G15gat), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n653), .B1(new_n642), .B2(new_n658), .ZN(G1326gat));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n440), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT43), .B(G22gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n452), .A2(new_n457), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n463), .B2(new_n487), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n477), .A2(new_n486), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n656), .A2(KEYINPUT108), .A3(new_n667), .A4(new_n461), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n664), .A2(new_n490), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n625), .A2(new_n627), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n663), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n663), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n489), .A2(new_n496), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n640), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n607), .B(KEYINPUT107), .ZN(new_n676));
  INV_X1    g475(.A(new_n549), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n672), .A2(new_n674), .A3(new_n675), .A4(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n643), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n609), .A2(new_n640), .A3(new_n671), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n497), .A3(new_n643), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(KEYINPUT45), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(KEYINPUT45), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n681), .B1(new_n684), .B2(new_n685), .ZN(G1328gat));
  NAND3_X1  g485(.A1(new_n682), .A2(new_n498), .A3(new_n328), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n687), .A2(KEYINPUT46), .ZN(new_n688));
  OAI21_X1  g487(.A(G36gat), .B1(new_n679), .B2(new_n327), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(KEYINPUT46), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(G1329gat));
  OAI21_X1  g490(.A(G43gat), .B1(new_n679), .B2(new_n656), .ZN(new_n692));
  INV_X1    g491(.A(G43gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n682), .A2(new_n693), .A3(new_n652), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT47), .Z(G1330gat));
  AND3_X1   g495(.A1(new_n489), .A2(new_n496), .A3(new_n673), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n666), .A2(new_n668), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n671), .B1(new_n698), .B2(new_n494), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n675), .B1(new_n699), .B2(KEYINPUT44), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n701), .A2(KEYINPUT110), .A3(new_n440), .A4(new_n678), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n679), .B2(new_n441), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(new_n510), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n441), .A2(new_n510), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT109), .Z(new_n707));
  NAND2_X1  g506(.A1(new_n682), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT48), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT111), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n510), .B1(new_n679), .B2(new_n441), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT48), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n713), .A3(new_n708), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n710), .A2(new_n711), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n705), .B2(new_n708), .ZN(new_n716));
  INV_X1    g515(.A(new_n714), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT111), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(G1331gat));
  INV_X1    g518(.A(new_n676), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n641), .A2(new_n549), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n669), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n643), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT112), .B(G57gat), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1332gat));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n328), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT49), .B(G64gat), .Z(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(G1333gat));
  INV_X1    g529(.A(new_n723), .ZN(new_n731));
  OAI21_X1  g530(.A(G71gat), .B1(new_n731), .B2(new_n656), .ZN(new_n732));
  INV_X1    g531(.A(G71gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n723), .A2(new_n733), .A3(new_n652), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g535(.A1(new_n723), .A2(new_n440), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g537(.A1(new_n701), .A2(new_n677), .A3(new_n607), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n680), .ZN(new_n740));
  INV_X1    g539(.A(new_n699), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n549), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n742), .A2(KEYINPUT51), .A3(new_n675), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT51), .B1(new_n742), .B2(new_n675), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(new_n394), .A3(new_n607), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n740), .B1(new_n746), .B2(new_n680), .ZN(G1336gat));
  OAI21_X1  g546(.A(G92gat), .B1(new_n739), .B2(new_n327), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n327), .A2(G92gat), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n676), .B(new_n749), .C1(new_n743), .C2(new_n744), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g551(.A(G99gat), .B1(new_n739), .B2(new_n656), .ZN(new_n753));
  INV_X1    g552(.A(G99gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n745), .A2(new_n754), .A3(new_n652), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n755), .B2(new_n608), .ZN(G1338gat));
  OAI21_X1  g555(.A(G106gat), .B1(new_n739), .B2(new_n441), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT53), .B1(new_n757), .B2(KEYINPUT113), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n441), .A2(G106gat), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n676), .B(new_n759), .C1(new_n743), .C2(new_n744), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n757), .B(new_n760), .C1(KEYINPUT113), .C2(KEYINPUT53), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(G1339gat));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n527), .B1(new_n524), .B2(new_n526), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n532), .A2(new_n533), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n540), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT115), .ZN(new_n769));
  INV_X1    g568(.A(new_n548), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(new_n546), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n607), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT54), .B1(new_n594), .B2(new_n600), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n596), .A2(new_n593), .A3(new_n589), .A4(new_n597), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n604), .A2(KEYINPUT54), .A3(new_n774), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n773), .A2(new_n775), .A3(new_n605), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n549), .B1(new_n776), .B2(KEYINPUT55), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n601), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n604), .A2(KEYINPUT54), .A3(new_n774), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n779), .A2(KEYINPUT55), .A3(new_n552), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n606), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n772), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n671), .ZN(new_n784));
  INV_X1    g583(.A(new_n782), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n779), .A2(new_n552), .A3(new_n780), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n785), .A2(new_n670), .A3(new_n771), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n640), .B1(new_n784), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n721), .A2(new_n608), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT114), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n765), .B1(new_n793), .B2(new_n440), .ZN(new_n794));
  INV_X1    g593(.A(new_n792), .ZN(new_n795));
  INV_X1    g594(.A(new_n789), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n788), .A2(new_n549), .A3(new_n606), .A4(new_n781), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n670), .B1(new_n797), .B2(new_n772), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n675), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(KEYINPUT116), .A3(new_n441), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n680), .A2(new_n328), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n794), .A2(new_n801), .A3(new_n652), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G113gat), .B1(new_n803), .B2(new_n677), .ZN(new_n804));
  INV_X1    g603(.A(new_n491), .ZN(new_n805));
  INV_X1    g604(.A(new_n802), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n793), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(G113gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n808), .A3(new_n549), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n804), .A2(new_n809), .ZN(G1340gat));
  OAI21_X1  g609(.A(G120gat), .B1(new_n803), .B2(new_n720), .ZN(new_n811));
  INV_X1    g610(.A(G120gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n807), .A2(new_n812), .A3(new_n607), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1341gat));
  NOR3_X1   g613(.A1(new_n803), .A2(new_n242), .A3(new_n675), .ZN(new_n815));
  AOI21_X1  g614(.A(G127gat), .B1(new_n807), .B2(new_n640), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(G1342gat));
  NAND2_X1  g616(.A1(new_n670), .A2(new_n327), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT117), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n800), .A2(new_n819), .A3(new_n643), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n820), .A2(G134gat), .A3(new_n805), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT56), .ZN(new_n822));
  OAI21_X1  g621(.A(G134gat), .B1(new_n803), .B2(new_n671), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1343gat));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n783), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n797), .A2(KEYINPUT118), .A3(new_n772), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(new_n671), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n640), .B1(new_n828), .B2(new_n789), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n440), .B1(new_n829), .B2(new_n792), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT57), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n793), .A2(new_n441), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n657), .A2(new_n806), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n677), .A2(new_n329), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n831), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n656), .A2(new_n440), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT119), .Z(new_n839));
  NAND3_X1  g638(.A1(new_n800), .A2(new_n802), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n329), .B1(new_n840), .B2(new_n677), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT121), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT58), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n837), .A2(new_n841), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n843), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n844), .B1(new_n845), .B2(new_n848), .ZN(G1344gat));
  OR3_X1    g648(.A1(new_n840), .A2(new_n345), .A3(new_n608), .ZN(new_n850));
  INV_X1    g649(.A(new_n791), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n833), .B(new_n440), .C1(new_n829), .C2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT57), .B1(new_n793), .B2(new_n441), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n835), .A2(new_n607), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT59), .B(G148gat), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n345), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n831), .A2(new_n834), .A3(new_n835), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n859), .B2(new_n607), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n850), .B(new_n856), .C1(new_n860), .C2(KEYINPUT59), .ZN(G1345gat));
  NOR3_X1   g660(.A1(new_n858), .A2(new_n341), .A3(new_n675), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n840), .A2(new_n675), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT122), .Z(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n864), .B2(new_n341), .ZN(G1346gat));
  OAI21_X1  g664(.A(G162gat), .B1(new_n858), .B2(new_n671), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n839), .A2(new_n342), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n820), .B2(new_n867), .ZN(G1347gat));
  NOR2_X1   g667(.A1(new_n643), .A2(new_n327), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n794), .A2(new_n801), .A3(new_n652), .A4(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G169gat), .B1(new_n870), .B2(new_n677), .ZN(new_n871));
  INV_X1    g670(.A(new_n869), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n793), .A2(new_n805), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n214), .A3(new_n549), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(G1348gat));
  NOR3_X1   g674(.A1(new_n870), .A2(new_n215), .A3(new_n720), .ZN(new_n876));
  AOI21_X1  g675(.A(G176gat), .B1(new_n873), .B2(new_n607), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(G1349gat));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n879));
  OAI21_X1  g678(.A(G183gat), .B1(new_n870), .B2(new_n675), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n873), .A2(new_n640), .A3(new_n209), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n880), .A2(new_n882), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT123), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(KEYINPUT60), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n885), .A2(new_n889), .ZN(G1350gat));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n891));
  OAI221_X1 g690(.A(G190gat), .B1(KEYINPUT124), .B2(new_n891), .C1(new_n870), .C2(new_n671), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(KEYINPUT124), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n210), .A3(new_n670), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1351gat));
  NOR2_X1   g695(.A1(new_n657), .A2(new_n872), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n832), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT125), .Z(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n298), .A3(new_n549), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n854), .A2(new_n657), .A3(new_n872), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n901), .A2(new_n549), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n298), .B2(new_n902), .ZN(G1352gat));
  XNOR2_X1  g702(.A(KEYINPUT126), .B(G204gat), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n898), .A2(new_n608), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT62), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n852), .A2(new_n853), .A3(new_n676), .A4(new_n897), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT127), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(KEYINPUT127), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n906), .A2(new_n910), .ZN(G1353gat));
  NAND3_X1  g710(.A1(new_n899), .A2(new_n305), .A3(new_n640), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n901), .A2(new_n640), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n913), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT63), .B1(new_n913), .B2(G211gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(G1354gat));
  AOI21_X1  g715(.A(G218gat), .B1(new_n899), .B2(new_n670), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n671), .A2(new_n306), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n901), .B2(new_n918), .ZN(G1355gat));
endmodule


