

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X2 U327 ( .A(KEYINPUT122), .B(n449), .ZN(n566) );
  INV_X1 U328 ( .A(G204GAT), .ZN(n296) );
  XNOR2_X1 U329 ( .A(n297), .B(n296), .ZN(n298) );
  NOR2_X1 U330 ( .A1(n415), .A2(n414), .ZN(n527) );
  XNOR2_X1 U331 ( .A(n299), .B(n298), .ZN(n332) );
  XNOR2_X1 U332 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U333 ( .A(n308), .B(n307), .ZN(n368) );
  XOR2_X1 U334 ( .A(n459), .B(KEYINPUT28), .Z(n529) );
  XNOR2_X1 U335 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U336 ( .A(n453), .B(n452), .ZN(G1349GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n301) );
  XNOR2_X1 U338 ( .A(G148GAT), .B(KEYINPUT73), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n295), .B(KEYINPUT74), .ZN(n299) );
  XNOR2_X1 U340 ( .A(G78GAT), .B(G106GAT), .ZN(n297) );
  XOR2_X1 U341 ( .A(G120GAT), .B(G57GAT), .Z(n431) );
  XNOR2_X1 U342 ( .A(n332), .B(n431), .ZN(n300) );
  XNOR2_X1 U343 ( .A(n301), .B(n300), .ZN(n308) );
  XNOR2_X1 U344 ( .A(G176GAT), .B(G92GAT), .ZN(n302) );
  XNOR2_X1 U345 ( .A(n302), .B(G64GAT), .ZN(n421) );
  XOR2_X1 U346 ( .A(n421), .B(KEYINPUT32), .Z(n304) );
  NAND2_X1 U347 ( .A1(G230GAT), .A2(G233GAT), .ZN(n303) );
  XOR2_X1 U348 ( .A(n304), .B(n303), .Z(n306) );
  XOR2_X1 U349 ( .A(G99GAT), .B(G85GAT), .Z(n371) );
  XOR2_X1 U350 ( .A(G71GAT), .B(KEYINPUT13), .Z(n395) );
  XNOR2_X1 U351 ( .A(n371), .B(n395), .ZN(n305) );
  XOR2_X1 U352 ( .A(n368), .B(KEYINPUT41), .Z(n555) );
  XOR2_X1 U353 ( .A(KEYINPUT82), .B(G176GAT), .Z(n310) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n310), .B(n309), .ZN(n329) );
  XOR2_X1 U356 ( .A(G134GAT), .B(G190GAT), .Z(n312) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G99GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U359 ( .A(KEYINPUT20), .B(G120GAT), .Z(n314) );
  XNOR2_X1 U360 ( .A(G15GAT), .B(KEYINPUT83), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U362 ( .A(n316), .B(n315), .Z(n327) );
  XNOR2_X1 U363 ( .A(KEYINPUT85), .B(KEYINPUT17), .ZN(n317) );
  XNOR2_X1 U364 ( .A(n317), .B(G183GAT), .ZN(n318) );
  XOR2_X1 U365 ( .A(n318), .B(KEYINPUT86), .Z(n320) );
  XNOR2_X1 U366 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n320), .B(n319), .ZN(n426) );
  XOR2_X1 U368 ( .A(G127GAT), .B(KEYINPUT0), .Z(n322) );
  XNOR2_X1 U369 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n321) );
  XNOR2_X1 U370 ( .A(n322), .B(n321), .ZN(n436) );
  XOR2_X1 U371 ( .A(n436), .B(G71GAT), .Z(n324) );
  NAND2_X1 U372 ( .A1(G227GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n426), .B(n325), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U376 ( .A(n329), .B(n328), .Z(n455) );
  INV_X1 U377 ( .A(n455), .ZN(n535) );
  XOR2_X1 U378 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n334) );
  XOR2_X1 U379 ( .A(G211GAT), .B(KEYINPUT21), .Z(n331) );
  XNOR2_X1 U380 ( .A(G197GAT), .B(G218GAT), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n416) );
  XNOR2_X1 U382 ( .A(n332), .B(n416), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n334), .B(n333), .ZN(n339) );
  XOR2_X1 U384 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n336) );
  XNOR2_X1 U385 ( .A(G141GAT), .B(G155GAT), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n338) );
  XOR2_X1 U387 ( .A(G162GAT), .B(KEYINPUT87), .Z(n337) );
  XNOR2_X1 U388 ( .A(n338), .B(n337), .ZN(n444) );
  XNOR2_X1 U389 ( .A(n339), .B(n444), .ZN(n347) );
  NAND2_X1 U390 ( .A1(G228GAT), .A2(G233GAT), .ZN(n345) );
  XOR2_X1 U391 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n341) );
  XNOR2_X1 U392 ( .A(G22GAT), .B(KEYINPUT89), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n343) );
  XOR2_X1 U394 ( .A(G50GAT), .B(KEYINPUT90), .Z(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U397 ( .A(n347), .B(n346), .ZN(n459) );
  XOR2_X1 U398 ( .A(KEYINPUT8), .B(KEYINPUT71), .Z(n349) );
  XNOR2_X1 U399 ( .A(G50GAT), .B(G43GAT), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U401 ( .A(KEYINPUT7), .B(n350), .ZN(n382) );
  XNOR2_X1 U402 ( .A(G15GAT), .B(G22GAT), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n351), .B(G1GAT), .ZN(n384) );
  XOR2_X1 U404 ( .A(G169GAT), .B(G8GAT), .Z(n422) );
  XOR2_X1 U405 ( .A(n384), .B(n422), .Z(n353) );
  XNOR2_X1 U406 ( .A(G36GAT), .B(G29GAT), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U408 ( .A(n382), .B(n354), .Z(n367) );
  XOR2_X1 U409 ( .A(KEYINPUT69), .B(G197GAT), .Z(n356) );
  XNOR2_X1 U410 ( .A(G113GAT), .B(G141GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U412 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n358) );
  XNOR2_X1 U413 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U415 ( .A(n360), .B(n359), .Z(n365) );
  XOR2_X1 U416 ( .A(KEYINPUT66), .B(KEYINPUT72), .Z(n362) );
  NAND2_X1 U417 ( .A1(G229GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U419 ( .A(KEYINPUT67), .B(n363), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U421 ( .A(n367), .B(n366), .Z(n504) );
  INV_X1 U422 ( .A(n504), .ZN(n574) );
  XOR2_X1 U423 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n370) );
  XNOR2_X1 U424 ( .A(KEYINPUT65), .B(KEYINPUT9), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n381) );
  XOR2_X1 U426 ( .A(G36GAT), .B(G190GAT), .Z(n419) );
  XOR2_X1 U427 ( .A(KEYINPUT75), .B(n419), .Z(n373) );
  XNOR2_X1 U428 ( .A(G218GAT), .B(n371), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U430 ( .A(G92GAT), .B(G106GAT), .Z(n375) );
  NAND2_X1 U431 ( .A1(G232GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U433 ( .A(n377), .B(n376), .Z(n379) );
  XOR2_X1 U434 ( .A(G29GAT), .B(G134GAT), .Z(n432) );
  XNOR2_X1 U435 ( .A(G162GAT), .B(n432), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n547) );
  XNOR2_X1 U439 ( .A(KEYINPUT36), .B(n547), .ZN(n585) );
  XOR2_X1 U440 ( .A(n384), .B(KEYINPUT78), .Z(n386) );
  NAND2_X1 U441 ( .A1(G231GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n402) );
  XOR2_X1 U443 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n388) );
  XNOR2_X1 U444 ( .A(G57GAT), .B(G64GAT), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U446 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n390) );
  XNOR2_X1 U447 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n400) );
  XOR2_X1 U450 ( .A(G211GAT), .B(G155GAT), .Z(n394) );
  XNOR2_X1 U451 ( .A(G183GAT), .B(G127GAT), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U453 ( .A(n396), .B(n395), .Z(n398) );
  XNOR2_X1 U454 ( .A(G8GAT), .B(G78GAT), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U457 ( .A(n402), .B(n401), .Z(n580) );
  INV_X1 U458 ( .A(n580), .ZN(n490) );
  NOR2_X1 U459 ( .A1(n585), .A2(n490), .ZN(n403) );
  XOR2_X1 U460 ( .A(KEYINPUT45), .B(n403), .Z(n404) );
  NOR2_X1 U461 ( .A1(n368), .A2(n404), .ZN(n405) );
  XOR2_X1 U462 ( .A(KEYINPUT114), .B(n405), .Z(n406) );
  NOR2_X1 U463 ( .A1(n574), .A2(n406), .ZN(n415) );
  NAND2_X1 U464 ( .A1(n574), .A2(n555), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n407), .B(KEYINPUT46), .ZN(n408) );
  NAND2_X1 U466 ( .A1(n408), .A2(n490), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n409), .B(KEYINPUT111), .ZN(n410) );
  BUF_X1 U468 ( .A(n547), .Z(n470) );
  NAND2_X1 U469 ( .A1(n410), .A2(n470), .ZN(n413) );
  XOR2_X1 U470 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n411) );
  XNOR2_X1 U471 ( .A(KEYINPUT47), .B(n411), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U473 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n526) );
  XNOR2_X1 U474 ( .A(n527), .B(n526), .ZN(n427) );
  XOR2_X1 U475 ( .A(n416), .B(G204GAT), .Z(n418) );
  NAND2_X1 U476 ( .A1(G226GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U478 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n519) );
  NOR2_X1 U482 ( .A1(n427), .A2(n519), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n428), .B(KEYINPUT54), .ZN(n446) );
  XOR2_X1 U484 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n430) );
  XNOR2_X1 U485 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n443) );
  XOR2_X1 U487 ( .A(G85GAT), .B(n431), .Z(n434) );
  XNOR2_X1 U488 ( .A(G148GAT), .B(n432), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U490 ( .A(n435), .B(KEYINPUT5), .Z(n441) );
  XOR2_X1 U491 ( .A(n436), .B(KEYINPUT1), .Z(n438) );
  NAND2_X1 U492 ( .A1(G225GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U494 ( .A(G1GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n467) );
  XNOR2_X1 U498 ( .A(KEYINPUT93), .B(n467), .ZN(n517) );
  NAND2_X1 U499 ( .A1(n446), .A2(n517), .ZN(n573) );
  NOR2_X1 U500 ( .A1(n459), .A2(n573), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n447), .B(KEYINPUT55), .ZN(n448) );
  NOR2_X1 U502 ( .A1(n535), .A2(n448), .ZN(n449) );
  NAND2_X1 U503 ( .A1(n555), .A2(n566), .ZN(n453) );
  XOR2_X1 U504 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n451) );
  XOR2_X1 U505 ( .A(G176GAT), .B(KEYINPUT56), .Z(n450) );
  XNOR2_X1 U506 ( .A(KEYINPUT27), .B(n519), .ZN(n463) );
  NOR2_X1 U507 ( .A1(n517), .A2(n463), .ZN(n528) );
  NAND2_X1 U508 ( .A1(n529), .A2(n528), .ZN(n533) );
  XNOR2_X1 U509 ( .A(KEYINPUT94), .B(n533), .ZN(n454) );
  NOR2_X1 U510 ( .A1(n455), .A2(n454), .ZN(n469) );
  NOR2_X1 U511 ( .A1(n535), .A2(n519), .ZN(n456) );
  XOR2_X1 U512 ( .A(KEYINPUT97), .B(n456), .Z(n457) );
  NOR2_X1 U513 ( .A1(n459), .A2(n457), .ZN(n458) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(n458), .Z(n465) );
  XOR2_X1 U515 ( .A(KEYINPUT96), .B(KEYINPUT26), .Z(n461) );
  NAND2_X1 U516 ( .A1(n459), .A2(n535), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U518 ( .A(KEYINPUT95), .B(n462), .ZN(n572) );
  NOR2_X1 U519 ( .A1(n463), .A2(n572), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U522 ( .A1(n469), .A2(n468), .ZN(n488) );
  NAND2_X1 U523 ( .A1(n470), .A2(n580), .ZN(n471) );
  XNOR2_X1 U524 ( .A(n471), .B(KEYINPUT80), .ZN(n472) );
  XNOR2_X1 U525 ( .A(n472), .B(KEYINPUT16), .ZN(n473) );
  NOR2_X1 U526 ( .A1(n488), .A2(n473), .ZN(n474) );
  XNOR2_X1 U527 ( .A(KEYINPUT98), .B(n474), .ZN(n505) );
  NOR2_X1 U528 ( .A1(n368), .A2(n504), .ZN(n492) );
  NAND2_X1 U529 ( .A1(n505), .A2(n492), .ZN(n475) );
  XOR2_X1 U530 ( .A(KEYINPUT99), .B(n475), .Z(n484) );
  NOR2_X1 U531 ( .A1(n517), .A2(n484), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT34), .B(n476), .Z(n477) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U534 ( .A1(n519), .A2(n484), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT100), .B(n478), .Z(n479) );
  XNOR2_X1 U536 ( .A(G8GAT), .B(n479), .ZN(G1325GAT) );
  NOR2_X1 U537 ( .A1(n484), .A2(n535), .ZN(n483) );
  XOR2_X1 U538 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n481) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n529), .A2(n484), .ZN(n486) );
  XNOR2_X1 U543 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(n487), .ZN(G1327GAT) );
  XNOR2_X1 U546 ( .A(KEYINPUT107), .B(KEYINPUT39), .ZN(n498) );
  NOR2_X1 U547 ( .A1(n585), .A2(n488), .ZN(n489) );
  NAND2_X1 U548 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n491), .B(KEYINPUT37), .ZN(n516) );
  NAND2_X1 U550 ( .A1(n516), .A2(n492), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n493), .B(KEYINPUT38), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT106), .B(n494), .ZN(n502) );
  NOR2_X1 U553 ( .A1(n517), .A2(n502), .ZN(n496) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n519), .A2(n502), .ZN(n499) );
  XOR2_X1 U558 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  NOR2_X1 U559 ( .A1(n535), .A2(n502), .ZN(n500) );
  XOR2_X1 U560 ( .A(KEYINPUT40), .B(n500), .Z(n501) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NOR2_X1 U562 ( .A1(n529), .A2(n502), .ZN(n503) );
  XOR2_X1 U563 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  AND2_X1 U564 ( .A1(n504), .A2(n555), .ZN(n515) );
  NAND2_X1 U565 ( .A1(n515), .A2(n505), .ZN(n512) );
  NOR2_X1 U566 ( .A1(n517), .A2(n512), .ZN(n507) );
  XNOR2_X1 U567 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  NOR2_X1 U570 ( .A1(n519), .A2(n512), .ZN(n509) );
  XOR2_X1 U571 ( .A(G64GAT), .B(n509), .Z(G1333GAT) );
  NOR2_X1 U572 ( .A1(n535), .A2(n512), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  NOR2_X1 U575 ( .A1(n529), .A2(n512), .ZN(n514) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n516), .A2(n515), .ZN(n523) );
  NOR2_X1 U579 ( .A1(n517), .A2(n523), .ZN(n518) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n519), .A2(n523), .ZN(n520) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n535), .A2(n523), .ZN(n521) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(n521), .Z(n522) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n522), .ZN(G1338GAT) );
  NOR2_X1 U586 ( .A1(n529), .A2(n523), .ZN(n524) );
  XOR2_X1 U587 ( .A(KEYINPUT44), .B(n524), .Z(n525) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  XOR2_X1 U589 ( .A(n527), .B(n526), .Z(n534) );
  NAND2_X1 U590 ( .A1(n528), .A2(n534), .ZN(n551) );
  NOR2_X1 U591 ( .A1(n535), .A2(n551), .ZN(n531) );
  INV_X1 U592 ( .A(n529), .ZN(n530) );
  NOR2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U594 ( .A1(KEYINPUT115), .A2(n532), .ZN(n539) );
  NOR2_X1 U595 ( .A1(KEYINPUT115), .A2(n533), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n427), .A2(n535), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n539), .A2(n538), .ZN(n548) );
  NAND2_X1 U599 ( .A1(n548), .A2(n574), .ZN(n540) );
  XNOR2_X1 U600 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U602 ( .A1(n555), .A2(n548), .ZN(n541) );
  XNOR2_X1 U603 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n546) );
  XOR2_X1 U605 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n544) );
  NAND2_X1 U606 ( .A1(n580), .A2(n548), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U608 ( .A(n546), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  INV_X1 U610 ( .A(n547), .ZN(n567) );
  NAND2_X1 U611 ( .A1(n567), .A2(n548), .ZN(n549) );
  XNOR2_X1 U612 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  XOR2_X1 U613 ( .A(G141GAT), .B(KEYINPUT119), .Z(n554) );
  NOR2_X1 U614 ( .A1(n551), .A2(n572), .ZN(n552) );
  XNOR2_X1 U615 ( .A(n552), .B(KEYINPUT118), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n574), .A2(n561), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U619 ( .A1(n555), .A2(n561), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n561), .A2(n580), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n559), .B(KEYINPUT120), .ZN(n560) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(n560), .ZN(G1346GAT) );
  XOR2_X1 U625 ( .A(G162GAT), .B(KEYINPUT121), .Z(n563) );
  NAND2_X1 U626 ( .A1(n567), .A2(n561), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n566), .A2(n574), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n580), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1351GAT) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT124), .ZN(n571) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(n571), .Z(n576) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n583) );
  NAND2_X1 U639 ( .A1(n583), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n578) );
  NAND2_X1 U642 ( .A1(n583), .A2(n368), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(G204GAT), .B(n579), .Z(G1353GAT) );
  NAND2_X1 U645 ( .A1(n583), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
  INV_X1 U648 ( .A(n583), .ZN(n584) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

