//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT74), .Z(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT66), .A2(G953), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT66), .A2(G953), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G227), .ZN(new_n194));
  XOR2_X1   g008(.A(G110), .B(G140), .Z(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT79), .ZN(new_n198));
  OR2_X1    g012(.A1(new_n198), .A2(KEYINPUT4), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(KEYINPUT4), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT78), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G104), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT77), .A3(G107), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n206), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT75), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g025(.A(KEYINPUT75), .B(KEYINPUT3), .C1(new_n206), .C2(G107), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n204), .A3(G104), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n214), .A2(new_n204), .A3(KEYINPUT76), .A4(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n202), .B1(new_n213), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n211), .A2(new_n212), .ZN(new_n221));
  INV_X1    g035(.A(new_n208), .ZN(new_n222));
  AND4_X1   g036(.A1(new_n202), .A2(new_n221), .A3(new_n219), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n201), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G143), .B(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G143), .ZN(new_n231));
  INV_X1    g045(.A(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n228), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n226), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n229), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n221), .A2(new_n219), .A3(new_n222), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT78), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n213), .A2(new_n202), .A3(new_n219), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n197), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n221), .A2(new_n219), .A3(new_n222), .A4(new_n197), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT4), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n224), .B(new_n237), .C1(new_n241), .C2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT11), .ZN(new_n245));
  INV_X1    g059(.A(G134), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(G137), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT11), .A3(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(G137), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G131), .ZN(new_n252));
  INV_X1    g066(.A(G131), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n247), .A2(new_n249), .A3(new_n253), .A4(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT1), .B1(new_n232), .B2(G146), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n232), .A2(G146), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n230), .A2(G143), .ZN(new_n259));
  OAI211_X1 g073(.A(G128), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n231), .B(new_n233), .C1(KEYINPUT1), .C2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n206), .A2(G107), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n204), .A2(G104), .ZN(new_n264));
  OAI21_X1  g078(.A(G101), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n260), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n242), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT10), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT80), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n269), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n244), .A2(new_n256), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n242), .A2(new_n266), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n260), .A2(new_n262), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n242), .B2(new_n265), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n255), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT12), .B1(new_n255), .B2(KEYINPUT81), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n255), .B(new_n278), .C1(new_n274), .C2(new_n276), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n196), .B1(new_n273), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n224), .A2(new_n237), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n239), .A2(new_n240), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n243), .B1(new_n285), .B2(G101), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n272), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n255), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n244), .A2(new_n256), .A3(new_n272), .ZN(new_n289));
  INV_X1    g103(.A(new_n196), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT82), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n283), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n283), .B2(new_n291), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n190), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G469), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n256), .B1(new_n244), .B2(new_n272), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n196), .B1(new_n273), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n280), .A2(new_n281), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n289), .A3(new_n290), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT83), .B(G469), .Z(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n190), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n189), .B1(new_n296), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n242), .A2(new_n265), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G116), .B(G119), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT2), .B(G113), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT5), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(G116), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT84), .ZN(new_n316));
  INV_X1    g130(.A(G113), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n309), .B2(KEYINPUT5), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n312), .B1(new_n319), .B2(KEYINPUT85), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT85), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n316), .A2(new_n321), .A3(new_n318), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n308), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n309), .B(new_n311), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n224), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n323), .B1(new_n326), .B2(new_n286), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT6), .ZN(new_n328));
  XNOR2_X1  g142(.A(G110), .B(G122), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT87), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT87), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n327), .A2(new_n333), .A3(new_n328), .A4(new_n330), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n328), .B1(new_n327), .B2(new_n330), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT86), .ZN(new_n337));
  OAI21_X1  g151(.A(G101), .B1(new_n220), .B2(new_n223), .ZN(new_n338));
  INV_X1    g152(.A(new_n243), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n324), .B1(new_n285), .B2(new_n201), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n320), .A2(new_n322), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n340), .A2(new_n341), .B1(new_n342), .B2(new_n308), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n337), .B1(new_n343), .B2(new_n329), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n224), .B(new_n325), .C1(new_n241), .C2(new_n243), .ZN(new_n345));
  AND4_X1   g159(.A1(new_n337), .A2(new_n345), .A3(new_n323), .A4(new_n329), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n336), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G125), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n275), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n227), .B1(new_n225), .B2(new_n228), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n234), .A2(new_n226), .A3(new_n235), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n349), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G953), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G224), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT88), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n353), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n335), .A2(new_n347), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n345), .A2(new_n323), .A3(new_n329), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(KEYINPUT86), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(KEYINPUT7), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n353), .B(new_n361), .Z(new_n362));
  INV_X1    g176(.A(new_n319), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n308), .B1(new_n312), .B2(new_n363), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n329), .B(KEYINPUT8), .Z(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n342), .B2(new_n307), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n362), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(G902), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n358), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(G210), .B1(G237), .B2(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n358), .A2(new_n368), .A3(new_n370), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n306), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G234), .ZN(new_n375));
  OAI21_X1  g189(.A(G217), .B1(new_n375), .B2(G902), .ZN(new_n376));
  XOR2_X1   g190(.A(G119), .B(G128), .Z(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT24), .B(G110), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT23), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n314), .B2(G128), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n261), .A2(KEYINPUT23), .A3(G119), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n381), .B(new_n382), .C1(G119), .C2(new_n261), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n379), .B1(new_n383), .B2(G110), .ZN(new_n384));
  INV_X1    g198(.A(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G125), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n386), .A2(KEYINPUT16), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n348), .A2(G140), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n388), .A3(KEYINPUT16), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(G146), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n388), .A3(new_n230), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n384), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT70), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n387), .A2(new_n389), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n230), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n390), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n383), .A2(G110), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n397), .B(new_n398), .C1(new_n377), .C2(new_n378), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT22), .B(G137), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n394), .A2(new_n399), .A3(new_n403), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n190), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT72), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT25), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(KEYINPUT71), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n376), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n408), .B2(new_n409), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n405), .A2(new_n190), .A3(new_n406), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n376), .A2(new_n190), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT73), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n405), .A2(new_n406), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n411), .A2(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n246), .A2(G137), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n248), .A2(G134), .ZN(new_n421));
  OAI21_X1  g235(.A(G131), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n254), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n237), .A2(new_n255), .B1(new_n275), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT30), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n352), .A2(KEYINPUT65), .B1(new_n254), .B2(new_n252), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n350), .A2(new_n351), .A3(new_n427), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n426), .A2(new_n428), .B1(new_n275), .B2(new_n423), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n425), .B(new_n325), .C1(new_n429), .C2(KEYINPUT30), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n255), .A2(new_n350), .A3(new_n351), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n275), .A2(new_n423), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n431), .A2(new_n324), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G237), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n193), .A2(G210), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT27), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT26), .B(G101), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n430), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT31), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n430), .A2(KEYINPUT31), .A3(new_n434), .A4(new_n439), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT28), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT67), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n324), .B1(new_n424), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n431), .A2(new_n446), .A3(new_n432), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT65), .B1(new_n229), .B2(new_n236), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n255), .A3(new_n428), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n324), .B1(new_n451), .B2(new_n432), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT28), .B1(new_n452), .B2(new_n433), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n439), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n444), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT32), .ZN(new_n458));
  NOR2_X1   g272(.A1(G472), .A2(G902), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n442), .A2(new_n443), .B1(new_n454), .B2(new_n455), .ZN(new_n461));
  INV_X1    g275(.A(new_n459), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT32), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT30), .B1(new_n451), .B2(new_n432), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n431), .A2(KEYINPUT30), .A3(new_n432), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n465), .A2(new_n466), .A3(new_n324), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n455), .B1(new_n467), .B2(new_n433), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT29), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n449), .A2(new_n453), .A3(new_n439), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n468), .A2(new_n470), .A3(new_n473), .A4(new_n469), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT69), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n324), .B1(new_n431), .B2(new_n432), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n475), .B(KEYINPUT28), .C1(new_n433), .C2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT28), .B1(new_n433), .B2(new_n476), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT69), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n431), .A2(new_n432), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n325), .B1(new_n480), .B2(KEYINPUT67), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n424), .A2(new_n446), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT28), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n477), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n455), .A2(new_n469), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n472), .A2(new_n474), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G472), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n419), .B1(new_n464), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g303(.A1(KEYINPUT66), .A2(G953), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT66), .A2(G953), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n490), .A2(G214), .A3(new_n435), .A4(new_n491), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n232), .A2(KEYINPUT89), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT89), .B(G143), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT18), .B(G131), .C1(new_n494), .C2(new_n496), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT89), .B(G143), .Z(new_n498));
  NAND4_X1  g312(.A1(new_n498), .A2(G214), .A3(new_n435), .A4(new_n193), .ZN(new_n499));
  NAND2_X1  g313(.A1(KEYINPUT18), .A2(G131), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n492), .A2(new_n493), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n386), .A2(new_n388), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G146), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n391), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n497), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(G113), .B(G122), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(G104), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n508), .B(KEYINPUT91), .Z(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n494), .B2(new_n496), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT17), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n499), .A2(new_n253), .A3(new_n501), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n390), .B(new_n396), .C1(new_n510), .C2(new_n511), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n506), .B(new_n509), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n386), .A2(new_n388), .A3(KEYINPUT19), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT19), .B1(new_n386), .B2(new_n388), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n230), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n519), .A2(new_n390), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n494), .A2(new_n496), .A3(G131), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n253), .B1(new_n499), .B2(new_n501), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n506), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n508), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n524), .B1(new_n523), .B2(new_n506), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n516), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(G475), .A2(G902), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(KEYINPUT92), .A3(KEYINPUT20), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n532));
  INV_X1    g346(.A(new_n529), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n500), .B1(new_n499), .B2(new_n501), .ZN(new_n535));
  INV_X1    g349(.A(new_n505), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n519), .A2(new_n390), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n510), .B2(new_n512), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT90), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n508), .A3(new_n525), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n533), .B1(new_n541), .B2(new_n516), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n532), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n531), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n397), .B1(new_n522), .B2(KEYINPUT17), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n537), .B1(new_n513), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n508), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT93), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n506), .B1(new_n514), .B2(new_n515), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n508), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n553), .A3(new_n516), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n190), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G475), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n546), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n354), .A2(G952), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n375), .B2(new_n435), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AOI211_X1 g374(.A(new_n190), .B(new_n193), .C1(G234), .C2(G237), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT21), .B(G898), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(G116), .B(G122), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(KEYINPUT96), .A3(new_n204), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT14), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G122), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(G116), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n204), .B1(new_n569), .B2(KEYINPUT14), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(G116), .ZN(new_n572));
  INV_X1    g386(.A(G116), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G122), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n574), .A3(new_n204), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n567), .A2(new_n570), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n232), .A2(G128), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n261), .A2(G143), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT95), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT95), .B1(new_n577), .B2(new_n578), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n580), .A2(new_n581), .A3(new_n246), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n577), .A2(new_n578), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(G134), .B1(new_n585), .B2(new_n579), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n565), .B(new_n576), .C1(new_n582), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n578), .A2(KEYINPUT13), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(new_n577), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n261), .A2(G143), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(KEYINPUT13), .B2(new_n578), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT13), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT94), .B1(new_n577), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n590), .B(G134), .C1(new_n592), .C2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n564), .B(new_n204), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n246), .B1(new_n580), .B2(new_n581), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n587), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n187), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(G217), .A3(new_n354), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n603));
  INV_X1    g417(.A(new_n601), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n587), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n587), .A2(KEYINPUT97), .A3(new_n598), .A4(new_n604), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n190), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(G478), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(KEYINPUT15), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n608), .B(new_n610), .Z(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n557), .A2(new_n563), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n304), .A2(new_n374), .A3(new_n489), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  OAI21_X1  g429(.A(G472), .B1(new_n461), .B2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT98), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n457), .A2(new_n459), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n619), .B(G472), .C1(new_n461), .C2(G902), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n273), .A2(new_n297), .A3(new_n196), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n290), .B1(new_n299), .B2(new_n289), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT82), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n283), .A2(new_n291), .A3(new_n292), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(G469), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n303), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n189), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n621), .A2(new_n418), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n563), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n374), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n608), .A2(G478), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n587), .A2(new_n598), .A3(new_n604), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n604), .B1(new_n587), .B2(new_n598), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT97), .ZN(new_n639));
  INV_X1    g453(.A(new_n607), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n638), .B1(KEYINPUT99), .B2(new_n605), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n599), .A2(KEYINPUT99), .A3(new_n601), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT33), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(G902), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n635), .B1(new_n646), .B2(new_n609), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT100), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n602), .B1(new_n637), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n636), .B1(new_n650), .B2(new_n643), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT33), .B1(new_n606), .B2(new_n607), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n190), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(G478), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT100), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(new_n635), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n557), .A2(new_n648), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n633), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  AOI21_X1  g475(.A(KEYINPUT102), .B1(new_n555), .B2(G475), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n663));
  INV_X1    g477(.A(G475), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n663), .B(new_n664), .C1(new_n554), .C2(new_n190), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n545), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n542), .A2(KEYINPUT101), .A3(new_n543), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n668), .A2(new_n544), .A3(new_n531), .A4(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n666), .A2(new_n612), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n633), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  NAND2_X1  g488(.A1(new_n411), .A2(new_n413), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n404), .A2(KEYINPUT36), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n400), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n416), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n618), .A2(new_n617), .A3(new_n620), .A4(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n304), .A2(new_n680), .A3(new_n374), .A4(new_n613), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n560), .B1(new_n561), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  AND4_X1   g500(.A1(new_n612), .A2(new_n666), .A3(new_n670), .A4(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n675), .A2(new_n678), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n464), .B2(new_n488), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n304), .A2(new_n687), .A3(new_n374), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XOR2_X1   g505(.A(new_n685), .B(KEYINPUT39), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n304), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n372), .A2(new_n373), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT38), .ZN(new_n697));
  INV_X1    g511(.A(new_n557), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n611), .ZN(new_n699));
  INV_X1    g513(.A(G472), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n455), .B1(new_n433), .B2(new_n476), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n440), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(G902), .B1(new_n702), .B2(KEYINPUT103), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n440), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n700), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n460), .B2(new_n463), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n305), .A2(new_n699), .A3(new_n688), .A4(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n694), .A2(new_n695), .A3(new_n697), .A4(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NAND2_X1  g527(.A1(new_n628), .A2(new_n629), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n358), .A2(new_n368), .A3(new_n370), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n370), .B1(new_n358), .B2(new_n368), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n305), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  AND4_X1   g532(.A1(new_n557), .A2(new_n648), .A3(new_n656), .A4(new_n686), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n718), .A2(KEYINPUT105), .A3(new_n689), .A4(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n304), .A2(new_n374), .A3(new_n689), .A4(new_n719), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  AOI22_X1  g539(.A1(new_n463), .A2(new_n460), .B1(new_n487), .B2(G472), .ZN(new_n726));
  AOI21_X1  g540(.A(G902), .B1(new_n298), .B2(new_n300), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n303), .B(new_n188), .C1(new_n627), .C2(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n726), .A2(new_n419), .A3(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n631), .A3(new_n374), .A4(new_n658), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT41), .B(G113), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT106), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n730), .B(new_n732), .ZN(G15));
  NAND4_X1  g547(.A1(new_n729), .A2(new_n631), .A3(new_n374), .A4(new_n671), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  INV_X1    g549(.A(new_n728), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n374), .A2(new_n689), .A3(new_n613), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT107), .B(G119), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G21));
  OAI21_X1  g553(.A(new_n444), .B1(new_n439), .B2(new_n484), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n459), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n418), .A3(new_n616), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n742), .A2(new_n728), .A3(new_n563), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n374), .A3(new_n699), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  AND3_X1   g559(.A1(new_n679), .A2(new_n616), .A3(new_n741), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n374), .A2(new_n719), .A3(new_n736), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  OAI21_X1  g562(.A(KEYINPUT108), .B1(new_n622), .B2(new_n623), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n291), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(G469), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT109), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n749), .A2(new_n754), .A3(G469), .A4(new_n751), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n627), .A2(new_n190), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n727), .B2(new_n302), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n372), .A2(new_n305), .A3(new_n373), .A4(new_n188), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(KEYINPUT42), .A3(new_n489), .A4(new_n719), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n715), .A2(new_n716), .A3(new_n306), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n758), .A3(new_n489), .A4(new_n188), .ZN(new_n765));
  INV_X1    g579(.A(new_n719), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(KEYINPUT110), .B(G131), .Z(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G33));
  INV_X1    g584(.A(new_n765), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n687), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NAND2_X1  g587(.A1(new_n624), .A2(new_n625), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n627), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n749), .A2(KEYINPUT45), .A3(new_n751), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n756), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT46), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n303), .B1(new_n778), .B2(KEYINPUT46), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n188), .B(new_n692), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n655), .B1(new_n654), .B2(new_n635), .ZN(new_n785));
  AOI211_X1 g599(.A(KEYINPUT100), .B(new_n634), .C1(new_n653), .C2(G478), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n698), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT43), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(KEYINPUT43), .A3(new_n698), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n790), .A2(KEYINPUT112), .A3(new_n791), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n621), .A2(new_n688), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT44), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n372), .A2(new_n305), .A3(new_n373), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n797), .B2(new_n798), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n784), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  NAND4_X1  g617(.A1(new_n764), .A2(new_n719), .A3(new_n726), .A4(new_n419), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n188), .ZN(new_n806));
  INV_X1    g620(.A(new_n781), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n806), .B1(new_n807), .B2(new_n779), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(KEYINPUT47), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(KEYINPUT47), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n805), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n686), .A2(new_n188), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n707), .A2(new_n679), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n374), .A3(new_n758), .A4(new_n699), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n690), .A2(new_n816), .A3(new_n747), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n724), .A2(KEYINPUT52), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(new_n724), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n762), .A2(new_n767), .B1(new_n687), .B2(new_n771), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n612), .A2(new_n546), .A3(new_n556), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(new_n657), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT113), .B1(new_n787), .B2(new_n557), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n826), .A2(new_n632), .A3(new_n630), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n614), .A2(new_n744), .A3(new_n737), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n730), .A2(new_n734), .A3(new_n681), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n719), .A2(new_n746), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n666), .A2(new_n611), .A3(new_n670), .A4(new_n686), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n714), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n464), .A2(new_n488), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n679), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n800), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n831), .A2(new_n761), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n821), .A2(new_n829), .A3(new_n830), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n813), .B1(new_n820), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n724), .A2(new_n817), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n724), .A2(new_n817), .A3(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n826), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n633), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n614), .A2(new_n744), .A3(new_n737), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n830), .A2(new_n847), .A3(new_n848), .A4(new_n837), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n768), .A2(new_n772), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n845), .A2(new_n851), .A3(KEYINPUT53), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n839), .A2(new_n840), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n840), .B1(new_n839), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n559), .B1(new_n790), .B2(new_n791), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n800), .A2(new_n728), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n489), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT48), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n857), .A2(new_n418), .A3(new_n560), .A4(new_n707), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT116), .Z(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n658), .ZN(new_n863));
  INV_X1    g677(.A(new_n742), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n856), .A2(new_n374), .A3(new_n736), .A4(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n860), .A2(new_n558), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n809), .A2(new_n810), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n727), .A2(new_n627), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n303), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n629), .B1(new_n870), .B2(KEYINPUT115), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(KEYINPUT115), .B2(new_n870), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n856), .A2(new_n864), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n800), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT114), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n736), .A2(new_n306), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n874), .A2(new_n697), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT50), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n787), .A2(new_n557), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n862), .A2(new_n881), .B1(new_n746), .B2(new_n858), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n866), .B1(new_n884), .B2(KEYINPUT51), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(KEYINPUT51), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n884), .A2(KEYINPUT117), .A3(KEYINPUT51), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n855), .B(new_n885), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(G952), .B2(G953), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n869), .A2(KEYINPUT49), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n869), .A2(KEYINPUT49), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n419), .A2(new_n306), .A3(new_n189), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OR4_X1    g709(.A1(new_n697), .A2(new_n895), .A3(new_n708), .A4(new_n788), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n891), .A2(new_n896), .ZN(G75));
  NOR2_X1   g711(.A1(new_n193), .A2(G952), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n190), .B1(new_n839), .B2(new_n852), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n900), .B2(G210), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n335), .A2(new_n347), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n357), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n899), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n901), .B2(new_n905), .ZN(G51));
  AND3_X1   g721(.A1(new_n900), .A2(new_n777), .A3(new_n776), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n756), .B(KEYINPUT57), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n820), .A2(new_n813), .A3(new_n838), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT53), .B1(new_n845), .B2(new_n851), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT54), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n839), .A2(new_n840), .A3(new_n852), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n909), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n908), .B1(new_n917), .B2(new_n301), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT119), .B1(new_n918), .B2(new_n898), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n920));
  INV_X1    g734(.A(new_n301), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT118), .B1(new_n853), .B2(new_n854), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n913), .A2(new_n910), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n921), .B1(new_n924), .B2(new_n909), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n920), .B(new_n899), .C1(new_n925), .C2(new_n908), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n919), .A2(new_n926), .ZN(G54));
  NAND2_X1  g741(.A1(KEYINPUT58), .A2(G475), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT120), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n900), .A2(new_n528), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n528), .B1(new_n900), .B2(new_n929), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n898), .ZN(G60));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT59), .Z(new_n934));
  NOR2_X1   g748(.A1(new_n855), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n641), .A2(new_n645), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n899), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n934), .B1(new_n641), .B2(new_n645), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n924), .B2(new_n938), .ZN(G63));
  INV_X1    g753(.A(KEYINPUT121), .ZN(new_n940));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT122), .Z(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n839), .B2(new_n852), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n944), .A2(new_n417), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n898), .B1(new_n944), .B2(new_n677), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n940), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT61), .Z(G66));
  INV_X1    g762(.A(G224), .ZN(new_n949));
  OAI21_X1  g763(.A(G953), .B1(new_n562), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n829), .A2(new_n830), .ZN(new_n951));
  INV_X1    g765(.A(new_n193), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(G898), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n902), .B1(new_n954), .B2(new_n952), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n953), .B(new_n955), .Z(G69));
  AND2_X1   g770(.A1(new_n811), .A2(new_n821), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n374), .A2(new_n489), .A3(new_n699), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n784), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n958), .B1(new_n784), .B2(new_n959), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n957), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n690), .A2(new_n747), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n724), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT123), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n802), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT124), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n802), .A2(new_n966), .A3(KEYINPUT124), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n465), .A2(new_n466), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n517), .A2(new_n518), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n972), .B(new_n973), .Z(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OR3_X1    g789(.A1(new_n971), .A2(new_n952), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(G227), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n952), .B1(new_n977), .B2(new_n684), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n193), .A2(G900), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n975), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n966), .A2(new_n712), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n764), .A2(new_n489), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n826), .A2(new_n693), .A3(new_n984), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n802), .A2(new_n811), .A3(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT62), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n966), .A2(new_n987), .A3(new_n712), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n983), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n981), .B1(new_n989), .B2(new_n193), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n976), .A2(KEYINPUT126), .A3(new_n979), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n979), .A2(KEYINPUT126), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n979), .A2(KEYINPUT126), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n971), .A2(new_n952), .A3(new_n975), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n993), .B(new_n994), .C1(new_n995), .C2(new_n990), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n992), .A2(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  INV_X1    g813(.A(new_n951), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n989), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n455), .B1(new_n430), .B2(new_n434), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n839), .A2(new_n852), .ZN(new_n1004));
  INV_X1    g818(.A(new_n999), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n468), .B2(new_n440), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n898), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1005), .B1(new_n971), .B2(new_n951), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n430), .A2(new_n434), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1009), .A2(new_n439), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1003), .B(new_n1007), .C1(new_n1008), .C2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(KEYINPUT127), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n969), .A2(new_n970), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n961), .A2(new_n962), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1014), .A2(new_n951), .A3(new_n1015), .A4(new_n957), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1010), .B1(new_n1017), .B2(new_n1005), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1018), .A2(new_n1019), .A3(new_n1003), .A4(new_n1007), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1013), .A2(new_n1020), .ZN(G57));
endmodule


