//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n204));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(G218gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n205), .B1(KEYINPUT22), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n204), .B1(new_n211), .B2(KEYINPUT29), .ZN(new_n212));
  AND2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(G155gat), .B2(G162gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G141gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G148gat), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G141gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G155gat), .B(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(G155gat), .ZN(new_n226));
  INV_X1    g025(.A(G162gat), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT2), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G228gat), .ZN(new_n232));
  INV_X1    g031(.A(G233gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n229), .A3(new_n204), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n211), .B1(new_n236), .B2(KEYINPUT29), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n231), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT77), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n230), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n219), .A2(new_n229), .A3(KEYINPUT77), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n212), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n234), .B1(new_n244), .B2(new_n237), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n203), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  INV_X1    g046(.A(new_n203), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(new_n238), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n246), .A2(new_n249), .B1(new_n202), .B2(G22gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(G78gat), .B(G106gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT31), .ZN(new_n252));
  INV_X1    g051(.A(G50gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(KEYINPUT80), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n239), .A2(new_n245), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(new_n239), .B2(new_n245), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n254), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT81), .B1(new_n256), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n262), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n255), .B1(new_n265), .B2(new_n260), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n266), .B(new_n267), .C1(new_n255), .C2(new_n250), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT64), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n275), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n274), .A2(KEYINPUT71), .A3(new_n276), .A4(new_n277), .ZN(new_n281));
  NOR2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n283), .A2(KEYINPUT26), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n280), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT28), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT27), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G183gat), .ZN(new_n288));
  INV_X1    g087(.A(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT27), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT68), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT68), .B1(new_n289), .B2(KEYINPUT27), .ZN(new_n292));
  INV_X1    g091(.A(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n286), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n289), .A2(KEYINPUT27), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n287), .A2(G183gat), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT69), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n288), .A2(new_n290), .A3(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n286), .A2(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n285), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT23), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(G169gat), .ZN(new_n308));
  INV_X1    g107(.A(G176gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT65), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT65), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G176gat), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n308), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n277), .B1(new_n282), .B2(KEYINPUT23), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n306), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT24), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(G183gat), .A3(G190gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(G183gat), .B(G190gat), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n316), .B(new_n318), .C1(new_n319), .C2(new_n317), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT65), .B(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n308), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n283), .A2(new_n307), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n323), .A2(KEYINPUT66), .A3(new_n277), .A4(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n315), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n327), .B(new_n277), .C1(new_n283), .C2(new_n307), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n307), .A2(G169gat), .A3(G176gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n277), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT67), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n324), .B(new_n318), .C1(new_n319), .C2(new_n317), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT25), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G113gat), .ZN(new_n336));
  INV_X1    g135(.A(G120gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(G113gat), .B2(G120gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G127gat), .B(G134gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G127gat), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n344), .A2(G134gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(G134gat), .ZN(new_n346));
  OAI22_X1  g145(.A1(new_n338), .A2(new_n340), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n305), .A2(new_n335), .A3(new_n348), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n343), .A2(new_n347), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n314), .B1(new_n322), .B2(new_n308), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n320), .B1(new_n351), .B2(KEYINPUT66), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n304), .A2(KEYINPUT24), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n289), .A2(G190gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n293), .A2(G183gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n353), .B1(new_n356), .B2(KEYINPUT24), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n357), .A2(new_n324), .A3(new_n331), .A4(new_n328), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n352), .A2(new_n315), .B1(new_n358), .B2(KEYINPUT25), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n285), .A2(new_n303), .A3(new_n304), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n350), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n272), .B1(new_n349), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT32), .ZN(new_n363));
  XOR2_X1   g162(.A(G71gat), .B(G99gat), .Z(new_n364));
  XNOR2_X1  g163(.A(G15gat), .B(G43gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n363), .B1(new_n366), .B2(KEYINPUT33), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n363), .A2(KEYINPUT33), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n371), .B2(new_n366), .ZN(new_n372));
  INV_X1    g171(.A(new_n272), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n348), .B1(new_n305), .B2(new_n335), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n350), .A3(new_n360), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n370), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n369), .B(new_n366), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n368), .B1(new_n372), .B2(new_n379), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n349), .A2(new_n361), .A3(new_n272), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n381), .A2(KEYINPUT34), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(KEYINPUT34), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n384), .B(new_n368), .C1(new_n372), .C2(new_n379), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n270), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n305), .B2(new_n335), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n359), .A2(KEYINPUT75), .A3(new_n360), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G226gat), .A2(G233gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n305), .A2(new_n335), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n394), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n211), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(G64gat), .ZN(new_n405));
  INV_X1    g204(.A(G92gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n399), .A3(new_n392), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT76), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n408), .A2(new_n409), .A3(new_n394), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n408), .B2(new_n394), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n397), .A2(new_n394), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n403), .B(new_n407), .C1(new_n413), .C2(new_n402), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n397), .A2(KEYINPUT29), .A3(new_n395), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n395), .B2(new_n393), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(new_n211), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n408), .A2(new_n394), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n412), .B1(new_n420), .B2(KEYINPUT76), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n408), .A2(new_n409), .A3(new_n394), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n419), .B1(new_n423), .B2(new_n211), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(KEYINPUT30), .A3(new_n407), .ZN(new_n425));
  XNOR2_X1  g224(.A(G1gat), .B(G29gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT0), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(G57gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n428), .B(G85gat), .Z(new_n429));
  INV_X1    g228(.A(KEYINPUT5), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n348), .B(new_n230), .ZN(new_n431));
  NAND2_X1  g230(.A1(G225gat), .A2(G233gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n243), .A2(new_n435), .A3(new_n348), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n435), .B1(new_n348), .B2(new_n230), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n204), .B1(new_n219), .B2(new_n229), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n235), .A2(new_n348), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n437), .B(new_n432), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n434), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n241), .A2(new_n350), .A3(new_n435), .A4(new_n242), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT4), .B1(new_n348), .B2(new_n230), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n430), .B(new_n432), .C1(new_n439), .C2(new_n438), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n444), .A2(KEYINPUT78), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n447));
  INV_X1    g246(.A(new_n445), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n442), .A2(new_n443), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n429), .B(new_n441), .C1(new_n446), .C2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT78), .B1(new_n444), .B2(new_n445), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n448), .A2(new_n447), .A3(new_n449), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n429), .B1(new_n456), .B2(new_n441), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  AOI211_X1 g257(.A(new_n452), .B(new_n429), .C1(new_n456), .C2(new_n441), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n407), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n402), .B1(new_n421), .B2(new_n422), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n461), .B1(new_n462), .B2(new_n419), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n416), .A2(new_n425), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT35), .B1(new_n389), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n458), .A2(new_n459), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n269), .A2(KEYINPUT35), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n416), .A2(new_n425), .A3(new_n463), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT74), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n387), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n386), .A2(new_n470), .A3(new_n387), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n467), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT38), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT37), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n407), .B1(new_n424), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n420), .A2(KEYINPUT76), .ZN(new_n479));
  INV_X1    g278(.A(new_n412), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n479), .A2(new_n402), .A3(new_n422), .A4(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n418), .A2(new_n482), .A3(new_n211), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT84), .B1(new_n401), .B2(new_n402), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT37), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n486), .B1(new_n485), .B2(KEYINPUT37), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n476), .B(new_n478), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n466), .A2(new_n414), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT37), .B1(new_n462), .B2(new_n419), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n477), .B(new_n403), .C1(new_n413), .C2(new_n402), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n461), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n490), .B1(new_n493), .B2(KEYINPUT38), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT39), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n439), .A2(new_n438), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n496), .B(new_n433), .C1(new_n444), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n429), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT83), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT83), .B1(new_n498), .B2(new_n429), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n433), .B1(new_n444), .B2(new_n497), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n504), .B(KEYINPUT39), .C1(new_n433), .C2(new_n431), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT40), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(KEYINPUT40), .B(new_n505), .C1(new_n501), .C2(new_n502), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n456), .A2(new_n441), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n429), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n269), .B1(new_n468), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT82), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n471), .A2(new_n472), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n388), .A2(KEYINPUT36), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n515), .A2(new_n516), .B1(new_n464), .B2(new_n269), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n512), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n516), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n464), .A2(new_n269), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(KEYINPUT82), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n475), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n524), .B(KEYINPUT13), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G8gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT90), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G1gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT16), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n532), .B(KEYINPUT91), .Z(new_n533));
  AOI21_X1  g332(.A(KEYINPUT92), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n528), .B(KEYINPUT90), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n531), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n527), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n527), .A3(new_n536), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G43gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n253), .ZN(new_n542));
  NAND2_X1  g341(.A1(G43gat), .A2(G50gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n545));
  OR3_X1    g344(.A1(KEYINPUT87), .A2(G29gat), .A3(G36gat), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT87), .B1(G29gat), .B2(G36gat), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n546), .A2(KEYINPUT14), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G29gat), .A2(G36gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n547), .B2(KEYINPUT14), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n545), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT88), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n542), .A2(new_n553), .A3(new_n543), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n545), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n546), .A2(KEYINPUT14), .A3(new_n547), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n547), .A2(KEYINPUT14), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n542), .A2(KEYINPUT88), .A3(new_n553), .A4(new_n543), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n556), .A2(new_n549), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n551), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT89), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n548), .A2(new_n550), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n552), .A3(new_n554), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(new_n558), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT89), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n565), .A3(new_n551), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n540), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n538), .A2(new_n561), .A3(new_n539), .A4(new_n566), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n526), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n539), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(new_n537), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n560), .A2(KEYINPUT17), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(new_n524), .A3(new_n568), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT18), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n570), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n538), .A2(new_n539), .B1(new_n561), .B2(new_n566), .ZN(new_n580));
  INV_X1    g379(.A(new_n575), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n567), .B2(new_n571), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n580), .B1(new_n582), .B2(new_n574), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n583), .A2(KEYINPUT93), .A3(KEYINPUT18), .A4(new_n524), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n576), .A2(KEYINPUT18), .A3(new_n524), .A4(new_n568), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT93), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n579), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT11), .ZN(new_n590));
  INV_X1    g389(.A(G169gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G197gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n594), .A2(KEYINPUT12), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(KEYINPUT12), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT86), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n597), .B1(new_n595), .B2(new_n596), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n588), .A2(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n595), .A2(new_n596), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n579), .A2(new_n587), .A3(new_n584), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G230gat), .A2(G233gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G71gat), .ZN(new_n608));
  INV_X1    g407(.A(G78gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G57gat), .B(G64gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT9), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n611), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G64gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(G57gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT94), .B(G57gat), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(new_n620), .B2(G64gat), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n610), .B1(KEYINPUT9), .B2(new_n612), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n616), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT95), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n616), .B(KEYINPUT95), .C1(new_n621), .C2(new_n622), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT8), .ZN(new_n628));
  NAND2_X1  g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(new_n630), .B2(new_n629), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT99), .B(G85gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n406), .ZN(new_n634));
  NAND2_X1  g433(.A1(G85gat), .A2(G92gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT7), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  OR2_X1    g436(.A1(G99gat), .A2(G106gat), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(new_n629), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n629), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n632), .A2(new_n634), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  INV_X1    g443(.A(new_n623), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(new_n641), .A3(new_n639), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n627), .ZN(new_n648));
  INV_X1    g447(.A(new_n642), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(KEYINPUT10), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n607), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n606), .B1(new_n643), .B2(new_n646), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n309), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G204gat), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n605), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n540), .B1(KEYINPUT21), .B2(new_n648), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G183gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G127gat), .B(G155gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT97), .ZN(new_n664));
  NAND2_X1  g463(.A1(G231gat), .A2(G233gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT96), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n664), .B(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n662), .A2(new_n668), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n648), .A2(KEYINPUT21), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(new_n206), .ZN(new_n674));
  OR3_X1    g473(.A1(new_n669), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n669), .B2(new_n670), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G134gat), .B(G162gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(G232gat), .A2(G233gat), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n679), .B(new_n682), .Z(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n582), .A2(new_n642), .ZN(new_n685));
  XNOR2_X1  g484(.A(G190gat), .B(G218gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT100), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(KEYINPUT101), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(KEYINPUT101), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n681), .B2(new_n680), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n567), .B2(new_n649), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n685), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n689), .B1(new_n685), .B2(new_n692), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n684), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n695), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(new_n683), .A3(new_n693), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n523), .A2(new_n660), .A3(new_n678), .A4(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n460), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n531), .ZN(G1324gat));
  NOR2_X1   g501(.A1(new_n700), .A2(new_n469), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT16), .B(G8gat), .Z(new_n704));
  AND2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n705), .A2(KEYINPUT42), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(KEYINPUT42), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n706), .B(new_n707), .C1(new_n527), .C2(new_n703), .ZN(G1325gat));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n519), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT102), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G15gat), .B1(new_n700), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n473), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(G15gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n700), .B2(new_n715), .ZN(G1326gat));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n270), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT43), .B(G22gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1327gat));
  NAND2_X1  g518(.A1(new_n521), .A2(KEYINPUT82), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n517), .A2(new_n513), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(new_n512), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n699), .B1(new_n722), .B2(new_n475), .ZN(new_n723));
  INV_X1    g522(.A(new_n660), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n678), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n726), .A2(G29gat), .A3(new_n460), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT45), .Z(new_n728));
  NAND4_X1  g527(.A1(new_n512), .A2(new_n710), .A3(new_n711), .A4(new_n520), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n475), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT103), .B1(new_n696), .B2(new_n698), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n696), .A2(new_n698), .A3(KEYINPUT103), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n730), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n723), .B2(new_n731), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n725), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n460), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n728), .A2(new_n739), .ZN(G1328gat));
  NOR3_X1   g539(.A1(new_n726), .A2(G36gat), .A3(new_n469), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT46), .ZN(new_n742));
  OAI21_X1  g541(.A(G36gat), .B1(new_n738), .B2(new_n469), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1329gat));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  INV_X1    g544(.A(new_n738), .ZN(new_n746));
  INV_X1    g545(.A(new_n712), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n541), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n473), .A2(new_n541), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n726), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n745), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G43gat), .B1(new_n738), .B2(new_n712), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n752), .B(KEYINPUT47), .C1(new_n726), .C2(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1330gat));
  OAI21_X1  g553(.A(G50gat), .B1(new_n738), .B2(new_n270), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n726), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n723), .A2(KEYINPUT104), .A3(new_n725), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n757), .A2(new_n253), .A3(new_n269), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n755), .A2(KEYINPUT48), .A3(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(G1331gat));
  NAND2_X1  g563(.A1(new_n678), .A2(new_n699), .ZN(new_n765));
  INV_X1    g564(.A(new_n659), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n765), .A2(new_n604), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n730), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n460), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(new_n620), .ZN(G1332gat));
  NOR2_X1   g569(.A1(new_n768), .A2(new_n469), .ZN(new_n771));
  NOR2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  AND2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n771), .B2(new_n772), .ZN(G1333gat));
  XNOR2_X1  g574(.A(new_n714), .B(KEYINPUT105), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n608), .B1(new_n768), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n747), .A2(G71gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n768), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g579(.A1(new_n768), .A2(new_n270), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(new_n609), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n678), .A2(new_n604), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n659), .ZN(new_n784));
  INV_X1    g583(.A(new_n699), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n523), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT44), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n784), .B1(new_n787), .B2(new_n736), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(new_n466), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n678), .A2(new_n604), .A3(new_n699), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n730), .A2(KEYINPUT51), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT51), .B1(new_n730), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n466), .A2(new_n633), .A3(new_n659), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT106), .Z(new_n795));
  OAI22_X1  g594(.A1(new_n789), .A2(new_n633), .B1(new_n793), .B2(new_n795), .ZN(G1336gat));
  OAI21_X1  g595(.A(new_n659), .B1(new_n791), .B2(new_n792), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n797), .A2(G92gat), .A3(new_n469), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(KEYINPUT52), .ZN(new_n799));
  INV_X1    g598(.A(new_n784), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n737), .A2(new_n468), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT107), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT107), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n737), .A2(new_n803), .A3(new_n468), .A4(new_n800), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(G92gat), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n406), .B1(new_n788), .B2(new_n468), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT52), .B1(new_n807), .B2(new_n798), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(G1337gat));
  NAND2_X1  g608(.A1(new_n788), .A2(new_n747), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G99gat), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n714), .A2(G99gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n797), .B2(new_n812), .ZN(G1338gat));
  NAND2_X1  g612(.A1(KEYINPUT53), .A2(G106gat), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n788), .B2(new_n269), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n270), .A2(G106gat), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n659), .B(new_n816), .C1(new_n791), .C2(new_n792), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(KEYINPUT108), .B2(KEYINPUT53), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n731), .B1(new_n523), .B2(new_n785), .ZN(new_n820));
  INV_X1    g619(.A(new_n734), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n732), .ZN(new_n822));
  AOI211_X1 g621(.A(KEYINPUT44), .B(new_n822), .C1(new_n729), .C2(new_n475), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n269), .B(new_n800), .C1(new_n820), .C2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n737), .A2(KEYINPUT109), .A3(new_n269), .A4(new_n800), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(G106gat), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n817), .A2(KEYINPUT108), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n819), .B1(new_n830), .B2(new_n831), .ZN(G1339gat));
  INV_X1    g631(.A(new_n658), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n647), .A2(new_n607), .A3(new_n650), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT110), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n647), .A2(new_n650), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n606), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT110), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n647), .A2(new_n650), .A3(new_n838), .A4(new_n607), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n835), .A2(new_n837), .A3(KEYINPUT54), .A4(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n656), .B1(new_n651), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n833), .B1(new_n845), .B2(KEYINPUT112), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n842), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT111), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT111), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n840), .A2(new_n849), .A3(KEYINPUT55), .A4(new_n842), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n843), .A2(new_n852), .A3(new_n844), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n604), .A2(new_n846), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n594), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n583), .A2(new_n524), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n568), .A2(new_n569), .A3(new_n526), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n603), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n659), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n822), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n859), .A3(new_n851), .A4(new_n853), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(new_n822), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(KEYINPUT113), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n735), .B1(new_n854), .B2(new_n860), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n863), .A2(new_n822), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n865), .A2(new_n677), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n678), .A2(new_n605), .A3(new_n766), .A4(new_n699), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n468), .A2(new_n460), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n872), .A2(new_n270), .A3(new_n473), .A4(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(new_n336), .A3(new_n605), .ZN(new_n875));
  INV_X1    g674(.A(new_n389), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n872), .A2(new_n466), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT114), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n460), .B1(new_n870), .B2(new_n871), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n880), .A3(new_n876), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n878), .A2(new_n469), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n604), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n875), .B1(new_n883), .B2(new_n336), .ZN(G1340gat));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n337), .A3(new_n659), .ZN(new_n885));
  OAI21_X1  g684(.A(G120gat), .B1(new_n874), .B2(new_n766), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(KEYINPUT115), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(KEYINPUT115), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(G1341gat));
  NAND3_X1  g688(.A1(new_n882), .A2(new_n344), .A3(new_n678), .ZN(new_n890));
  OAI21_X1  g689(.A(G127gat), .B1(new_n874), .B2(new_n677), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1342gat));
  NOR2_X1   g691(.A1(new_n699), .A2(G134gat), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n469), .A3(new_n881), .A4(new_n893), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n874), .B2(new_n699), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT116), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT117), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n894), .A2(new_n898), .A3(KEYINPUT56), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n894), .B2(KEYINPUT56), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n895), .B(new_n897), .C1(new_n899), .C2(new_n900), .ZN(G1343gat));
  NOR3_X1   g700(.A1(new_n747), .A2(new_n270), .A3(new_n468), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n605), .A2(G141gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n879), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT58), .B1(new_n904), .B2(KEYINPUT120), .ZN(new_n905));
  AOI211_X1 g704(.A(KEYINPUT57), .B(new_n270), .C1(new_n870), .C2(new_n871), .ZN(new_n906));
  XOR2_X1   g705(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n907));
  AOI21_X1  g706(.A(new_n833), .B1(new_n843), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n604), .A2(new_n851), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n785), .B1(new_n909), .B2(new_n860), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n677), .B1(new_n910), .B2(new_n868), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n270), .B1(new_n911), .B2(new_n871), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n712), .B(new_n873), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n906), .A2(new_n605), .A3(new_n914), .ZN(new_n915));
  OAI221_X1 g714(.A(new_n905), .B1(KEYINPUT120), .B2(new_n904), .C1(new_n915), .C2(new_n220), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT119), .B1(new_n906), .B2(new_n914), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n872), .A2(new_n913), .A3(new_n269), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n712), .A2(new_n873), .ZN(new_n919));
  INV_X1    g718(.A(new_n912), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(KEYINPUT57), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n917), .A2(new_n604), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n879), .A2(new_n902), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n924), .A2(G141gat), .B1(new_n926), .B2(new_n903), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT58), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n916), .B1(new_n927), .B2(new_n928), .ZN(G1344gat));
  NAND3_X1  g728(.A1(new_n917), .A2(new_n659), .A3(new_n923), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n931), .A3(G148gat), .ZN(new_n932));
  INV_X1    g731(.A(new_n910), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n863), .A2(new_n699), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n678), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n871), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n913), .B(new_n269), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n270), .B1(new_n870), .B2(new_n871), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n913), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n766), .B1(new_n919), .B2(KEYINPUT121), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n940), .B1(KEYINPUT121), .B2(new_n919), .ZN(new_n941));
  OAI21_X1  g740(.A(G148gat), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT59), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n932), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n222), .A3(new_n659), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1345gat));
  NAND3_X1  g745(.A1(new_n926), .A2(new_n226), .A3(new_n678), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n917), .A2(new_n678), .A3(new_n923), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n226), .ZN(G1346gat));
  NAND3_X1  g748(.A1(new_n917), .A2(new_n735), .A3(new_n923), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n917), .A2(new_n923), .A3(KEYINPUT122), .A4(new_n735), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(G162gat), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n926), .A2(new_n227), .A3(new_n785), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1347gat));
  NAND2_X1  g755(.A1(new_n468), .A2(new_n460), .ZN(new_n957));
  AOI211_X1 g756(.A(new_n389), .B(new_n957), .C1(new_n870), .C2(new_n871), .ZN(new_n958));
  AOI21_X1  g757(.A(G169gat), .B1(new_n958), .B2(new_n604), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n269), .B1(new_n870), .B2(new_n871), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n776), .A2(new_n957), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n605), .A2(new_n591), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1348gat));
  AOI21_X1  g763(.A(G176gat), .B1(new_n958), .B2(new_n659), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n766), .A2(new_n322), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n962), .B2(new_n966), .ZN(G1349gat));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n960), .A2(new_n678), .A3(new_n961), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(G183gat), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT123), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n678), .A2(new_n298), .A3(new_n300), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n958), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n958), .B2(new_n972), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n293), .A3(new_n735), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n785), .A3(new_n961), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(G190gat), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT125), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n978), .A2(new_n982), .A3(G190gat), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n981), .B1(new_n980), .B2(new_n983), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n977), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  NOR2_X1   g785(.A1(new_n747), .A2(new_n957), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n938), .A2(new_n987), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n988), .A2(new_n604), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n872), .A2(new_n269), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT57), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n991), .A2(new_n937), .A3(new_n987), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n604), .A2(G197gat), .ZN(new_n993));
  OAI22_X1  g792(.A1(new_n989), .A2(G197gat), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(G1352gat));
  XNOR2_X1  g794(.A(KEYINPUT126), .B(G204gat), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n766), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n988), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g797(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n996), .B1(new_n992), .B2(new_n766), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(G1353gat));
  NAND3_X1  g801(.A1(new_n988), .A2(new_n206), .A3(new_n678), .ZN(new_n1003));
  NAND4_X1  g802(.A1(new_n991), .A2(new_n678), .A3(new_n937), .A4(new_n987), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  INV_X1    g804(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1003), .B1(new_n1006), .B2(new_n1007), .ZN(G1354gat));
  NAND3_X1  g807(.A1(new_n938), .A2(new_n735), .A3(new_n987), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1009), .A2(new_n207), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n785), .A2(G218gat), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1010), .B1(new_n992), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g811(.A(new_n1012), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


