//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1173, new_n1174, new_n1175, new_n1176, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  AND3_X1   g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(new_n209));
  OR2_X1    g0009(.A1(new_n209), .A2(KEYINPUT0), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT66), .Z(new_n225));
  AOI22_X1  g0025(.A1(new_n220), .A2(KEYINPUT1), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n209), .A2(KEYINPUT0), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n210), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT68), .B(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n234), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT69), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n249), .A2(new_n250), .B1(G20), .B2(G77), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(KEYINPUT15), .B(G87), .Z(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n251), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n221), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n259), .B1(new_n261), .B2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G77), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n260), .B(new_n263), .C1(G77), .C2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G1698), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT72), .B(G107), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI22_X1  g0075(.A1(new_n273), .A2(new_n215), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n272), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n277), .A2(new_n213), .A3(G1698), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n281), .A2(new_n266), .ZN(new_n283));
  AOI211_X1 g0083(.A(new_n268), .B(new_n282), .C1(G244), .C2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n265), .B1(new_n284), .B2(G190), .ZN(new_n285));
  INV_X1    g0085(.A(G200), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(new_n284), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT71), .B(G179), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n289), .B(new_n265), .C1(G169), .C2(new_n284), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n250), .ZN(new_n292));
  INV_X1    g0092(.A(G150), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n222), .B1(new_n201), .B2(new_n203), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n212), .A2(KEYINPUT70), .ZN(new_n296));
  XOR2_X1   g0096(.A(new_n296), .B(KEYINPUT8), .Z(new_n297));
  AOI211_X1 g0097(.A(new_n294), .B(new_n295), .C1(new_n297), .C2(new_n253), .ZN(new_n298));
  INV_X1    g0098(.A(new_n259), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n264), .ZN(new_n301));
  INV_X1    g0101(.A(G50), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n262), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n302), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G1698), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n272), .A2(G222), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G223), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n309), .B1(new_n202), .B2(new_n272), .C1(new_n273), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n280), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n268), .B1(new_n283), .B2(G226), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n288), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n314), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n307), .B(new_n317), .C1(G169), .C2(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n306), .A2(KEYINPUT9), .B1(G190), .B2(new_n318), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n314), .A2(G200), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n321), .C1(KEYINPUT9), .C2(new_n306), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n322), .A2(KEYINPUT10), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(KEYINPUT10), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n291), .B(new_n319), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT18), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT76), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT16), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT7), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(G20), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT74), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT74), .A2(G33), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT3), .ZN(new_n333));
  INV_X1    g0133(.A(new_n271), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n330), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n329), .B1(new_n272), .B2(G20), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n214), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n212), .A2(new_n214), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n338), .A2(new_n203), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(G20), .B1(G159), .B2(new_n250), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n328), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT3), .B1(new_n331), .B2(new_n332), .ZN(new_n343));
  AOI21_X1  g0143(.A(G20), .B1(new_n343), .B2(new_n270), .ZN(new_n344));
  OAI21_X1  g0144(.A(G68), .B1(new_n344), .B2(new_n329), .ZN(new_n345));
  AOI211_X1 g0145(.A(KEYINPUT7), .B(G20), .C1(new_n343), .C2(new_n270), .ZN(new_n346));
  OAI211_X1 g0146(.A(KEYINPUT16), .B(new_n340), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n342), .A2(new_n347), .A3(new_n259), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n297), .A2(new_n301), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n297), .A2(new_n304), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT75), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT75), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n348), .A2(new_n354), .A3(new_n351), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n281), .A2(G232), .A3(new_n266), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n267), .B2(new_n266), .ZN(new_n358));
  MUX2_X1   g0158(.A(G223), .B(G226), .S(G1698), .Z(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(new_n343), .A3(new_n270), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n281), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n315), .ZN(new_n364));
  INV_X1    g0164(.A(G169), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n363), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n327), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n348), .A2(new_n354), .A3(new_n351), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n354), .B1(new_n348), .B2(new_n351), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n327), .B(new_n366), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n326), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n363), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT77), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n363), .A2(KEYINPUT77), .A3(new_n373), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n376), .B(new_n377), .C1(G200), .C2(new_n363), .ZN(new_n378));
  INV_X1    g0178(.A(new_n352), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT17), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT76), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(KEYINPUT18), .A3(new_n370), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n372), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n272), .A2(G226), .A3(new_n308), .ZN(new_n386));
  INV_X1    g0186(.A(G97), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n252), .B2(new_n387), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n277), .A2(new_n213), .A3(new_n308), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n280), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n268), .B1(new_n283), .B2(G238), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n394));
  OAI21_X1  g0194(.A(G169), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n393), .A2(new_n394), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n395), .A2(KEYINPUT14), .B1(new_n396), .B2(G179), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n395), .A2(KEYINPUT14), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n301), .A2(new_n214), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT12), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n253), .A2(G77), .B1(G20), .B2(new_n214), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n302), .B2(new_n292), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n401), .B(new_n404), .C1(new_n214), .C2(new_n304), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT11), .B1(new_n403), .B2(new_n259), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n399), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT73), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n396), .B2(new_n286), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n407), .B1(new_n396), .B2(G190), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT73), .B(G200), .C1(new_n393), .C2(new_n394), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n325), .A2(new_n385), .A3(new_n414), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n299), .B(new_n264), .C1(G1), .C2(new_n252), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G107), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT25), .B1(new_n301), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n301), .A2(KEYINPUT25), .A3(new_n418), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n417), .A2(G107), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n343), .A2(new_n270), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n423), .A2(KEYINPUT22), .A3(new_n222), .A4(G87), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT22), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n222), .A2(G87), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n277), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n331), .A2(new_n332), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G116), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT23), .ZN(new_n431));
  AOI21_X1  g0231(.A(G20), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n274), .A2(KEYINPUT23), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n418), .A3(G20), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(KEYINPUT83), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT83), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n432), .B2(new_n436), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n428), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n259), .B1(new_n441), .B2(KEYINPUT24), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT24), .ZN(new_n443));
  AOI211_X1 g0243(.A(new_n443), .B(new_n428), .C1(new_n440), .C2(new_n438), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n422), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT5), .B(G41), .ZN(new_n446));
  INV_X1    g0246(.A(G45), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G1), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(G274), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n280), .B1(new_n448), .B2(new_n446), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(G264), .ZN(new_n452));
  NOR2_X1   g0252(.A1(G250), .A2(G1698), .ZN(new_n453));
  INV_X1    g0253(.A(G257), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(G1698), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n423), .A2(new_n455), .B1(G294), .B2(new_n429), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n452), .B1(new_n456), .B2(new_n281), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G179), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n365), .B2(new_n457), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n445), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n343), .A2(G257), .A3(new_n308), .A4(new_n270), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n461), .A2(KEYINPUT80), .ZN(new_n462));
  AND2_X1   g0262(.A1(G264), .A2(G1698), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n423), .A2(new_n463), .B1(G303), .B2(new_n277), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(KEYINPUT80), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n280), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n450), .B1(new_n451), .B2(G270), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n417), .A2(G116), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n301), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n258), .A2(new_n221), .B1(G20), .B2(new_n471), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(new_n222), .C1(G33), .C2(new_n387), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT20), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n476), .A2(KEYINPUT81), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(KEYINPUT20), .A3(new_n475), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n476), .B2(KEYINPUT81), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n470), .B(new_n472), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT21), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n469), .A2(G169), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n468), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n466), .B2(new_n280), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G179), .A3(new_n480), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n469), .A2(G200), .ZN(new_n488));
  INV_X1    g0288(.A(new_n480), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n489), .C1(new_n373), .C2(new_n469), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n480), .A2(G169), .ZN(new_n491));
  OAI211_X1 g0291(.A(KEYINPUT82), .B(new_n481), .C1(new_n491), .C2(new_n485), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n460), .A2(new_n487), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n457), .A2(new_n286), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT84), .ZN(new_n495));
  INV_X1    g0295(.A(new_n457), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n373), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT84), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n457), .A2(new_n498), .A3(new_n286), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(new_n422), .C1(new_n444), .C2(new_n442), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n335), .A2(new_n336), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n274), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n418), .A2(KEYINPUT6), .A3(G97), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n387), .A2(new_n418), .ZN(new_n505));
  NOR2_X1   g0305(.A1(G97), .A2(G107), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n504), .B1(new_n507), .B2(KEYINPUT6), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n508), .A2(G20), .B1(G77), .B2(new_n250), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n299), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT78), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n264), .A2(G97), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n417), .B2(G97), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n514), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT78), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n451), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n454), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n423), .A2(G244), .A3(new_n308), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n272), .A2(KEYINPUT4), .A3(G244), .A4(new_n308), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n474), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n520), .B1(new_n528), .B2(new_n280), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(G190), .A3(new_n449), .ZN(new_n530));
  INV_X1    g0330(.A(new_n520), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n526), .B1(new_n522), .B2(new_n521), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n449), .B(new_n531), .C1(new_n532), .C2(new_n281), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G200), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n518), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n365), .B1(new_n529), .B2(new_n449), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n533), .A2(new_n288), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n536), .A2(new_n537), .B1(new_n510), .B2(new_n516), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n501), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n255), .A2(new_n264), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n423), .A2(new_n222), .A3(G68), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n254), .A2(new_n387), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n274), .A2(G87), .A3(G97), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n252), .A2(new_n387), .ZN(new_n544));
  AOI21_X1  g0344(.A(G20), .B1(new_n544), .B2(KEYINPUT19), .ZN(new_n545));
  OAI221_X1 g0345(.A(new_n541), .B1(KEYINPUT19), .B2(new_n542), .C1(new_n543), .C2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n540), .B1(new_n546), .B2(new_n259), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n417), .A2(new_n255), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n280), .A2(new_n448), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G250), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n448), .A2(G274), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n343), .A2(G244), .A3(G1698), .A4(new_n270), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n554), .A2(KEYINPUT79), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n423), .A2(G238), .A3(new_n308), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(KEYINPUT79), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(new_n430), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n553), .B1(new_n558), .B2(new_n280), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n288), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n549), .B(new_n560), .C1(G169), .C2(new_n559), .ZN(new_n561));
  INV_X1    g0361(.A(G87), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n416), .A2(new_n562), .ZN(new_n563));
  AOI211_X1 g0363(.A(new_n540), .B(new_n563), .C1(new_n546), .C2(new_n259), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(G190), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n286), .C2(new_n559), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n493), .A2(new_n539), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n415), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g0369(.A(new_n569), .B(KEYINPUT85), .Z(G372));
  INV_X1    g0370(.A(KEYINPUT87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n460), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n492), .A2(new_n483), .A3(new_n486), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT86), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT86), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n492), .A2(new_n483), .A3(new_n575), .A4(new_n486), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n445), .A2(KEYINPUT87), .A3(new_n459), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n572), .A2(new_n574), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n539), .A2(new_n567), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n567), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT26), .ZN(new_n582));
  INV_X1    g0382(.A(new_n537), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n533), .A2(G169), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n518), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n581), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n584), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n511), .A2(new_n514), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n587), .A2(new_n566), .A3(new_n561), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT26), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n561), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n415), .B1(new_n580), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n319), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n352), .A2(new_n366), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n594), .B(new_n326), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n408), .A2(new_n290), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n381), .A2(new_n413), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n323), .A2(new_n324), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n593), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n592), .A2(new_n600), .ZN(G369));
  INV_X1    g0401(.A(G13), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(G20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n261), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n604), .B(KEYINPUT88), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT27), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n606), .B(KEYINPUT89), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n605), .A2(KEYINPUT27), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n608), .A2(G213), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(G343), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n480), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n573), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n574), .A2(new_n576), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n490), .B(new_n614), .C1(new_n615), .C2(new_n613), .ZN(new_n616));
  INV_X1    g0416(.A(G330), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n445), .A2(new_n612), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n460), .A2(new_n619), .A3(new_n501), .ZN(new_n620));
  INV_X1    g0420(.A(new_n612), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n460), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n573), .A2(new_n621), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n612), .B1(new_n572), .B2(new_n577), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n627), .ZN(G399));
  INV_X1    g0428(.A(new_n207), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(G41), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G1), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n543), .A2(new_n471), .ZN(new_n633));
  INV_X1    g0433(.A(new_n225), .ZN(new_n634));
  OAI22_X1  g0434(.A1(new_n632), .A2(new_n633), .B1(new_n634), .B2(new_n631), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n635), .B(KEYINPUT28), .ZN(new_n636));
  INV_X1    g0436(.A(new_n585), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT26), .B1(new_n637), .B2(new_n567), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n638), .B(new_n561), .C1(KEYINPUT26), .C2(new_n589), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n573), .B1(new_n445), .B2(new_n459), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n640), .A2(new_n539), .A3(new_n567), .ZN(new_n641));
  OAI211_X1 g0441(.A(KEYINPUT29), .B(new_n621), .C1(new_n639), .C2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n580), .A2(new_n591), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(new_n612), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n644), .B2(KEYINPUT29), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n529), .A2(new_n559), .A3(new_n496), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(KEYINPUT30), .A3(G179), .A4(new_n485), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT30), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n529), .A2(new_n559), .A3(new_n496), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n485), .A2(G179), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n533), .A2(new_n457), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n558), .A2(new_n280), .ZN(new_n654));
  INV_X1    g0454(.A(new_n553), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n469), .A3(new_n288), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT90), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n656), .A2(new_n469), .A3(KEYINPUT90), .A4(new_n288), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n653), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(KEYINPUT31), .B(new_n612), .C1(new_n652), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT91), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n612), .B1(new_n652), .B2(new_n661), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT31), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(KEYINPUT91), .A3(new_n665), .ZN(new_n668));
  INV_X1    g0468(.A(new_n493), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n579), .A2(new_n669), .A3(new_n621), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n645), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n636), .B1(new_n674), .B2(G1), .ZN(G364));
  AOI21_X1  g0475(.A(new_n261), .B1(new_n603), .B2(G45), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n630), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n221), .B1(G20), .B2(new_n365), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n373), .A2(new_n286), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n222), .A2(G179), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n562), .ZN(new_n685));
  OR3_X1    g0485(.A1(new_n685), .A2(new_n277), .A3(KEYINPUT93), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT93), .B1(new_n685), .B2(new_n277), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n288), .A2(new_n222), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n373), .A2(G200), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n686), .B(new_n687), .C1(new_n212), .C2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n683), .A2(new_n373), .A3(new_n286), .ZN(new_n692));
  INV_X1    g0492(.A(G159), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT32), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n373), .A2(G179), .A3(G200), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n222), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n683), .A2(new_n373), .A3(G200), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n698), .A2(G97), .B1(new_n700), .B2(G107), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n688), .A2(new_n682), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n695), .B(new_n701), .C1(new_n302), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n688), .A2(new_n373), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G200), .ZN(new_n705));
  AOI211_X1 g0505(.A(new_n691), .B(new_n703), .C1(G77), .C2(new_n705), .ZN(new_n706));
  OR3_X1    g0506(.A1(new_n704), .A2(KEYINPUT94), .A3(new_n286), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT94), .B1(new_n704), .B2(new_n286), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n706), .B1(new_n214), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G322), .ZN(new_n712));
  INV_X1    g0512(.A(G326), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n712), .A2(new_n690), .B1(new_n702), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G303), .ZN(new_n715));
  INV_X1    g0515(.A(G283), .ZN(new_n716));
  OAI221_X1 g0516(.A(new_n277), .B1(new_n684), .B2(new_n715), .C1(new_n716), .C2(new_n699), .ZN(new_n717));
  INV_X1    g0517(.A(G294), .ZN(new_n718));
  INV_X1    g0518(.A(G329), .ZN(new_n719));
  OAI22_X1  g0519(.A1(new_n697), .A2(new_n718), .B1(new_n692), .B2(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n714), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G311), .ZN(new_n722));
  INV_X1    g0522(.A(new_n705), .ZN(new_n723));
  XNOR2_X1  g0523(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n724));
  INV_X1    g0524(.A(G317), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n721), .B1(new_n722), .B2(new_n723), .C1(new_n710), .C2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n681), .B1(new_n711), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT92), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n680), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n277), .A2(new_n629), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n734), .A2(G355), .B1(new_n471), .B2(new_n629), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n423), .A2(new_n629), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n634), .B2(G45), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n242), .A2(new_n447), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n679), .B(new_n728), .C1(new_n733), .C2(new_n739), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT96), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n616), .B2(new_n732), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n618), .A2(new_n678), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n616), .A2(new_n617), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(G396));
  NOR2_X1   g0546(.A1(new_n290), .A2(new_n612), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n612), .A2(new_n265), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n287), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(new_n749), .B2(new_n290), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n644), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n672), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n678), .B1(new_n751), .B2(new_n672), .ZN(new_n754));
  INV_X1    g0554(.A(new_n750), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n730), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n680), .A2(new_n729), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n678), .B1(new_n758), .B2(G77), .ZN(new_n759));
  INV_X1    g0559(.A(G137), .ZN(new_n760));
  INV_X1    g0560(.A(G143), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n702), .B1(new_n690), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n723), .A2(new_n693), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n762), .B(new_n763), .C1(G150), .C2(new_n709), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n343), .A2(new_n270), .ZN(new_n767));
  INV_X1    g0567(.A(new_n684), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(G50), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G132), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n214), .A2(new_n699), .B1(new_n692), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(G58), .B2(new_n698), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n766), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n764), .A2(new_n765), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n723), .A2(new_n471), .B1(new_n702), .B2(new_n715), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n709), .B2(G283), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(KEYINPUT97), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n562), .A2(new_n699), .B1(new_n692), .B2(new_n722), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n277), .B1(new_n684), .B2(new_n418), .C1(new_n697), .C2(new_n387), .ZN(new_n780));
  INV_X1    g0580(.A(new_n690), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n779), .B(new_n780), .C1(G294), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT97), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n776), .B2(new_n783), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n773), .A2(new_n774), .B1(new_n778), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n759), .B1(new_n785), .B2(new_n680), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n753), .A2(new_n754), .B1(new_n756), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G384));
  NOR3_X1   g0588(.A1(new_n634), .A2(new_n202), .A3(new_n338), .ZN(new_n789));
  INV_X1    g0589(.A(new_n201), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n214), .ZN(new_n791));
  OAI211_X1 g0591(.A(G1), .B(new_n602), .C1(new_n789), .C2(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(G116), .A3(new_n223), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(KEYINPUT35), .B2(new_n508), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n792), .B1(new_n795), .B2(KEYINPUT36), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(KEYINPUT36), .B2(new_n795), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT101), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n767), .A2(new_n222), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n214), .B1(new_n799), .B2(KEYINPUT7), .ZN(new_n800));
  INV_X1    g0600(.A(new_n346), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n340), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n328), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n347), .A2(new_n259), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n804), .A2(new_n805), .B1(new_n350), .B2(new_n349), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n798), .B1(new_n806), .B2(new_n610), .ZN(new_n807));
  INV_X1    g0607(.A(new_n610), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT16), .B1(new_n802), .B2(new_n340), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n347), .A2(new_n259), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n351), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n808), .A2(new_n811), .A3(KEYINPUT101), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n384), .A2(new_n381), .ZN(new_n814));
  AOI21_X1  g0614(.A(KEYINPUT18), .B1(new_n383), .B2(new_n370), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT37), .B1(new_n378), .B2(new_n379), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n817), .A2(new_n382), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n356), .A2(new_n808), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n811), .A2(new_n366), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n807), .A2(new_n380), .A3(new_n812), .A4(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n818), .A2(new_n819), .B1(new_n821), .B2(KEYINPUT37), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n816), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT38), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT102), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n822), .B1(new_n385), .B2(new_n813), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT38), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n827), .B1(new_n828), .B2(KEYINPUT38), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n816), .A2(KEYINPUT38), .A3(new_n823), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n830), .A2(new_n833), .A3(KEYINPUT39), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n819), .A2(new_n380), .A3(new_n594), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT37), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n819), .A2(new_n382), .A3(new_n817), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT104), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n818), .A2(KEYINPUT104), .A3(new_n819), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n819), .B1(new_n381), .B2(new_n595), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n825), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n829), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n834), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n408), .A2(new_n612), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT103), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n831), .A2(new_n832), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n824), .A2(new_n827), .A3(new_n825), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n830), .A2(new_n833), .A3(KEYINPUT103), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n612), .A2(new_n407), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n408), .A2(new_n413), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n399), .A2(new_n407), .A3(new_n612), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n621), .B(new_n750), .C1(new_n580), .C2(new_n591), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n747), .B(KEYINPUT99), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n857), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT100), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n852), .A2(new_n853), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n595), .A2(new_n808), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n848), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n642), .B(new_n415), .C1(new_n644), .C2(KEYINPUT29), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n868), .A2(new_n600), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n867), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n666), .A2(KEYINPUT105), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT105), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n664), .A2(new_n872), .A3(new_n665), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n871), .A2(new_n662), .A3(new_n670), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n855), .A2(new_n856), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n750), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n852), .A2(new_n853), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT106), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n879), .B1(new_n829), .B2(new_n843), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n874), .A2(KEYINPUT106), .A3(new_n750), .A4(new_n875), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(G330), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n415), .A2(G330), .A3(new_n874), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n885), .B1(new_n878), .B2(new_n879), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n890), .A2(new_n415), .A3(new_n874), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OAI22_X1  g0692(.A1(new_n870), .A2(new_n892), .B1(new_n261), .B2(new_n603), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n893), .A2(KEYINPUT107), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n870), .A2(new_n892), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n893), .B2(KEYINPUT107), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n797), .B1(new_n894), .B2(new_n896), .ZN(G367));
  OR2_X1    g0697(.A1(new_n621), .A2(new_n564), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n581), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n561), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n625), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n535), .B(new_n538), .C1(new_n518), .C2(new_n621), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(KEYINPUT42), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n906), .A2(KEYINPUT108), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n585), .A2(new_n612), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n538), .B1(new_n910), .B2(new_n460), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n621), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n905), .A2(KEYINPUT42), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n906), .A2(KEYINPUT108), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n907), .A2(new_n912), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n902), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n623), .A2(new_n910), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n915), .A2(new_n902), .A3(new_n916), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n630), .B(KEYINPUT41), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n627), .A2(new_n909), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT45), .Z(new_n925));
  NOR2_X1   g0725(.A1(new_n627), .A2(new_n909), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT44), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n623), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n623), .B1(new_n925), .B2(new_n927), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT109), .B1(new_n616), .B2(new_n617), .ZN(new_n932));
  INV_X1    g0732(.A(new_n624), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n903), .B1(new_n622), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n932), .B(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(new_n674), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n923), .B1(new_n937), .B2(new_n673), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n921), .B(new_n922), .C1(new_n938), .C2(new_n676), .ZN(new_n939));
  INV_X1    g0739(.A(new_n736), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n238), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n733), .B1(new_n207), .B2(new_n256), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n678), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n732), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n900), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n768), .A2(KEYINPUT46), .A3(G116), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT46), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n684), .B2(new_n471), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n946), .B(new_n948), .C1(new_n725), .C2(new_n692), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n767), .B1(new_n387), .B2(new_n699), .C1(new_n702), .C2(new_n722), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n949), .B(new_n950), .C1(G303), .C2(new_n781), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n705), .A2(G283), .B1(new_n274), .B2(new_n698), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT110), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n709), .A2(G294), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n951), .B(new_n954), .C1(new_n953), .C2(new_n952), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n709), .A2(G159), .B1(new_n790), .B2(new_n705), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT111), .Z(new_n957));
  OAI221_X1 g0757(.A(new_n272), .B1(new_n684), .B2(new_n212), .C1(new_n697), .C2(new_n214), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n202), .A2(new_n699), .B1(new_n692), .B2(new_n760), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n960), .B1(new_n761), .B2(new_n702), .C1(new_n293), .C2(new_n690), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n955), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT47), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n681), .B1(new_n962), .B2(new_n963), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n943), .B(new_n945), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n939), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(G387));
  AOI21_X1  g0768(.A(new_n940), .B1(new_n234), .B2(G45), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n633), .B2(new_n734), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n249), .A2(new_n302), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT50), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n447), .B1(new_n214), .B2(new_n202), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n972), .A2(new_n633), .A3(new_n973), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n970), .A2(new_n974), .B1(G107), .B2(new_n207), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n679), .B1(new_n975), .B2(new_n733), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n767), .B1(G77), .B2(new_n768), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n302), .B2(new_n690), .C1(new_n693), .C2(new_n702), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n256), .A2(new_n697), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G97), .B2(new_n700), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n293), .B2(new_n692), .C1(new_n723), .C2(new_n214), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n978), .B(new_n981), .C1(new_n297), .C2(new_n709), .ZN(new_n982));
  INV_X1    g0782(.A(new_n702), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n709), .A2(G311), .B1(G322), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT112), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n715), .B2(new_n723), .C1(new_n725), .C2(new_n690), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT48), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n716), .B2(new_n697), .C1(new_n718), .C2(new_n684), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT49), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n767), .B1(new_n471), .B2(new_n699), .C1(new_n713), .C2(new_n692), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n988), .B2(new_n989), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n982), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n976), .B1(new_n622), .B2(new_n944), .C1(new_n993), .C2(new_n681), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n935), .A2(new_n677), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n674), .A2(new_n935), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n630), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n674), .A2(new_n935), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n994), .B(new_n995), .C1(new_n997), .C2(new_n998), .ZN(G393));
  NAND2_X1  g0799(.A1(new_n910), .A2(new_n732), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n733), .B1(new_n387), .B2(new_n207), .C1(new_n246), .C2(new_n940), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n678), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n293), .A2(new_n702), .B1(new_n690), .B2(new_n693), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT51), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n692), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1005), .A2(G143), .B1(new_n768), .B2(G68), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1006), .A2(KEYINPUT113), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n698), .A2(G77), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1008), .B(new_n423), .C1(new_n562), .C2(new_n699), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n705), .A2(new_n249), .B1(new_n1006), .B2(KEYINPUT113), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1004), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n710), .A2(new_n201), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n710), .A2(new_n715), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n722), .A2(new_n690), .B1(new_n702), .B2(new_n725), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT52), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n697), .A2(new_n471), .B1(new_n692), .B2(new_n712), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n277), .B1(new_n684), .B2(new_n716), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(G107), .C2(new_n700), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n705), .A2(G294), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1012), .A2(new_n1013), .B1(new_n1014), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1002), .B1(new_n1024), .B2(new_n680), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n931), .A2(new_n677), .B1(new_n1000), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n936), .A2(new_n630), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n996), .B1(new_n929), .B2(new_n930), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1026), .B1(new_n1027), .B2(new_n1029), .ZN(G390));
  OAI211_X1 g0830(.A(new_n834), .B(new_n845), .C1(new_n861), .C2(new_n847), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n663), .A2(new_n666), .B1(new_n568), .B2(new_n621), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n617), .B1(new_n1032), .B2(new_n668), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(new_n750), .A3(new_n875), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n621), .B(new_n750), .C1(new_n639), .C2(new_n641), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n860), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n875), .B(KEYINPUT114), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n844), .B1(new_n408), .B2(new_n612), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1031), .A2(new_n1034), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n868), .A2(new_n600), .A3(new_n888), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n858), .A2(new_n860), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n875), .B1(new_n1033), .B2(new_n750), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n874), .A2(G330), .A3(new_n750), .A4(new_n875), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1042), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n874), .A2(G330), .A3(new_n750), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1038), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1041), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1031), .A2(new_n1039), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1040), .B(new_n1050), .C1(new_n1051), .C2(new_n1044), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1050), .ZN(new_n1053));
  AND3_X1   g0853(.A1(new_n1031), .A2(new_n1034), .A3(new_n1039), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1044), .B1(new_n1031), .B2(new_n1039), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n1056), .A3(new_n630), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n846), .A2(new_n731), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n690), .A2(new_n471), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n277), .B1(new_n684), .B2(new_n562), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT115), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n1060), .A2(new_n1061), .B1(new_n702), .B2(new_n716), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1059), .B(new_n1062), .C1(new_n1061), .C2(new_n1060), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1008), .B1(new_n214), .B2(new_n699), .C1(new_n718), .C2(new_n692), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G97), .B2(new_n705), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(new_n275), .C2(new_n710), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n684), .A2(new_n293), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT53), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1067), .A2(new_n1068), .B1(new_n1005), .B2(G125), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .C1(new_n201), .C2(new_n699), .ZN(new_n1070));
  XOR2_X1   g0870(.A(KEYINPUT54), .B(G143), .Z(new_n1071));
  AOI21_X1  g0871(.A(new_n1070), .B1(new_n705), .B2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n272), .B1(new_n693), .B2(new_n697), .C1(new_n690), .C2(new_n770), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G128), .B2(new_n983), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1072), .B(new_n1074), .C1(new_n760), .C2(new_n710), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n681), .B1(new_n1066), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n678), .B1(new_n758), .B2(new_n297), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1058), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n677), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1057), .A2(new_n1080), .ZN(G378));
  NAND2_X1  g0881(.A1(new_n599), .A2(new_n319), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n306), .A2(new_n610), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n1085));
  XNOR2_X1  g0885(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1086), .B(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n617), .B(new_n885), .C1(new_n878), .C2(new_n879), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(KEYINPUT120), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n848), .A2(new_n865), .A3(new_n866), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n1089), .B2(KEYINPUT120), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n880), .A2(KEYINPUT120), .A3(G330), .A4(new_n886), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(new_n867), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1090), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1052), .A2(new_n869), .A3(new_n888), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1093), .A2(new_n867), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT120), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n887), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1091), .A2(new_n890), .A3(KEYINPUT120), .A4(G330), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1097), .A2(new_n1099), .A3(new_n1100), .A4(new_n1088), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1095), .A2(new_n1096), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT57), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1095), .A2(KEYINPUT57), .A3(new_n1096), .A4(new_n1101), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n630), .A3(new_n1105), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1088), .A2(new_n731), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT119), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n678), .B1(new_n758), .B2(new_n790), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n423), .A2(G41), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n418), .B2(new_n690), .C1(new_n471), .C2(new_n702), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n700), .A2(G58), .B1(new_n1005), .B2(G283), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n214), .B2(new_n697), .C1(new_n202), .C2(new_n684), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1111), .B(new_n1113), .C1(new_n255), .C2(new_n705), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n387), .B2(new_n710), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT58), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n302), .B1(G33), .B2(G41), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1115), .A2(new_n1116), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1116), .B2(new_n1115), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1005), .A2(G124), .ZN(new_n1120));
  AOI211_X1 g0920(.A(G33), .B(G41), .C1(new_n700), .C2(G159), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n983), .A2(G125), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n781), .A2(G128), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n698), .A2(G150), .B1(new_n768), .B2(new_n1071), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n709), .A2(G132), .B1(G137), .B2(new_n705), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1127), .A2(KEYINPUT116), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(KEYINPUT116), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1125), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT59), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1120), .B(new_n1121), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1119), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1109), .B1(new_n1134), .B2(new_n680), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1107), .A2(new_n1108), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1108), .B1(new_n1107), .B2(new_n1135), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1095), .A2(new_n677), .A3(new_n1101), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1106), .A2(new_n1141), .ZN(G375));
  NAND3_X1  g0942(.A1(new_n1046), .A2(new_n1049), .A3(new_n1041), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1053), .A2(new_n923), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n710), .A2(new_n471), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n277), .B1(new_n684), .B2(new_n387), .C1(new_n202), .C2(new_n699), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n979), .B(new_n1146), .C1(G303), .C2(new_n1005), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n716), .B2(new_n690), .C1(new_n718), .C2(new_n702), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1145), .B(new_n1148), .C1(new_n274), .C2(new_n705), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n767), .B1(G159), .B2(new_n768), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n770), .B2(new_n702), .C1(new_n760), .C2(new_n690), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n700), .A2(G58), .B1(new_n1005), .B2(G128), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n302), .B2(new_n697), .C1(new_n723), .C2(new_n293), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(new_n709), .C2(new_n1071), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n680), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n679), .B1(new_n214), .B2(new_n757), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1038), .B2(new_n729), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n857), .B1(new_n672), .B2(new_n755), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1044), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1036), .B1(new_n1038), .B2(new_n1047), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1161), .A2(new_n1042), .B1(new_n1034), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1159), .B1(new_n1163), .B2(new_n676), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1144), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT121), .ZN(G381));
  NOR2_X1   g0967(.A1(G375), .A2(G378), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT122), .ZN(new_n1170));
  NOR4_X1   g0970(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n1171), .ZN(G407));
  AOI21_X1  g0972(.A(new_n631), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1140), .B1(new_n1173), .B2(new_n1105), .ZN(new_n1174));
  INV_X1    g0974(.A(G378), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(G407), .B(G213), .C1(G343), .C2(new_n1176), .ZN(G409));
  NAND4_X1  g0977(.A1(new_n1095), .A2(new_n923), .A3(new_n1096), .A4(new_n1101), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1107), .A2(new_n1135), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1057), .A2(new_n1179), .A3(new_n1080), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1139), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n611), .A2(G213), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n611), .A2(G213), .A3(G2897), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT60), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1143), .B1(new_n1050), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1163), .A2(KEYINPUT60), .A3(new_n1041), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n630), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT123), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1187), .A2(KEYINPUT123), .A3(new_n630), .A4(new_n1188), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G384), .B1(new_n1193), .B2(new_n1165), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n787), .B(new_n1164), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1182), .A2(KEYINPUT124), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1185), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1182), .A2(KEYINPUT124), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n611), .A2(G213), .A3(G2897), .ZN(new_n1200));
  NOR4_X1   g1000(.A1(new_n1194), .A2(new_n1195), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT61), .B1(new_n1184), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(G375), .A2(G378), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT62), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1204), .A2(new_n1205), .A3(new_n1196), .A4(new_n1183), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1183), .B(new_n1196), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT62), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1203), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(KEYINPUT125), .B1(new_n967), .B2(G390), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(G393), .B(G396), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n967), .B2(G390), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT125), .ZN(new_n1213));
  INV_X1    g1013(.A(G390), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n939), .C2(new_n966), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1210), .A2(new_n1212), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1214), .B1(new_n967), .B2(KEYINPUT126), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT126), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1218), .B(G390), .C1(new_n939), .C2(new_n966), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1219), .A3(new_n1211), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1216), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1209), .A2(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1204), .A2(KEYINPUT63), .A3(new_n1196), .A4(new_n1183), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT63), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1207), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1221), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1203), .A2(new_n1223), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1222), .A2(new_n1227), .ZN(G405));
  INV_X1    g1028(.A(new_n1196), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(KEYINPUT127), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1230), .B1(new_n1168), .B2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1204), .B(new_n1176), .C1(KEYINPUT127), .C2(new_n1229), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n1226), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1226), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(G402));
endmodule


