

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(KEYINPUT28), .ZN(n702) );
  XNOR2_X1 U555 ( .A(n581), .B(KEYINPUT15), .ZN(n895) );
  XNOR2_X1 U556 ( .A(n536), .B(KEYINPUT23), .ZN(n537) );
  AND2_X1 U557 ( .A1(n684), .A2(n958), .ZN(n517) );
  XOR2_X1 U558 ( .A(KEYINPUT95), .B(n687), .Z(n518) );
  AND2_X1 U559 ( .A1(n688), .A2(n518), .ZN(n519) );
  INV_X1 U560 ( .A(n723), .ZN(n708) );
  INV_X1 U561 ( .A(n966), .ZN(n743) );
  NOR2_X1 U562 ( .A1(G651), .A2(n628), .ZN(n646) );
  INV_X1 U563 ( .A(KEYINPUT64), .ZN(n536) );
  NOR2_X1 U564 ( .A1(n798), .A2(n797), .ZN(n799) );
  AND2_X1 U565 ( .A1(n542), .A2(G2104), .ZN(n877) );
  INV_X1 U566 ( .A(n895), .ZN(n964) );
  XOR2_X1 U567 ( .A(KEYINPUT1), .B(n527), .Z(n650) );
  XNOR2_X1 U568 ( .A(n538), .B(n537), .ZN(n541) );
  NOR2_X1 U569 ( .A1(n546), .A2(n545), .ZN(G160) );
  XNOR2_X1 U570 ( .A(KEYINPUT74), .B(KEYINPUT7), .ZN(n535) );
  XOR2_X1 U571 ( .A(KEYINPUT4), .B(KEYINPUT72), .Z(n521) );
  NOR2_X1 U572 ( .A1(G543), .A2(G651), .ZN(n642) );
  NAND2_X1 U573 ( .A1(G89), .A2(n642), .ZN(n520) );
  XNOR2_X1 U574 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U575 ( .A(KEYINPUT71), .B(n522), .ZN(n524) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  INV_X1 U577 ( .A(G651), .ZN(n526) );
  NOR2_X1 U578 ( .A1(n628), .A2(n526), .ZN(n643) );
  NAND2_X1 U579 ( .A1(n643), .A2(G76), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U581 ( .A(n525), .B(KEYINPUT5), .ZN(n533) );
  XNOR2_X1 U582 ( .A(KEYINPUT6), .B(KEYINPUT73), .ZN(n531) );
  NAND2_X1 U583 ( .A1(G51), .A2(n646), .ZN(n529) );
  NOR2_X1 U584 ( .A1(G543), .A2(n526), .ZN(n527) );
  NAND2_X1 U585 ( .A1(G63), .A2(n650), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U587 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U589 ( .A(n535), .B(n534), .ZN(G168) );
  XOR2_X1 U590 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  INV_X1 U591 ( .A(G2105), .ZN(n542) );
  NAND2_X1 U592 ( .A1(G101), .A2(n877), .ZN(n538) );
  NOR2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n539) );
  XOR2_X2 U594 ( .A(KEYINPUT17), .B(n539), .Z(n878) );
  NAND2_X1 U595 ( .A1(G137), .A2(n878), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n546) );
  AND2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  NAND2_X1 U598 ( .A1(G113), .A2(n881), .ZN(n544) );
  NOR2_X1 U599 ( .A1(G2104), .A2(n542), .ZN(n882) );
  NAND2_X1 U600 ( .A1(G125), .A2(n882), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G52), .A2(n646), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G64), .A2(n650), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U605 ( .A(KEYINPUT66), .B(n549), .ZN(n555) );
  NAND2_X1 U606 ( .A1(G90), .A2(n642), .ZN(n551) );
  NAND2_X1 U607 ( .A1(G77), .A2(n643), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U609 ( .A(KEYINPUT9), .B(n552), .ZN(n553) );
  XNOR2_X1 U610 ( .A(KEYINPUT67), .B(n553), .ZN(n554) );
  NOR2_X1 U611 ( .A1(n555), .A2(n554), .ZN(G171) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U613 ( .A(G132), .ZN(G219) );
  INV_X1 U614 ( .A(G82), .ZN(G220) );
  NAND2_X1 U615 ( .A1(n877), .A2(G102), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G114), .A2(n881), .ZN(n556) );
  XOR2_X1 U617 ( .A(KEYINPUT85), .B(n556), .Z(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G138), .A2(n878), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G126), .A2(n882), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U622 ( .A1(n562), .A2(n561), .ZN(G164) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U624 ( .A(n563), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U625 ( .A(G223), .ZN(n825) );
  NAND2_X1 U626 ( .A1(n825), .A2(G567), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U628 ( .A1(n642), .A2(G81), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G68), .A2(n643), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U632 ( .A(n568), .B(KEYINPUT13), .ZN(n570) );
  NAND2_X1 U633 ( .A1(G43), .A2(n646), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n650), .A2(G56), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n571), .Z(n572) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n958) );
  NAND2_X1 U638 ( .A1(n958), .A2(G860), .ZN(G153) );
  INV_X1 U639 ( .A(G171), .ZN(G301) );
  NAND2_X1 U640 ( .A1(G868), .A2(G301), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G92), .A2(n642), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G66), .A2(n650), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U644 ( .A(KEYINPUT70), .B(n576), .ZN(n580) );
  NAND2_X1 U645 ( .A1(G54), .A2(n646), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G79), .A2(n643), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  INV_X1 U649 ( .A(G868), .ZN(n663) );
  NAND2_X1 U650 ( .A1(n895), .A2(n663), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(G284) );
  NAND2_X1 U652 ( .A1(G53), .A2(n646), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G65), .A2(n650), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U655 ( .A(KEYINPUT68), .B(n586), .Z(n590) );
  NAND2_X1 U656 ( .A1(G91), .A2(n642), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G78), .A2(n643), .ZN(n587) );
  AND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(G299) );
  NAND2_X1 U660 ( .A1(G868), .A2(G286), .ZN(n592) );
  NAND2_X1 U661 ( .A1(G299), .A2(n663), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n592), .A2(n591), .ZN(G297) );
  INV_X1 U663 ( .A(G860), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n593), .A2(G559), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n594), .A2(n964), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n595), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U667 ( .A1(n964), .A2(G868), .ZN(n596) );
  NOR2_X1 U668 ( .A1(G559), .A2(n596), .ZN(n598) );
  AND2_X1 U669 ( .A1(n663), .A2(n958), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(G282) );
  NAND2_X1 U671 ( .A1(G99), .A2(n877), .ZN(n600) );
  NAND2_X1 U672 ( .A1(G111), .A2(n881), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n606) );
  NAND2_X1 U674 ( .A1(n882), .A2(G123), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT18), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G135), .A2(n878), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U678 ( .A(KEYINPUT75), .B(n604), .Z(n605) );
  NOR2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U680 ( .A(KEYINPUT76), .B(n607), .ZN(n912) );
  XOR2_X1 U681 ( .A(G2096), .B(KEYINPUT77), .Z(n608) );
  XNOR2_X1 U682 ( .A(n912), .B(n608), .ZN(n610) );
  INV_X1 U683 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U685 ( .A1(G93), .A2(n642), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G80), .A2(n643), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U688 ( .A(KEYINPUT78), .B(n613), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G55), .A2(n646), .ZN(n615) );
  NAND2_X1 U690 ( .A1(G67), .A2(n650), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n616) );
  OR2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n664) );
  NAND2_X1 U693 ( .A1(n964), .A2(G559), .ZN(n660) );
  XOR2_X1 U694 ( .A(n958), .B(n660), .Z(n618) );
  NOR2_X1 U695 ( .A1(G860), .A2(n618), .ZN(n619) );
  XOR2_X1 U696 ( .A(n664), .B(n619), .Z(G145) );
  NAND2_X1 U697 ( .A1(G61), .A2(n650), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n620), .B(KEYINPUT80), .ZN(n627) );
  NAND2_X1 U699 ( .A1(G48), .A2(n646), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G86), .A2(n642), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n643), .A2(G73), .ZN(n623) );
  XOR2_X1 U703 ( .A(KEYINPUT2), .B(n623), .Z(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(G305) );
  NAND2_X1 U706 ( .A1(G49), .A2(n646), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G87), .A2(n628), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n650), .A2(n631), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n632) );
  XOR2_X1 U711 ( .A(KEYINPUT79), .B(n632), .Z(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U713 ( .A1(G50), .A2(n646), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G62), .A2(n650), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G88), .A2(n642), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G75), .A2(n643), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U719 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U720 ( .A(n641), .B(KEYINPUT81), .ZN(G303) );
  INV_X1 U721 ( .A(G303), .ZN(G166) );
  NAND2_X1 U722 ( .A1(G85), .A2(n642), .ZN(n645) );
  NAND2_X1 U723 ( .A1(G72), .A2(n643), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U725 ( .A1(G47), .A2(n646), .ZN(n647) );
  XNOR2_X1 U726 ( .A(KEYINPUT65), .B(n647), .ZN(n648) );
  NOR2_X1 U727 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n650), .A2(G60), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(G290) );
  XOR2_X1 U730 ( .A(KEYINPUT19), .B(KEYINPUT82), .Z(n653) );
  XNOR2_X1 U731 ( .A(G288), .B(n653), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(n664), .ZN(n656) );
  INV_X1 U733 ( .A(G299), .ZN(n701) );
  XNOR2_X1 U734 ( .A(n701), .B(G166), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U736 ( .A(n657), .B(G290), .Z(n658) );
  XNOR2_X1 U737 ( .A(G305), .B(n658), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n958), .B(n659), .ZN(n896) );
  XNOR2_X1 U739 ( .A(n896), .B(n660), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n661), .A2(G868), .ZN(n662) );
  XOR2_X1 U741 ( .A(KEYINPUT83), .B(n662), .Z(n666) );
  NAND2_X1 U742 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U743 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U748 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U750 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U753 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U754 ( .A1(G96), .A2(n673), .ZN(n829) );
  NAND2_X1 U755 ( .A1(G2106), .A2(n829), .ZN(n674) );
  XNOR2_X1 U756 ( .A(n674), .B(KEYINPUT84), .ZN(n678) );
  NAND2_X1 U757 ( .A1(G120), .A2(G69), .ZN(n675) );
  NOR2_X1 U758 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U759 ( .A1(G108), .A2(n676), .ZN(n830) );
  NAND2_X1 U760 ( .A1(G567), .A2(n830), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n678), .A2(n677), .ZN(n831) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U763 ( .A1(n831), .A2(n679), .ZN(n828) );
  NAND2_X1 U764 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n762) );
  INV_X1 U766 ( .A(n762), .ZN(n693) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n763) );
  NAND2_X1 U768 ( .A1(n693), .A2(n763), .ZN(n723) );
  NAND2_X1 U769 ( .A1(G8), .A2(n723), .ZN(n757) );
  NOR2_X1 U770 ( .A1(G1981), .A2(G305), .ZN(n680) );
  XOR2_X1 U771 ( .A(n680), .B(KEYINPUT24), .Z(n681) );
  NOR2_X1 U772 ( .A1(n757), .A2(n681), .ZN(n761) );
  XNOR2_X1 U773 ( .A(G1981), .B(KEYINPUT100), .ZN(n682) );
  XNOR2_X1 U774 ( .A(n682), .B(G305), .ZN(n977) );
  NAND2_X1 U775 ( .A1(G1996), .A2(n708), .ZN(n683) );
  XNOR2_X1 U776 ( .A(KEYINPUT26), .B(n683), .ZN(n684) );
  NOR2_X1 U777 ( .A1(n708), .A2(G1348), .ZN(n686) );
  NOR2_X1 U778 ( .A1(G2067), .A2(n723), .ZN(n685) );
  NOR2_X1 U779 ( .A1(n686), .A2(n685), .ZN(n689) );
  NAND2_X1 U780 ( .A1(n689), .A2(n895), .ZN(n688) );
  NAND2_X1 U781 ( .A1(G1341), .A2(n723), .ZN(n687) );
  NAND2_X1 U782 ( .A1(n517), .A2(n519), .ZN(n691) );
  OR2_X1 U783 ( .A1(n689), .A2(n895), .ZN(n690) );
  AND2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n699) );
  AND2_X1 U785 ( .A1(G2072), .A2(n763), .ZN(n692) );
  NAND2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(KEYINPUT27), .ZN(n695) );
  XNOR2_X1 U788 ( .A(KEYINPUT94), .B(n695), .ZN(n697) );
  INV_X1 U789 ( .A(G1956), .ZN(n990) );
  NOR2_X1 U790 ( .A1(n708), .A2(n990), .ZN(n696) );
  NOR2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n698) );
  NAND2_X1 U793 ( .A1(n699), .A2(n698), .ZN(n705) );
  NOR2_X1 U794 ( .A1(n701), .A2(n700), .ZN(n703) );
  XNOR2_X1 U795 ( .A(n703), .B(n702), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U797 ( .A(KEYINPUT29), .B(n706), .Z(n712) );
  NOR2_X1 U798 ( .A1(n708), .A2(G1961), .ZN(n707) );
  XNOR2_X1 U799 ( .A(n707), .B(KEYINPUT93), .ZN(n710) );
  XNOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .ZN(n935) );
  NAND2_X1 U801 ( .A1(n708), .A2(n935), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n716) );
  NAND2_X1 U803 ( .A1(n716), .A2(G171), .ZN(n711) );
  NAND2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n721) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n757), .ZN(n734) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n723), .ZN(n731) );
  NOR2_X1 U807 ( .A1(n734), .A2(n731), .ZN(n713) );
  NAND2_X1 U808 ( .A1(G8), .A2(n713), .ZN(n714) );
  XNOR2_X1 U809 ( .A(KEYINPUT30), .B(n714), .ZN(n715) );
  NOR2_X1 U810 ( .A1(G168), .A2(n715), .ZN(n718) );
  NOR2_X1 U811 ( .A1(G171), .A2(n716), .ZN(n717) );
  NOR2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U813 ( .A(KEYINPUT31), .B(n719), .Z(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n732) );
  NAND2_X1 U815 ( .A1(n732), .A2(G286), .ZN(n728) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n757), .ZN(n722) );
  XNOR2_X1 U817 ( .A(n722), .B(KEYINPUT96), .ZN(n725) );
  NOR2_X1 U818 ( .A1(n723), .A2(G2090), .ZN(n724) );
  NOR2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n726), .A2(G303), .ZN(n727) );
  NAND2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U822 ( .A1(n729), .A2(G8), .ZN(n730) );
  XNOR2_X1 U823 ( .A(n730), .B(KEYINPUT32), .ZN(n738) );
  NAND2_X1 U824 ( .A1(G8), .A2(n731), .ZN(n736) );
  INV_X1 U825 ( .A(n732), .ZN(n733) );
  NOR2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n753) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n739) );
  XOR2_X1 U830 ( .A(KEYINPUT97), .B(n739), .Z(n748) );
  NOR2_X1 U831 ( .A1(G1971), .A2(G303), .ZN(n740) );
  NOR2_X1 U832 ( .A1(n748), .A2(n740), .ZN(n962) );
  NAND2_X1 U833 ( .A1(n753), .A2(n962), .ZN(n741) );
  XNOR2_X1 U834 ( .A(n741), .B(KEYINPUT98), .ZN(n745) );
  NAND2_X1 U835 ( .A1(G288), .A2(G1976), .ZN(n742) );
  XOR2_X1 U836 ( .A(KEYINPUT99), .B(n742), .Z(n966) );
  NOR2_X1 U837 ( .A1(n757), .A2(n743), .ZN(n744) );
  AND2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U839 ( .A1(KEYINPUT33), .A2(n746), .ZN(n747) );
  NOR2_X1 U840 ( .A1(n977), .A2(n747), .ZN(n752) );
  INV_X1 U841 ( .A(n748), .ZN(n749) );
  NOR2_X1 U842 ( .A1(n757), .A2(n749), .ZN(n750) );
  NAND2_X1 U843 ( .A1(KEYINPUT33), .A2(n750), .ZN(n751) );
  NAND2_X1 U844 ( .A1(n752), .A2(n751), .ZN(n759) );
  NOR2_X1 U845 ( .A1(G2090), .A2(G303), .ZN(n754) );
  NAND2_X1 U846 ( .A1(G8), .A2(n754), .ZN(n755) );
  NAND2_X1 U847 ( .A1(n753), .A2(n755), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n798) );
  NOR2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n811) );
  XOR2_X1 U852 ( .A(G2067), .B(KEYINPUT37), .Z(n764) );
  XNOR2_X1 U853 ( .A(KEYINPUT87), .B(n764), .ZN(n808) );
  NAND2_X1 U854 ( .A1(G104), .A2(n877), .ZN(n766) );
  NAND2_X1 U855 ( .A1(G140), .A2(n878), .ZN(n765) );
  NAND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U857 ( .A(KEYINPUT34), .B(n767), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n882), .A2(G128), .ZN(n768) );
  XNOR2_X1 U859 ( .A(n768), .B(KEYINPUT88), .ZN(n770) );
  NAND2_X1 U860 ( .A1(G116), .A2(n881), .ZN(n769) );
  NAND2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U862 ( .A(n771), .B(KEYINPUT35), .Z(n772) );
  NOR2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U864 ( .A(KEYINPUT36), .B(n774), .Z(n775) );
  XNOR2_X1 U865 ( .A(KEYINPUT89), .B(n775), .ZN(n891) );
  NOR2_X1 U866 ( .A1(n808), .A2(n891), .ZN(n925) );
  NAND2_X1 U867 ( .A1(n811), .A2(n925), .ZN(n806) );
  NAND2_X1 U868 ( .A1(G105), .A2(n877), .ZN(n776) );
  XNOR2_X1 U869 ( .A(n776), .B(KEYINPUT38), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G117), .A2(n881), .ZN(n778) );
  NAND2_X1 U871 ( .A1(G141), .A2(n878), .ZN(n777) );
  NAND2_X1 U872 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U873 ( .A1(G129), .A2(n882), .ZN(n779) );
  XNOR2_X1 U874 ( .A(KEYINPUT91), .B(n779), .ZN(n780) );
  NOR2_X1 U875 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n874) );
  NAND2_X1 U877 ( .A1(G1996), .A2(n874), .ZN(n792) );
  NAND2_X1 U878 ( .A1(G107), .A2(n881), .ZN(n785) );
  NAND2_X1 U879 ( .A1(G119), .A2(n882), .ZN(n784) );
  NAND2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U881 ( .A(KEYINPUT90), .B(n786), .Z(n790) );
  NAND2_X1 U882 ( .A1(G95), .A2(n877), .ZN(n788) );
  NAND2_X1 U883 ( .A1(G131), .A2(n878), .ZN(n787) );
  AND2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n888) );
  NAND2_X1 U886 ( .A1(G1991), .A2(n888), .ZN(n791) );
  NAND2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n913) );
  NAND2_X1 U888 ( .A1(n811), .A2(n913), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n806), .A2(n800), .ZN(n793) );
  XOR2_X1 U890 ( .A(KEYINPUT92), .B(n793), .Z(n796) );
  XNOR2_X1 U891 ( .A(G1986), .B(KEYINPUT86), .ZN(n794) );
  XNOR2_X1 U892 ( .A(n794), .B(G290), .ZN(n961) );
  NAND2_X1 U893 ( .A1(n811), .A2(n961), .ZN(n795) );
  NAND2_X1 U894 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U895 ( .A(n799), .B(KEYINPUT101), .ZN(n813) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n874), .ZN(n918) );
  INV_X1 U897 ( .A(n800), .ZN(n803) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n888), .ZN(n914) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n801) );
  NOR2_X1 U900 ( .A1(n914), .A2(n801), .ZN(n802) );
  NOR2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U902 ( .A1(n918), .A2(n804), .ZN(n805) );
  XNOR2_X1 U903 ( .A(n805), .B(KEYINPUT39), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n808), .A2(n891), .ZN(n922) );
  NAND2_X1 U906 ( .A1(n809), .A2(n922), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U909 ( .A(n814), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U910 ( .A(G2454), .B(G2446), .ZN(n823) );
  XNOR2_X1 U911 ( .A(G2430), .B(G2443), .ZN(n821) );
  XOR2_X1 U912 ( .A(G2435), .B(KEYINPUT102), .Z(n816) );
  XNOR2_X1 U913 ( .A(G2451), .B(G2438), .ZN(n815) );
  XNOR2_X1 U914 ( .A(n816), .B(n815), .ZN(n817) );
  XOR2_X1 U915 ( .A(n817), .B(G2427), .Z(n819) );
  XNOR2_X1 U916 ( .A(G1348), .B(G1341), .ZN(n818) );
  XNOR2_X1 U917 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U918 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U919 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n824), .A2(G14), .ZN(n900) );
  XNOR2_X1 U921 ( .A(KEYINPUT103), .B(n900), .ZN(G401) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U924 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U926 ( .A1(n828), .A2(n827), .ZN(G188) );
  XOR2_X1 U927 ( .A(G69), .B(KEYINPUT104), .Z(G235) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G108), .ZN(G238) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U934 ( .A(KEYINPUT105), .B(n831), .ZN(G319) );
  XOR2_X1 U935 ( .A(G2096), .B(KEYINPUT43), .Z(n833) );
  XNOR2_X1 U936 ( .A(G2072), .B(KEYINPUT106), .ZN(n832) );
  XNOR2_X1 U937 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U938 ( .A(n834), .B(G2678), .Z(n836) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2090), .ZN(n835) );
  XNOR2_X1 U940 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U941 ( .A(KEYINPUT42), .B(G2100), .Z(n838) );
  XNOR2_X1 U942 ( .A(G2078), .B(G2084), .ZN(n837) );
  XNOR2_X1 U943 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U944 ( .A(n840), .B(n839), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1976), .B(G1971), .Z(n842) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1961), .ZN(n841) );
  XNOR2_X1 U947 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U948 ( .A(G1981), .B(G1966), .Z(n844) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U950 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U951 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U952 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n847) );
  XNOR2_X1 U953 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U954 ( .A(G2474), .B(n849), .ZN(n850) );
  XNOR2_X1 U955 ( .A(n850), .B(n990), .ZN(G229) );
  NAND2_X1 U956 ( .A1(n882), .A2(G124), .ZN(n851) );
  XNOR2_X1 U957 ( .A(n851), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U958 ( .A1(G136), .A2(n878), .ZN(n852) );
  NAND2_X1 U959 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U960 ( .A(KEYINPUT108), .B(n854), .ZN(n858) );
  NAND2_X1 U961 ( .A1(G100), .A2(n877), .ZN(n856) );
  NAND2_X1 U962 ( .A1(G112), .A2(n881), .ZN(n855) );
  NAND2_X1 U963 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U964 ( .A1(n858), .A2(n857), .ZN(G162) );
  NAND2_X1 U965 ( .A1(G106), .A2(n877), .ZN(n860) );
  NAND2_X1 U966 ( .A1(G142), .A2(n878), .ZN(n859) );
  NAND2_X1 U967 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U968 ( .A(n861), .B(KEYINPUT45), .ZN(n863) );
  NAND2_X1 U969 ( .A1(G118), .A2(n881), .ZN(n862) );
  NAND2_X1 U970 ( .A1(n863), .A2(n862), .ZN(n866) );
  NAND2_X1 U971 ( .A1(G130), .A2(n882), .ZN(n864) );
  XNOR2_X1 U972 ( .A(KEYINPUT109), .B(n864), .ZN(n865) );
  NOR2_X1 U973 ( .A1(n866), .A2(n865), .ZN(n876) );
  XOR2_X1 U974 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n868) );
  XNOR2_X1 U975 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n867) );
  XNOR2_X1 U976 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U977 ( .A(n869), .B(KEYINPUT110), .Z(n871) );
  XNOR2_X1 U978 ( .A(G160), .B(G162), .ZN(n870) );
  XNOR2_X1 U979 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U980 ( .A(G164), .B(n872), .Z(n873) );
  XNOR2_X1 U981 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U982 ( .A(n876), .B(n875), .ZN(n890) );
  NAND2_X1 U983 ( .A1(G103), .A2(n877), .ZN(n880) );
  NAND2_X1 U984 ( .A1(G139), .A2(n878), .ZN(n879) );
  NAND2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G115), .A2(n881), .ZN(n884) );
  NAND2_X1 U987 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U988 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n907) );
  XNOR2_X1 U991 ( .A(n888), .B(n907), .ZN(n889) );
  XNOR2_X1 U992 ( .A(n890), .B(n889), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n893), .B(n912), .ZN(n894) );
  NOR2_X1 U995 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n897), .B(G286), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n898), .B(G171), .ZN(n899) );
  NOR2_X1 U999 ( .A1(G37), .A2(n899), .ZN(G397) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n900), .ZN(n903) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n901), .B(KEYINPUT49), .ZN(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(KEYINPUT113), .B(n904), .Z(n906) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n905) );
  NAND2_X1 U1006 ( .A1(n906), .A2(n905), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1008 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1018) );
  XNOR2_X1 U1009 ( .A(KEYINPUT52), .B(KEYINPUT115), .ZN(n930) );
  XOR2_X1 U1010 ( .A(G2072), .B(n907), .Z(n909) );
  XOR2_X1 U1011 ( .A(G164), .B(G2078), .Z(n908) );
  NOR2_X1 U1012 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1013 ( .A(KEYINPUT50), .B(n910), .ZN(n928) );
  XOR2_X1 U1014 ( .A(G160), .B(G2084), .Z(n911) );
  NOR2_X1 U1015 ( .A1(n912), .A2(n911), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n921) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(n919), .B(KEYINPUT51), .ZN(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT114), .B(n926), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n930), .B(n929), .ZN(n931) );
  INV_X1 U1027 ( .A(KEYINPUT55), .ZN(n953) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n953), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n932), .A2(G29), .ZN(n1016) );
  XNOR2_X1 U1030 ( .A(G2090), .B(G35), .ZN(n948) );
  XOR2_X1 U1031 ( .A(G1991), .B(G25), .Z(n933) );
  NAND2_X1 U1032 ( .A1(G28), .A2(n933), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(KEYINPUT116), .B(n934), .ZN(n945) );
  XNOR2_X1 U1034 ( .A(G27), .B(n935), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(G2072), .B(G33), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1038 ( .A(KEYINPUT117), .B(n938), .Z(n939) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G32), .B(G1996), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1042 ( .A(KEYINPUT118), .B(n943), .Z(n944) );
  NOR2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(KEYINPUT53), .B(n946), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1046 ( .A(G2084), .B(G34), .Z(n949) );
  XNOR2_X1 U1047 ( .A(KEYINPUT54), .B(n949), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(n953), .B(n952), .ZN(n955) );
  INV_X1 U1050 ( .A(G29), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(G11), .A2(n956), .ZN(n1014) );
  INV_X1 U1053 ( .A(G16), .ZN(n1010) );
  XNOR2_X1 U1054 ( .A(KEYINPUT56), .B(KEYINPUT119), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(n1010), .B(n957), .ZN(n982) );
  XOR2_X1 U1056 ( .A(n958), .B(G1341), .Z(n959) );
  XNOR2_X1 U1057 ( .A(KEYINPUT120), .B(n959), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n974) );
  XNOR2_X1 U1059 ( .A(G171), .B(G1961), .ZN(n963) );
  NAND2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(G1348), .B(n964), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(G1971), .A2(G303), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(G1956), .B(G299), .ZN(n967) );
  NOR2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(KEYINPUT121), .B(n975), .ZN(n980) );
  XOR2_X1 U1070 ( .A(G1966), .B(G168), .Z(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1072 ( .A(KEYINPUT57), .B(n978), .Z(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n1012) );
  XOR2_X1 U1075 ( .A(G1986), .B(G24), .Z(n984) );
  XOR2_X1 U1076 ( .A(G1971), .B(G22), .Z(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(G23), .B(G1976), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1080 ( .A(KEYINPUT58), .B(n987), .Z(n1007) );
  XOR2_X1 U1081 ( .A(G1961), .B(G5), .Z(n1002) );
  XOR2_X1 U1082 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n1000) );
  XOR2_X1 U1083 ( .A(KEYINPUT124), .B(G4), .Z(n989) );
  XNOR2_X1 U1084 ( .A(G1348), .B(KEYINPUT59), .ZN(n988) );
  XNOR2_X1 U1085 ( .A(n989), .B(n988), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G20), .B(n990), .ZN(n993) );
  XOR2_X1 U1087 ( .A(G1341), .B(G19), .Z(n991) );
  XNOR2_X1 U1088 ( .A(KEYINPUT122), .B(n991), .ZN(n992) );
  NAND2_X1 U1089 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1090 ( .A(G6), .B(G1981), .ZN(n994) );
  NOR2_X1 U1091 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1092 ( .A(n996), .B(KEYINPUT123), .ZN(n997) );
  NOR2_X1 U1093 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1094 ( .A(n1000), .B(n999), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1096 ( .A(G21), .B(G1966), .ZN(n1003) );
  NOR2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1098 ( .A(KEYINPUT126), .B(n1005), .Z(n1006) );
  NOR2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1100 ( .A(KEYINPUT61), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(n1018), .B(n1017), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

