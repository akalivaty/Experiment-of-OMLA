

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X4 U550 ( .A1(n520), .A2(G2105), .ZN(n884) );
  OR2_X1 U551 ( .A1(n698), .A2(n697), .ZN(n696) );
  NOR2_X1 U552 ( .A1(G651), .A2(n628), .ZN(n636) );
  NOR2_X1 U553 ( .A1(G2105), .A2(G2104), .ZN(n516) );
  XOR2_X1 U554 ( .A(KEYINPUT17), .B(n516), .Z(n883) );
  NAND2_X1 U555 ( .A1(n883), .A2(G137), .ZN(n519) );
  XOR2_X1 U556 ( .A(G2104), .B(KEYINPUT66), .Z(n520) );
  NAND2_X1 U557 ( .A1(G101), .A2(n884), .ZN(n517) );
  XOR2_X1 U558 ( .A(KEYINPUT23), .B(n517), .Z(n518) );
  NAND2_X1 U559 ( .A1(n519), .A2(n518), .ZN(n524) );
  AND2_X1 U560 ( .A1(G2105), .A2(n520), .ZN(n879) );
  NAND2_X1 U561 ( .A1(G125), .A2(n879), .ZN(n522) );
  AND2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n880) );
  NAND2_X1 U563 ( .A1(G113), .A2(n880), .ZN(n521) );
  NAND2_X1 U564 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X2 U565 ( .A1(n524), .A2(n523), .ZN(G160) );
  INV_X1 U566 ( .A(G651), .ZN(n529) );
  NOR2_X1 U567 ( .A1(G543), .A2(n529), .ZN(n525) );
  XOR2_X1 U568 ( .A(KEYINPUT1), .B(n525), .Z(n635) );
  NAND2_X1 U569 ( .A1(G64), .A2(n635), .ZN(n527) );
  XOR2_X1 U570 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  NAND2_X1 U571 ( .A1(G52), .A2(n636), .ZN(n526) );
  NAND2_X1 U572 ( .A1(n527), .A2(n526), .ZN(n534) );
  NOR2_X1 U573 ( .A1(G651), .A2(G543), .ZN(n631) );
  NAND2_X1 U574 ( .A1(n631), .A2(G90), .ZN(n528) );
  XOR2_X1 U575 ( .A(KEYINPUT69), .B(n528), .Z(n531) );
  NOR2_X1 U576 ( .A1(n628), .A2(n529), .ZN(n632) );
  NAND2_X1 U577 ( .A1(n632), .A2(G77), .ZN(n530) );
  NAND2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U579 ( .A(KEYINPUT9), .B(n532), .Z(n533) );
  NOR2_X1 U580 ( .A1(n534), .A2(n533), .ZN(G171) );
  AND2_X1 U581 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U582 ( .A1(n883), .A2(G135), .ZN(n535) );
  XNOR2_X1 U583 ( .A(KEYINPUT80), .B(n535), .ZN(n538) );
  NAND2_X1 U584 ( .A1(n879), .A2(G123), .ZN(n536) );
  XNOR2_X1 U585 ( .A(KEYINPUT18), .B(n536), .ZN(n537) );
  NAND2_X1 U586 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U587 ( .A(KEYINPUT81), .B(n539), .ZN(n544) );
  NAND2_X1 U588 ( .A1(G111), .A2(n880), .ZN(n541) );
  NAND2_X1 U589 ( .A1(G99), .A2(n884), .ZN(n540) );
  NAND2_X1 U590 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U591 ( .A(KEYINPUT82), .B(n542), .Z(n543) );
  NAND2_X1 U592 ( .A1(n544), .A2(n543), .ZN(n974) );
  XNOR2_X1 U593 ( .A(G2096), .B(n974), .ZN(n545) );
  OR2_X1 U594 ( .A1(G2100), .A2(n545), .ZN(G156) );
  INV_X1 U595 ( .A(G57), .ZN(G237) );
  INV_X1 U596 ( .A(G132), .ZN(G219) );
  INV_X1 U597 ( .A(G82), .ZN(G220) );
  NAND2_X1 U598 ( .A1(G63), .A2(n635), .ZN(n547) );
  NAND2_X1 U599 ( .A1(G51), .A2(n636), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U601 ( .A(KEYINPUT6), .B(n548), .ZN(n555) );
  NAND2_X1 U602 ( .A1(n631), .A2(G89), .ZN(n549) );
  XNOR2_X1 U603 ( .A(KEYINPUT4), .B(n549), .ZN(n552) );
  NAND2_X1 U604 ( .A1(n632), .A2(G76), .ZN(n550) );
  XOR2_X1 U605 ( .A(KEYINPUT77), .B(n550), .Z(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U607 ( .A(n553), .B(KEYINPUT5), .Z(n554) );
  NOR2_X1 U608 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U609 ( .A(KEYINPUT78), .B(n556), .Z(n557) );
  XNOR2_X1 U610 ( .A(KEYINPUT7), .B(n557), .ZN(G168) );
  XOR2_X1 U611 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U612 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U613 ( .A(n558), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U614 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n560) );
  INV_X1 U615 ( .A(G223), .ZN(n825) );
  NAND2_X1 U616 ( .A1(G567), .A2(n825), .ZN(n559) );
  XNOR2_X1 U617 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U618 ( .A(KEYINPUT72), .B(n561), .Z(G234) );
  INV_X1 U619 ( .A(G860), .ZN(n593) );
  NAND2_X1 U620 ( .A1(n631), .A2(G81), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G68), .A2(n632), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n564), .A2(n563), .ZN(n566) );
  XOR2_X1 U624 ( .A(KEYINPUT74), .B(KEYINPUT13), .Z(n565) );
  XNOR2_X1 U625 ( .A(n566), .B(n565), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n635), .A2(G56), .ZN(n567) );
  XOR2_X1 U627 ( .A(KEYINPUT14), .B(n567), .Z(n568) );
  NOR2_X1 U628 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n636), .A2(G43), .ZN(n570) );
  NAND2_X1 U630 ( .A1(n571), .A2(n570), .ZN(n937) );
  NOR2_X1 U631 ( .A1(n593), .A2(n937), .ZN(n572) );
  XNOR2_X1 U632 ( .A(n572), .B(KEYINPUT75), .ZN(G153) );
  INV_X1 U633 ( .A(G171), .ZN(G301) );
  NAND2_X1 U634 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U635 ( .A1(G54), .A2(n636), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G92), .A2(n631), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G66), .A2(n635), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n632), .A2(G79), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT76), .B(n575), .Z(n576) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U643 ( .A(n580), .B(KEYINPUT15), .ZN(n943) );
  INV_X1 U644 ( .A(n943), .ZN(n698) );
  INV_X1 U645 ( .A(G868), .ZN(n596) );
  NAND2_X1 U646 ( .A1(n698), .A2(n596), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U648 ( .A1(G91), .A2(n631), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n583), .B(KEYINPUT70), .ZN(n590) );
  NAND2_X1 U650 ( .A1(G65), .A2(n635), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G53), .A2(n636), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G78), .A2(n632), .ZN(n586) );
  XNOR2_X1 U654 ( .A(KEYINPUT71), .B(n586), .ZN(n587) );
  NOR2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(G299) );
  NAND2_X1 U657 ( .A1(G868), .A2(G286), .ZN(n592) );
  NAND2_X1 U658 ( .A1(G299), .A2(n596), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n592), .A2(n591), .ZN(G297) );
  NAND2_X1 U660 ( .A1(n593), .A2(G559), .ZN(n594) );
  NAND2_X1 U661 ( .A1(n594), .A2(n943), .ZN(n595) );
  XNOR2_X1 U662 ( .A(n595), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U663 ( .A1(G559), .A2(n596), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n943), .A2(n597), .ZN(n598) );
  XNOR2_X1 U665 ( .A(n598), .B(KEYINPUT79), .ZN(n600) );
  NOR2_X1 U666 ( .A1(n937), .A2(G868), .ZN(n599) );
  NOR2_X1 U667 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U668 ( .A1(G86), .A2(n631), .ZN(n602) );
  NAND2_X1 U669 ( .A1(G61), .A2(n635), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U671 ( .A1(n632), .A2(G73), .ZN(n603) );
  XOR2_X1 U672 ( .A(KEYINPUT2), .B(n603), .Z(n604) );
  NOR2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U674 ( .A1(n636), .A2(G48), .ZN(n606) );
  NAND2_X1 U675 ( .A1(n607), .A2(n606), .ZN(G305) );
  NAND2_X1 U676 ( .A1(n635), .A2(G62), .ZN(n614) );
  NAND2_X1 U677 ( .A1(G88), .A2(n631), .ZN(n609) );
  NAND2_X1 U678 ( .A1(G75), .A2(n632), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n636), .A2(G50), .ZN(n610) );
  XOR2_X1 U681 ( .A(KEYINPUT86), .B(n610), .Z(n611) );
  NOR2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U684 ( .A(KEYINPUT87), .B(n615), .Z(G303) );
  INV_X1 U685 ( .A(G303), .ZN(G166) );
  NAND2_X1 U686 ( .A1(n631), .A2(G85), .ZN(n616) );
  XOR2_X1 U687 ( .A(KEYINPUT67), .B(n616), .Z(n618) );
  NAND2_X1 U688 ( .A1(n632), .A2(G72), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U690 ( .A(KEYINPUT68), .B(n619), .Z(n623) );
  NAND2_X1 U691 ( .A1(G60), .A2(n635), .ZN(n621) );
  NAND2_X1 U692 ( .A1(G47), .A2(n636), .ZN(n620) );
  AND2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n623), .A2(n622), .ZN(G290) );
  NAND2_X1 U695 ( .A1(G49), .A2(n636), .ZN(n625) );
  NAND2_X1 U696 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U698 ( .A1(n635), .A2(n626), .ZN(n627) );
  XOR2_X1 U699 ( .A(KEYINPUT85), .B(n627), .Z(n630) );
  NAND2_X1 U700 ( .A1(n628), .A2(G87), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U702 ( .A1(G93), .A2(n631), .ZN(n634) );
  NAND2_X1 U703 ( .A1(G80), .A2(n632), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n640) );
  NAND2_X1 U705 ( .A1(G67), .A2(n635), .ZN(n638) );
  NAND2_X1 U706 ( .A1(G55), .A2(n636), .ZN(n637) );
  NAND2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U709 ( .A(KEYINPUT84), .B(n641), .ZN(n832) );
  NOR2_X1 U710 ( .A1(G868), .A2(n832), .ZN(n642) );
  XNOR2_X1 U711 ( .A(n642), .B(KEYINPUT91), .ZN(n654) );
  XNOR2_X1 U712 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n644) );
  XNOR2_X1 U713 ( .A(G305), .B(KEYINPUT19), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U715 ( .A(n645), .B(n832), .ZN(n647) );
  INV_X1 U716 ( .A(G299), .ZN(n702) );
  XNOR2_X1 U717 ( .A(n702), .B(G166), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n648), .B(G290), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n649), .B(G288), .ZN(n836) );
  NAND2_X1 U721 ( .A1(G559), .A2(n943), .ZN(n650) );
  XOR2_X1 U722 ( .A(n937), .B(n650), .Z(n830) );
  XNOR2_X1 U723 ( .A(n836), .B(n830), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n651), .B(KEYINPUT90), .ZN(n652) );
  NAND2_X1 U725 ( .A1(G868), .A2(n652), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(G295) );
  NAND2_X1 U727 ( .A1(G2078), .A2(G2084), .ZN(n655) );
  XOR2_X1 U728 ( .A(KEYINPUT20), .B(n655), .Z(n656) );
  NAND2_X1 U729 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U730 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n658), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U732 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U733 ( .A1(G661), .A2(G483), .ZN(n666) );
  NOR2_X1 U734 ( .A1(G220), .A2(G219), .ZN(n659) );
  XOR2_X1 U735 ( .A(KEYINPUT22), .B(n659), .Z(n660) );
  NOR2_X1 U736 ( .A1(G218), .A2(n660), .ZN(n661) );
  NAND2_X1 U737 ( .A1(G96), .A2(n661), .ZN(n834) );
  NAND2_X1 U738 ( .A1(n834), .A2(G2106), .ZN(n665) );
  NAND2_X1 U739 ( .A1(G69), .A2(G120), .ZN(n662) );
  NOR2_X1 U740 ( .A1(G237), .A2(n662), .ZN(n663) );
  NAND2_X1 U741 ( .A1(G108), .A2(n663), .ZN(n835) );
  NAND2_X1 U742 ( .A1(n835), .A2(G567), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n842) );
  NOR2_X1 U744 ( .A1(n666), .A2(n842), .ZN(n667) );
  XNOR2_X1 U745 ( .A(n667), .B(KEYINPUT92), .ZN(n829) );
  NAND2_X1 U746 ( .A1(G36), .A2(n829), .ZN(G176) );
  NAND2_X1 U747 ( .A1(G126), .A2(n879), .ZN(n669) );
  NAND2_X1 U748 ( .A1(G138), .A2(n883), .ZN(n668) );
  NAND2_X1 U749 ( .A1(n669), .A2(n668), .ZN(n673) );
  NAND2_X1 U750 ( .A1(G114), .A2(n880), .ZN(n671) );
  NAND2_X1 U751 ( .A1(G102), .A2(n884), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U753 ( .A1(n673), .A2(n672), .ZN(G164) );
  NOR2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n933) );
  NOR2_X1 U755 ( .A1(G1971), .A2(G303), .ZN(n674) );
  NOR2_X1 U756 ( .A1(n933), .A2(n674), .ZN(n739) );
  NAND2_X1 U757 ( .A1(G160), .A2(G40), .ZN(n749) );
  XNOR2_X1 U758 ( .A(n749), .B(KEYINPUT97), .ZN(n675) );
  NOR2_X1 U759 ( .A1(G164), .A2(G1384), .ZN(n750) );
  NAND2_X1 U760 ( .A1(n675), .A2(n750), .ZN(n676) );
  XNOR2_X1 U761 ( .A(n676), .B(KEYINPUT64), .ZN(n711) );
  INV_X1 U762 ( .A(n711), .ZN(n691) );
  INV_X2 U763 ( .A(n691), .ZN(n728) );
  NOR2_X1 U764 ( .A1(n728), .A2(G2084), .ZN(n712) );
  NAND2_X1 U765 ( .A1(G8), .A2(n712), .ZN(n726) );
  AND2_X1 U766 ( .A1(n728), .A2(G1961), .ZN(n678) );
  XNOR2_X1 U767 ( .A(G2078), .B(KEYINPUT25), .ZN(n919) );
  NOR2_X1 U768 ( .A1(n728), .A2(n919), .ZN(n677) );
  NOR2_X1 U769 ( .A1(n678), .A2(n677), .ZN(n717) );
  NAND2_X1 U770 ( .A1(n717), .A2(G171), .ZN(n710) );
  NAND2_X1 U771 ( .A1(n728), .A2(G1956), .ZN(n682) );
  INV_X1 U772 ( .A(KEYINPUT27), .ZN(n680) );
  NAND2_X1 U773 ( .A1(G2072), .A2(n691), .ZN(n679) );
  XNOR2_X1 U774 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U775 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U776 ( .A(n683), .B(KEYINPUT98), .Z(n701) );
  NOR2_X1 U777 ( .A1(n702), .A2(n701), .ZN(n684) );
  XOR2_X1 U778 ( .A(n684), .B(KEYINPUT28), .Z(n706) );
  INV_X1 U779 ( .A(G1996), .ZN(n916) );
  NOR2_X1 U780 ( .A1(n711), .A2(n916), .ZN(n686) );
  XNOR2_X1 U781 ( .A(KEYINPUT26), .B(KEYINPUT99), .ZN(n685) );
  XNOR2_X1 U782 ( .A(n686), .B(n685), .ZN(n688) );
  NAND2_X1 U783 ( .A1(n728), .A2(G1341), .ZN(n687) );
  NAND2_X1 U784 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U785 ( .A1(n937), .A2(n689), .ZN(n690) );
  XNOR2_X1 U786 ( .A(KEYINPUT65), .B(n690), .ZN(n697) );
  AND2_X1 U787 ( .A1(n691), .A2(G2067), .ZN(n692) );
  XOR2_X1 U788 ( .A(n692), .B(KEYINPUT100), .Z(n694) );
  NAND2_X1 U789 ( .A1(n728), .A2(G1348), .ZN(n693) );
  NAND2_X1 U790 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U791 ( .A1(n696), .A2(n695), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U793 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U797 ( .A(KEYINPUT29), .B(KEYINPUT101), .ZN(n707) );
  XNOR2_X1 U798 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n722) );
  NAND2_X1 U800 ( .A1(n711), .A2(G8), .ZN(n789) );
  NOR2_X1 U801 ( .A1(G1966), .A2(n789), .ZN(n723) );
  NOR2_X1 U802 ( .A1(n723), .A2(n712), .ZN(n713) );
  XNOR2_X1 U803 ( .A(KEYINPUT102), .B(n713), .ZN(n714) );
  NAND2_X1 U804 ( .A1(n714), .A2(G8), .ZN(n715) );
  XNOR2_X1 U805 ( .A(n715), .B(KEYINPUT30), .ZN(n716) );
  NOR2_X1 U806 ( .A1(n716), .A2(G168), .ZN(n719) );
  NOR2_X1 U807 ( .A1(G171), .A2(n717), .ZN(n718) );
  NOR2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U809 ( .A(KEYINPUT31), .B(n720), .Z(n721) );
  NAND2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n727) );
  INV_X1 U811 ( .A(n727), .ZN(n724) );
  NOR2_X1 U812 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n738) );
  NAND2_X1 U814 ( .A1(n727), .A2(G286), .ZN(n735) );
  INV_X1 U815 ( .A(G8), .ZN(n733) );
  NOR2_X1 U816 ( .A1(n728), .A2(G2090), .ZN(n730) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n789), .ZN(n729) );
  NOR2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U819 ( .A1(n731), .A2(G303), .ZN(n732) );
  OR2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n734) );
  AND2_X1 U821 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U822 ( .A(n736), .B(KEYINPUT32), .ZN(n737) );
  NAND2_X1 U823 ( .A1(n738), .A2(n737), .ZN(n784) );
  NAND2_X1 U824 ( .A1(n739), .A2(n784), .ZN(n740) );
  XNOR2_X1 U825 ( .A(KEYINPUT103), .B(n740), .ZN(n744) );
  NAND2_X1 U826 ( .A1(G288), .A2(G1976), .ZN(n741) );
  XNOR2_X1 U827 ( .A(n741), .B(KEYINPUT104), .ZN(n934) );
  INV_X1 U828 ( .A(n934), .ZN(n742) );
  OR2_X1 U829 ( .A1(n742), .A2(n789), .ZN(n743) );
  NOR2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U831 ( .A1(n745), .A2(KEYINPUT33), .ZN(n748) );
  NAND2_X1 U832 ( .A1(n933), .A2(KEYINPUT33), .ZN(n746) );
  NOR2_X1 U833 ( .A1(n746), .A2(n789), .ZN(n747) );
  NOR2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n780) );
  XOR2_X1 U835 ( .A(G1981), .B(G305), .Z(n948) );
  NOR2_X1 U836 ( .A1(n750), .A2(n749), .ZN(n808) );
  NAND2_X1 U837 ( .A1(G140), .A2(n883), .ZN(n752) );
  NAND2_X1 U838 ( .A1(G104), .A2(n884), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U840 ( .A(KEYINPUT34), .B(n753), .ZN(n759) );
  NAND2_X1 U841 ( .A1(G128), .A2(n879), .ZN(n755) );
  NAND2_X1 U842 ( .A1(G116), .A2(n880), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U844 ( .A(KEYINPUT35), .B(n756), .Z(n757) );
  XNOR2_X1 U845 ( .A(KEYINPUT94), .B(n757), .ZN(n758) );
  NOR2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U847 ( .A(KEYINPUT36), .B(n760), .ZN(n897) );
  XNOR2_X1 U848 ( .A(G2067), .B(KEYINPUT37), .ZN(n805) );
  NOR2_X1 U849 ( .A1(n897), .A2(n805), .ZN(n971) );
  NAND2_X1 U850 ( .A1(n808), .A2(n971), .ZN(n803) );
  NAND2_X1 U851 ( .A1(G129), .A2(n879), .ZN(n762) );
  NAND2_X1 U852 ( .A1(G117), .A2(n880), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n884), .A2(G105), .ZN(n763) );
  XOR2_X1 U855 ( .A(KEYINPUT38), .B(n763), .Z(n764) );
  NOR2_X1 U856 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U857 ( .A(n766), .B(KEYINPUT96), .ZN(n768) );
  NAND2_X1 U858 ( .A1(G141), .A2(n883), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n900) );
  AND2_X1 U860 ( .A1(n900), .A2(G1996), .ZN(n970) );
  NAND2_X1 U861 ( .A1(G119), .A2(n879), .ZN(n770) );
  NAND2_X1 U862 ( .A1(G107), .A2(n880), .ZN(n769) );
  NAND2_X1 U863 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U864 ( .A(KEYINPUT95), .B(n771), .ZN(n775) );
  NAND2_X1 U865 ( .A1(G131), .A2(n883), .ZN(n773) );
  NAND2_X1 U866 ( .A1(G95), .A2(n884), .ZN(n772) );
  AND2_X1 U867 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n896) );
  AND2_X1 U869 ( .A1(n896), .A2(G1991), .ZN(n973) );
  OR2_X1 U870 ( .A1(n970), .A2(n973), .ZN(n776) );
  NAND2_X1 U871 ( .A1(n808), .A2(n776), .ZN(n796) );
  AND2_X1 U872 ( .A1(n803), .A2(n796), .ZN(n791) );
  AND2_X1 U873 ( .A1(n948), .A2(n791), .ZN(n778) );
  XOR2_X1 U874 ( .A(G1986), .B(KEYINPUT93), .Z(n777) );
  XNOR2_X1 U875 ( .A(G290), .B(n777), .ZN(n956) );
  NAND2_X1 U876 ( .A1(n956), .A2(n808), .ZN(n781) );
  AND2_X1 U877 ( .A1(n778), .A2(n781), .ZN(n779) );
  NAND2_X1 U878 ( .A1(n780), .A2(n779), .ZN(n813) );
  INV_X1 U879 ( .A(n781), .ZN(n795) );
  NOR2_X1 U880 ( .A1(G2090), .A2(G303), .ZN(n782) );
  NAND2_X1 U881 ( .A1(G8), .A2(n782), .ZN(n783) );
  NAND2_X1 U882 ( .A1(n784), .A2(n783), .ZN(n786) );
  AND2_X1 U883 ( .A1(n789), .A2(n791), .ZN(n785) );
  AND2_X1 U884 ( .A1(n786), .A2(n785), .ZN(n793) );
  NOR2_X1 U885 ( .A1(G1981), .A2(G305), .ZN(n787) );
  XOR2_X1 U886 ( .A(n787), .B(KEYINPUT24), .Z(n788) );
  NOR2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U889 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U890 ( .A1(n795), .A2(n794), .ZN(n811) );
  NOR2_X1 U891 ( .A1(G1996), .A2(n900), .ZN(n977) );
  INV_X1 U892 ( .A(n796), .ZN(n800) );
  NOR2_X1 U893 ( .A1(G1991), .A2(n896), .ZN(n797) );
  XOR2_X1 U894 ( .A(KEYINPUT105), .B(n797), .Z(n967) );
  NOR2_X1 U895 ( .A1(G1986), .A2(G290), .ZN(n798) );
  NOR2_X1 U896 ( .A1(n967), .A2(n798), .ZN(n799) );
  NOR2_X1 U897 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U898 ( .A1(n977), .A2(n801), .ZN(n802) );
  XNOR2_X1 U899 ( .A(n802), .B(KEYINPUT39), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n897), .A2(n805), .ZN(n969) );
  NAND2_X1 U902 ( .A1(n806), .A2(n969), .ZN(n807) );
  XNOR2_X1 U903 ( .A(KEYINPUT106), .B(n807), .ZN(n809) );
  AND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U907 ( .A(n814), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U908 ( .A(G2454), .B(G2430), .Z(n816) );
  XNOR2_X1 U909 ( .A(G2451), .B(G2446), .ZN(n815) );
  XNOR2_X1 U910 ( .A(n816), .B(n815), .ZN(n823) );
  XOR2_X1 U911 ( .A(G2443), .B(G2427), .Z(n818) );
  XNOR2_X1 U912 ( .A(G2438), .B(KEYINPUT107), .ZN(n817) );
  XNOR2_X1 U913 ( .A(n818), .B(n817), .ZN(n819) );
  XOR2_X1 U914 ( .A(n819), .B(G2435), .Z(n821) );
  XNOR2_X1 U915 ( .A(G1348), .B(G1341), .ZN(n820) );
  XNOR2_X1 U916 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n824), .A2(G14), .ZN(n904) );
  XOR2_X1 U919 ( .A(KEYINPUT108), .B(n904), .Z(G401) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n825), .ZN(G217) );
  NAND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n826) );
  XNOR2_X1 U922 ( .A(KEYINPUT109), .B(n826), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n827), .A2(G661), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(G188) );
  XNOR2_X1 U927 ( .A(KEYINPUT83), .B(n830), .ZN(n831) );
  NOR2_X1 U928 ( .A1(G860), .A2(n831), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(G145) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U935 ( .A(G286), .B(n836), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n943), .B(G171), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n840) );
  XOR2_X1 U938 ( .A(n937), .B(KEYINPUT115), .Z(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n841) );
  NOR2_X1 U940 ( .A1(G37), .A2(n841), .ZN(G397) );
  INV_X1 U941 ( .A(n842), .ZN(G319) );
  XOR2_X1 U942 ( .A(G2096), .B(KEYINPUT43), .Z(n844) );
  XNOR2_X1 U943 ( .A(G2072), .B(KEYINPUT110), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U945 ( .A(n845), .B(KEYINPUT42), .Z(n847) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2090), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U948 ( .A(G2678), .B(G2100), .Z(n849) );
  XNOR2_X1 U949 ( .A(G2078), .B(G2084), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U952 ( .A(KEYINPUT41), .B(G1981), .Z(n853) );
  XNOR2_X1 U953 ( .A(G1966), .B(G1956), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(n854), .B(KEYINPUT112), .Z(n856) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U958 ( .A(G1976), .B(G1971), .Z(n858) );
  XNOR2_X1 U959 ( .A(G1986), .B(G1961), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U961 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U962 ( .A(KEYINPUT111), .B(G2474), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G136), .A2(n883), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G112), .A2(n880), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n869) );
  NAND2_X1 U967 ( .A1(n879), .A2(G124), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G100), .A2(n884), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U971 ( .A1(n869), .A2(n868), .ZN(G162) );
  NAND2_X1 U972 ( .A1(G139), .A2(n883), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G103), .A2(n884), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G127), .A2(n879), .ZN(n873) );
  NAND2_X1 U976 ( .A1(G115), .A2(n880), .ZN(n872) );
  NAND2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n874), .Z(n875) );
  NOR2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n963) );
  XOR2_X1 U980 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n878) );
  XNOR2_X1 U981 ( .A(G164), .B(KEYINPUT48), .ZN(n877) );
  XNOR2_X1 U982 ( .A(n878), .B(n877), .ZN(n892) );
  NAND2_X1 U983 ( .A1(G130), .A2(n879), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G118), .A2(n880), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G142), .A2(n883), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G106), .A2(n884), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U989 ( .A(KEYINPUT45), .B(n887), .ZN(n888) );
  XNOR2_X1 U990 ( .A(KEYINPUT113), .B(n888), .ZN(n889) );
  NOR2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U992 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U993 ( .A(G160), .B(G162), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n963), .B(n895), .ZN(n899) );
  XOR2_X1 U996 ( .A(n897), .B(n896), .Z(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n974), .B(n900), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n903), .ZN(G395) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n904), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(KEYINPUT116), .B(n905), .ZN(n906) );
  NOR2_X1 U1003 ( .A1(G397), .A2(n906), .ZN(n909) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n907) );
  XOR2_X1 U1005 ( .A(KEYINPUT49), .B(n907), .Z(n908) );
  NAND2_X1 U1006 ( .A1(n909), .A2(n908), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(n910), .A2(G395), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n911), .B(KEYINPUT117), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1011 ( .A(G2072), .B(G33), .Z(n912) );
  NAND2_X1 U1012 ( .A1(n912), .A2(G28), .ZN(n915) );
  XOR2_X1 U1013 ( .A(G26), .B(G2067), .Z(n913) );
  XNOR2_X1 U1014 ( .A(KEYINPUT119), .B(n913), .ZN(n914) );
  NOR2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n923) );
  XOR2_X1 U1016 ( .A(G1991), .B(G25), .Z(n918) );
  XNOR2_X1 U1017 ( .A(n916), .B(G32), .ZN(n917) );
  NAND2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n921) );
  XOR2_X1 U1019 ( .A(G27), .B(n919), .Z(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(n924), .B(KEYINPUT53), .ZN(n927) );
  XOR2_X1 U1023 ( .A(G2084), .B(G34), .Z(n925) );
  XNOR2_X1 U1024 ( .A(KEYINPUT54), .B(n925), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(G35), .B(G2090), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(n930), .B(KEYINPUT120), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(G29), .A2(n931), .ZN(n932) );
  XOR2_X1 U1030 ( .A(KEYINPUT55), .B(n932), .Z(n962) );
  XOR2_X1 U1031 ( .A(G16), .B(KEYINPUT56), .Z(n959) );
  INV_X1 U1032 ( .A(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(n936), .B(KEYINPUT121), .ZN(n954) );
  XNOR2_X1 U1035 ( .A(G1341), .B(KEYINPUT122), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(n938), .B(n937), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(G1956), .B(G299), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(G166), .B(G1971), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G171), .B(G1961), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1042 ( .A(G1348), .B(n943), .Z(n944) );
  NOR2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G1966), .B(G168), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1047 ( .A(KEYINPUT57), .B(n950), .Z(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1051 ( .A(KEYINPUT123), .B(n957), .Z(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(KEYINPUT124), .B(n960), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n991) );
  XOR2_X1 U1055 ( .A(G2072), .B(n963), .Z(n965) );
  XOR2_X1 U1056 ( .A(G164), .B(G2078), .Z(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(KEYINPUT50), .B(n966), .ZN(n987) );
  INV_X1 U1059 ( .A(n967), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n984) );
  NOR2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n982) );
  XOR2_X1 U1062 ( .A(G160), .B(G2084), .Z(n972) );
  NOR2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n975) );
  NAND2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n980) );
  XOR2_X1 U1065 ( .A(G2090), .B(G162), .Z(n976) );
  NOR2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(n978), .B(KEYINPUT51), .ZN(n979) );
  NOR2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1069 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1070 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1071 ( .A(KEYINPUT118), .B(n985), .ZN(n986) );
  NAND2_X1 U1072 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(KEYINPUT52), .B(n988), .ZN(n989) );
  NAND2_X1 U1074 ( .A1(n989), .A2(G29), .ZN(n990) );
  NAND2_X1 U1075 ( .A1(n991), .A2(n990), .ZN(n1018) );
  XOR2_X1 U1076 ( .A(G1986), .B(G24), .Z(n995) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n993) );
  XNOR2_X1 U1078 ( .A(G23), .B(G1976), .ZN(n992) );
  NOR2_X1 U1079 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1080 ( .A1(n995), .A2(n994), .ZN(n997) );
  XNOR2_X1 U1081 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(n997), .B(n996), .ZN(n1001) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G21), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(G5), .B(G1961), .ZN(n998) );
  NOR2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1011) );
  XOR2_X1 U1087 ( .A(G1348), .B(KEYINPUT59), .Z(n1002) );
  XNOR2_X1 U1088 ( .A(G4), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(G20), .B(G1956), .ZN(n1003) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(G1341), .B(G19), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G1981), .B(G6), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(KEYINPUT60), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(KEYINPUT126), .B(n1012), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(n1013), .B(KEYINPUT61), .ZN(n1015) );
  INV_X1 U1099 ( .A(G16), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1101 ( .A1(G11), .A2(n1016), .ZN(n1017) );
  NOR2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(n1019), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

