//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G128), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G110), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(new_n191), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT24), .B(G110), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n194), .A2(new_n195), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n199), .B(KEYINPUT76), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n205));
  OR3_X1    g019(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G146), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n202), .A2(new_n204), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n200), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(G146), .B1(new_n205), .B2(new_n206), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  OAI221_X1 g028(.A(new_n214), .B1(new_n195), .B2(new_n194), .C1(new_n197), .C2(new_n198), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT22), .B(G137), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n216), .B(KEYINPUT77), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT71), .A2(G953), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT71), .A2(G953), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(G221), .A3(G234), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n217), .B(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n211), .A2(new_n215), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n211), .A2(new_n215), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n222), .B(KEYINPUT78), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n187), .B(new_n223), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n226), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n224), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n231), .A2(KEYINPUT25), .A3(new_n187), .A4(new_n223), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G217), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(G234), .B2(new_n187), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n223), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n235), .A2(G902), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n233), .A2(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT74), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT11), .A2(G134), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT67), .B1(new_n242), .B2(G137), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT11), .A4(G134), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  AOI21_X1  g062(.A(G131), .B1(new_n248), .B2(G137), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(G134), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT11), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT66), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI211_X1 g066(.A(KEYINPUT66), .B(new_n251), .C1(new_n248), .C2(G137), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n247), .B(new_n249), .C1(new_n252), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n248), .A2(G137), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n250), .A3(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n258), .B(G131), .C1(new_n257), .C2(new_n256), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n259), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT65), .B1(new_n265), .B2(G146), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT64), .B(G143), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(G146), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(KEYINPUT64), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT64), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G143), .ZN(new_n272));
  AND4_X1   g086(.A1(new_n269), .A2(new_n270), .A3(new_n272), .A4(G146), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n264), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT1), .B1(new_n265), .B2(G146), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G128), .ZN(new_n276));
  AOI21_X1  g090(.A(G146), .B1(new_n270), .B2(new_n272), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n209), .A2(G143), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n262), .A2(new_n263), .A3(new_n280), .ZN(new_n281));
  OR2_X1    g095(.A1(new_n189), .A2(G116), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n189), .A2(G116), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT2), .B(G113), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n247), .B(new_n256), .C1(new_n252), .C2(new_n254), .ZN(new_n288));
  NAND2_X1  g102(.A1(KEYINPUT68), .A2(G131), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n251), .B1(new_n248), .B2(G137), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n294), .A2(new_n253), .B1(new_n243), .B2(new_n246), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n256), .A3(new_n289), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n270), .A2(new_n272), .A3(G146), .ZN(new_n298));
  INV_X1    g112(.A(new_n266), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n267), .A2(new_n269), .A3(G146), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g116(.A1(KEYINPUT0), .A2(G128), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n270), .A2(new_n272), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n209), .ZN(new_n305));
  INV_X1    g119(.A(new_n278), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(KEYINPUT0), .A2(G128), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n302), .A2(new_n303), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n297), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n281), .A2(new_n287), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G237), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n220), .A2(G210), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT27), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT27), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n220), .A2(new_n316), .A3(G210), .A4(new_n313), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT26), .B(G101), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n315), .B2(new_n317), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n280), .A2(new_n255), .A3(new_n259), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n311), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n260), .A2(new_n261), .B1(new_n274), .B2(new_n279), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n326), .A2(new_n263), .B1(new_n297), .B2(new_n310), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n327), .B2(new_n324), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n322), .B1(new_n328), .B2(new_n286), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT31), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n287), .B1(new_n311), .B2(new_n323), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n312), .A2(KEYINPUT28), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n281), .A2(new_n311), .A3(new_n333), .A4(new_n287), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI22_X1  g149(.A1(new_n329), .A2(new_n330), .B1(new_n335), .B2(new_n321), .ZN(new_n336));
  INV_X1    g150(.A(new_n325), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n324), .B1(new_n281), .B2(new_n311), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n286), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n322), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n330), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n329), .A2(KEYINPUT72), .A3(new_n330), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n336), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(G472), .A2(G902), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n346), .B(KEYINPUT73), .Z(new_n347));
  OAI21_X1  g161(.A(new_n241), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT32), .ZN(new_n349));
  INV_X1    g163(.A(new_n347), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT72), .B1(new_n329), .B2(new_n330), .ZN(new_n351));
  AND4_X1   g165(.A1(KEYINPUT72), .A2(new_n339), .A3(new_n330), .A4(new_n340), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(KEYINPUT74), .B(new_n350), .C1(new_n353), .C2(new_n336), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n348), .A2(new_n349), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n343), .A2(new_n344), .ZN(new_n356));
  INV_X1    g170(.A(new_n336), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n347), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n335), .A2(new_n321), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n360));
  INV_X1    g174(.A(new_n312), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n328), .B2(new_n286), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n359), .B(new_n360), .C1(new_n321), .C2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT75), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n287), .B1(new_n281), .B2(new_n311), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n321), .A2(KEYINPUT29), .ZN(new_n366));
  AOI211_X1 g180(.A(new_n365), .B(new_n366), .C1(new_n332), .C2(new_n334), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n364), .B1(new_n367), .B2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n332), .A2(new_n334), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n327), .A2(new_n287), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT75), .B(new_n187), .C1(new_n371), .C2(new_n366), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n363), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n358), .A2(KEYINPUT32), .B1(new_n373), .B2(G472), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n240), .B1(new_n355), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G140), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT79), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n220), .A2(G227), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G107), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n381), .A2(G107), .ZN(new_n384));
  OAI21_X1  g198(.A(G101), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(new_n381), .B2(G107), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G104), .ZN(new_n389));
  INV_X1    g203(.A(G101), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n386), .A2(new_n389), .A3(new_n390), .A4(new_n382), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n280), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n192), .B1(new_n305), .B2(KEYINPUT1), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT82), .B1(new_n395), .B2(new_n302), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT1), .ZN(new_n397));
  OAI21_X1  g211(.A(G128), .B1(new_n277), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n398), .A2(new_n399), .A3(new_n300), .A4(new_n301), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n274), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n394), .B1(new_n401), .B2(new_n393), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n297), .A2(KEYINPUT83), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT12), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT12), .ZN(new_n405));
  INV_X1    g219(.A(new_n403), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n398), .A2(new_n300), .A3(new_n301), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n407), .A2(KEYINPUT82), .B1(new_n302), .B2(new_n264), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n392), .B1(new_n408), .B2(new_n400), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n405), .B(new_n406), .C1(new_n409), .C2(new_n394), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT10), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n401), .A2(new_n412), .A3(new_n393), .ZN(new_n413));
  INV_X1    g227(.A(new_n280), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT10), .B1(new_n414), .B2(new_n392), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n297), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n302), .A2(new_n303), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n307), .A2(new_n309), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n386), .A2(new_n389), .A3(new_n382), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G101), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n425), .A3(G101), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT80), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n418), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n426), .B(KEYINPUT80), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n430), .A2(KEYINPUT81), .A3(new_n310), .A4(new_n423), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n416), .A2(new_n417), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT84), .B1(new_n411), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n433), .A2(KEYINPUT84), .A3(new_n404), .A4(new_n410), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n380), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n380), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n413), .A2(new_n415), .B1(new_n429), .B2(new_n431), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n441), .B2(new_n417), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n416), .A2(new_n432), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT85), .A3(new_n297), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n439), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n437), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G469), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n376), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n404), .A2(new_n410), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n416), .A2(new_n417), .A3(new_n432), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n435), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n445), .B1(new_n454), .B2(new_n380), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT86), .B(G469), .C1(new_n455), .C2(G902), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n442), .A2(new_n444), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n438), .B1(new_n457), .B2(new_n433), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n439), .A2(new_n451), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n448), .B(new_n187), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n449), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT9), .B(G234), .ZN(new_n462));
  OAI21_X1  g276(.A(G221), .B1(new_n462), .B2(G902), .ZN(new_n463));
  OAI21_X1  g277(.A(G210), .B1(G237), .B2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n310), .A2(new_n203), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n414), .A2(new_n203), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G224), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n469), .A2(G953), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n468), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n286), .A2(new_n423), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT88), .B1(new_n428), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n430), .A2(new_n474), .A3(new_n286), .A4(new_n423), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n283), .A2(KEYINPUT5), .ZN(new_n476));
  INV_X1    g290(.A(G113), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n283), .A2(new_n282), .A3(KEYINPUT5), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n284), .A2(new_n285), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n393), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(G110), .B(G122), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n473), .A2(new_n475), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT6), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n473), .A2(new_n475), .A3(new_n482), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n483), .B(KEYINPUT89), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(KEYINPUT6), .A3(new_n487), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n471), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n481), .A2(new_n480), .A3(new_n392), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n483), .B(KEYINPUT8), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n478), .A2(KEYINPUT90), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n478), .A2(KEYINPUT90), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n479), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n481), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n494), .B1(new_n393), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n310), .A2(new_n203), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n280), .A2(G125), .ZN(new_n501));
  OAI211_X1 g315(.A(KEYINPUT7), .B(new_n470), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n470), .A2(KEYINPUT7), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n466), .A2(new_n467), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n499), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n484), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n187), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n465), .B1(new_n491), .B2(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n468), .B(new_n470), .Z(new_n509));
  AOI22_X1  g323(.A1(new_n484), .A2(KEYINPUT6), .B1(new_n486), .B2(new_n487), .ZN(new_n510));
  INV_X1    g324(.A(new_n490), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(G902), .B1(new_n505), .B2(new_n484), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n464), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT18), .A2(G131), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n220), .A2(G143), .A3(G214), .A4(new_n313), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n218), .A2(G214), .A3(new_n313), .A4(new_n219), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n267), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n208), .B(G146), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n516), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n519), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G131), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n517), .B2(new_n519), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT17), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n213), .A2(KEYINPUT91), .A3(new_n207), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT91), .ZN(new_n530));
  INV_X1    g344(.A(new_n207), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(new_n212), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n517), .A2(new_n526), .A3(new_n519), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n534), .A2(new_n527), .A3(KEYINPUT17), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n525), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(G113), .B(G122), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n381), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT92), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n525), .B(new_n539), .C1(new_n533), .C2(new_n535), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n187), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G475), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n208), .B(KEYINPUT19), .Z(new_n545));
  OAI221_X1 g359(.A(new_n207), .B1(new_n545), .B2(G146), .C1(new_n527), .C2(new_n534), .ZN(new_n546));
  INV_X1    g360(.A(new_n538), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n525), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(G475), .A2(G902), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n524), .A2(new_n523), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n550), .A2(new_n520), .A3(new_n521), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n552));
  OR3_X1    g366(.A1(new_n534), .A2(new_n527), .A3(KEYINPUT17), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n548), .B(new_n549), .C1(new_n554), .C2(new_n547), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n536), .A2(new_n538), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n558), .A2(KEYINPUT20), .A3(new_n548), .A4(new_n549), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n544), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n267), .A2(G128), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n192), .A2(G143), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n248), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(G116), .B(G122), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(new_n388), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n561), .A2(new_n566), .A3(new_n562), .ZN(new_n567));
  OAI21_X1  g381(.A(G134), .B1(new_n561), .B2(new_n566), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n563), .B(new_n565), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G122), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G116), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n388), .B1(new_n571), .B2(KEYINPUT14), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(new_n564), .ZN(new_n573));
  INV_X1    g387(.A(new_n563), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n248), .B1(new_n561), .B2(new_n562), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n462), .A2(new_n234), .A3(G953), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n569), .A2(new_n576), .A3(new_n578), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n577), .A2(KEYINPUT94), .A3(new_n579), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n187), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G478), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(KEYINPUT15), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n587), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n583), .A2(new_n187), .A3(new_n584), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G952), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(G953), .ZN(new_n593));
  INV_X1    g407(.A(G234), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n593), .B1(new_n594), .B2(new_n313), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n187), .B(new_n220), .C1(G234), .C2(G237), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT21), .B(G898), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n560), .A2(new_n591), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(G214), .B1(G237), .B2(G902), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT87), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n515), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n375), .A2(new_n461), .A3(new_n463), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  AND2_X1   g419(.A1(new_n461), .A2(new_n463), .ZN(new_n606));
  OAI21_X1  g420(.A(G472), .B1(new_n345), .B2(G902), .ZN(new_n607));
  AND4_X1   g421(.A1(new_n348), .A2(new_n607), .A3(new_n354), .A4(new_n239), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n515), .A2(new_n601), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n585), .A2(new_n586), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n577), .A2(KEYINPUT95), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n579), .A2(KEYINPUT96), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n582), .B2(KEYINPUT96), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n612), .A2(new_n613), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n583), .A2(new_n615), .A3(new_n584), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n187), .A2(G478), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n611), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n560), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n610), .A2(new_n599), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n609), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  NAND4_X1  g441(.A1(new_n591), .A2(new_n559), .A3(new_n544), .A4(new_n557), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n610), .A2(new_n599), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n609), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT98), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NAND2_X1  g448(.A1(new_n233), .A2(new_n235), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT36), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n226), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(new_n224), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n238), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  AND4_X1   g455(.A1(new_n348), .A2(new_n607), .A3(new_n354), .A4(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n461), .A2(new_n463), .A3(new_n603), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  NAND2_X1  g459(.A1(new_n355), .A2(new_n374), .ZN(new_n646));
  INV_X1    g460(.A(new_n641), .ZN(new_n647));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n596), .B1(new_n597), .B2(new_n648), .ZN(new_n649));
  NOR4_X1   g463(.A1(new_n647), .A2(new_n610), .A3(new_n628), .A4(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n606), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  XOR2_X1   g466(.A(new_n649), .B(KEYINPUT39), .Z(new_n653));
  NAND2_X1  g467(.A1(new_n606), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n358), .A2(KEYINPUT32), .ZN(new_n657));
  INV_X1    g471(.A(G472), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n339), .A2(new_n340), .ZN(new_n659));
  INV_X1    g473(.A(new_n321), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n660), .B1(new_n361), .B2(new_n365), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n355), .B(new_n657), .C1(new_n658), .C2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n515), .B(KEYINPUT38), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n560), .A2(new_n601), .A3(new_n591), .ZN(new_n665));
  AND4_X1   g479(.A1(new_n647), .A2(new_n663), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n655), .A2(new_n656), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n304), .ZN(G45));
  OR2_X1    g482(.A1(new_n623), .A2(new_n649), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n610), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT99), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n647), .B1(new_n355), .B2(new_n374), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n606), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  AOI21_X1  g488(.A(KEYINPUT85), .B1(new_n443), .B2(new_n297), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n441), .A2(new_n440), .A3(new_n417), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n433), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n459), .B1(new_n677), .B2(new_n380), .ZN(new_n678));
  OAI21_X1  g492(.A(G469), .B1(new_n678), .B2(G902), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n463), .A3(new_n460), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n679), .A2(KEYINPUT100), .A3(new_n463), .A4(new_n460), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n375), .A2(new_n624), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NAND2_X1  g500(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n688), .A2(KEYINPUT101), .A3(new_n375), .A4(new_n629), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n375), .A2(new_n629), .A3(new_n682), .A4(new_n683), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  NAND4_X1  g508(.A1(new_n682), .A2(new_n515), .A3(new_n601), .A4(new_n683), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n672), .A2(new_n600), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n189), .ZN(G21));
  NAND2_X1  g512(.A1(new_n665), .A2(new_n515), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n665), .A2(new_n515), .A3(KEYINPUT102), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n599), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n356), .A2(new_n357), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n658), .B1(new_n704), .B2(new_n187), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n660), .A2(new_n371), .B1(new_n659), .B2(KEYINPUT31), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n347), .B1(new_n356), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n705), .A2(new_n240), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n703), .A2(new_n682), .A3(new_n683), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G122), .ZN(G24));
  INV_X1    g524(.A(new_n695), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n647), .A2(new_n705), .A3(new_n707), .ZN(new_n712));
  INV_X1    g526(.A(new_n669), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  INV_X1    g530(.A(new_n463), .ZN(new_n717));
  OAI21_X1  g531(.A(G469), .B1(new_n455), .B2(G902), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n717), .B1(new_n718), .B2(new_n460), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n508), .A2(new_n514), .A3(new_n601), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT103), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n508), .A2(new_n514), .A3(new_n722), .A4(new_n601), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n719), .A2(new_n724), .A3(new_n713), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n726), .B1(new_n358), .B2(KEYINPUT32), .ZN(new_n727));
  OAI211_X1 g541(.A(KEYINPUT104), .B(new_n349), .C1(new_n345), .C2(new_n347), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n374), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n239), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT42), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n669), .A2(KEYINPUT42), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n375), .A2(new_n724), .A3(new_n719), .A4(new_n732), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G131), .ZN(G33));
  NOR2_X1   g549(.A1(new_n628), .A2(new_n649), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n375), .A2(new_n736), .A3(new_n724), .A4(new_n719), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT105), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n719), .A2(new_n724), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n375), .A4(new_n736), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NAND2_X1  g557(.A1(G469), .A2(G902), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n455), .A2(KEYINPUT45), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT106), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n455), .A2(new_n747), .A3(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n455), .A2(KEYINPUT45), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n448), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n750), .B1(new_n749), .B2(new_n752), .ZN(new_n755));
  OAI211_X1 g569(.A(KEYINPUT46), .B(new_n744), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n744), .B1(new_n754), .B2(new_n755), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n749), .A2(new_n752), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT107), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n753), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(KEYINPUT108), .A3(KEYINPUT46), .A4(new_n744), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n758), .A2(new_n761), .A3(new_n765), .A4(new_n460), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n766), .A2(new_n463), .A3(new_n653), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n348), .A2(new_n607), .A3(new_n354), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n641), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(KEYINPUT109), .Z(new_n770));
  NAND4_X1  g584(.A1(new_n622), .A2(new_n559), .A3(new_n544), .A4(new_n557), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT43), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(KEYINPUT44), .ZN(new_n774));
  INV_X1    g588(.A(new_n724), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n773), .B2(KEYINPUT44), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n767), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  NAND2_X1  g592(.A1(new_n766), .A2(new_n463), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT47), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n775), .A2(new_n646), .A3(new_n239), .A4(new_n669), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n201), .ZN(G42));
  NAND3_X1  g598(.A1(new_n239), .A2(new_n463), .A3(new_n602), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT110), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n679), .A2(new_n460), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n771), .B(new_n786), .C1(KEYINPUT49), .C2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT111), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(KEYINPUT49), .ZN(new_n790));
  OR4_X1    g604(.A1(new_n663), .A2(new_n789), .A3(new_n664), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n690), .B(KEYINPUT101), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n709), .B(new_n684), .C1(new_n695), .C2(new_n696), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n793), .A2(KEYINPUT112), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n796));
  INV_X1    g610(.A(new_n794), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n796), .B1(new_n797), .B2(new_n693), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n623), .A2(new_n628), .ZN(new_n800));
  INV_X1    g614(.A(new_n599), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n515), .A2(new_n800), .A3(new_n602), .A4(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n461), .A2(new_n463), .A3(new_n802), .A4(new_n608), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n604), .A2(new_n643), .A3(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n560), .A2(new_n591), .A3(new_n649), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n721), .A2(new_n723), .A3(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n461), .A2(new_n463), .A3(new_n806), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n807), .A2(new_n672), .B1(new_n714), .B2(new_n739), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n734), .A2(new_n742), .A3(new_n804), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT113), .B1(new_n799), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT112), .B1(new_n793), .B2(new_n794), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n797), .A2(new_n693), .A3(new_n796), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(new_n811), .A3(KEYINPUT113), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n649), .B1(new_n701), .B2(new_n702), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n663), .A2(new_n814), .A3(new_n647), .A4(new_n719), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n715), .A2(new_n673), .A3(new_n651), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n792), .B1(new_n810), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n793), .A2(new_n792), .A3(new_n794), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n818), .A2(new_n809), .A3(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n826), .B(new_n792), .C1(new_n810), .C2(new_n819), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n810), .A2(new_n819), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n825), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n824), .B1(new_n830), .B2(KEYINPUT54), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n687), .A2(new_n775), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n833), .A2(new_n240), .A3(new_n595), .A4(new_n663), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n622), .A2(new_n560), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n772), .A2(new_n595), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n834), .A2(new_n835), .B1(new_n712), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n708), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n840), .A2(new_n687), .A3(new_n601), .A4(new_n664), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT50), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT118), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n787), .B(KEYINPUT116), .Z(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n463), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT117), .Z(new_n846));
  AND2_X1   g660(.A1(new_n780), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n840), .A2(new_n775), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n839), .B(new_n843), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n837), .A2(new_n730), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT119), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT48), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT120), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n855), .A2(KEYINPUT120), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n834), .A2(new_n560), .A3(new_n622), .ZN(new_n859));
  INV_X1    g673(.A(new_n840), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n592), .B(G953), .C1(new_n711), .C2(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n859), .B(new_n861), .C1(new_n854), .C2(new_n856), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n779), .B(KEYINPUT47), .Z(new_n863));
  OAI21_X1  g677(.A(new_n848), .B1(new_n863), .B2(new_n845), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n839), .A2(KEYINPUT51), .A3(new_n842), .ZN(new_n865));
  AOI211_X1 g679(.A(new_n858), .B(new_n862), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n831), .A2(new_n852), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(G952), .A2(G953), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n791), .B1(new_n867), .B2(new_n868), .ZN(G75));
  NOR2_X1   g683(.A1(new_n220), .A2(G952), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n187), .B1(new_n820), .B2(new_n823), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(G210), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n510), .A2(new_n511), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n471), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n512), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT55), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n871), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n875), .A2(new_n879), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT121), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n875), .A2(new_n883), .A3(new_n879), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n880), .B1(new_n882), .B2(new_n884), .ZN(G51));
  AOI21_X1  g699(.A(new_n821), .B1(new_n820), .B2(new_n823), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n824), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n744), .B(KEYINPUT57), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n887), .A2(new_n888), .B1(new_n458), .B2(new_n459), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n872), .A2(new_n753), .A3(new_n763), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n870), .B1(new_n889), .B2(new_n890), .ZN(G54));
  NAND3_X1  g705(.A1(new_n872), .A2(KEYINPUT58), .A3(G475), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n558), .A2(new_n548), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n870), .ZN(G60));
  XNOR2_X1  g710(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n897));
  NAND2_X1  g711(.A1(G478), .A2(G902), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n620), .B1(new_n831), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n620), .A2(new_n899), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n820), .A2(new_n823), .ZN(new_n904));
  INV_X1    g718(.A(new_n821), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n901), .B1(new_n908), .B2(new_n870), .ZN(new_n909));
  OAI211_X1 g723(.A(KEYINPUT123), .B(new_n871), .C1(new_n887), .C2(new_n903), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n900), .A2(new_n909), .A3(new_n910), .ZN(G63));
  AND2_X1   g725(.A1(new_n820), .A2(new_n823), .ZN(new_n912));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT60), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n912), .A2(new_n638), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n236), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n871), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n915), .A2(KEYINPUT61), .A3(new_n871), .A4(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(G66));
  OAI21_X1  g735(.A(G953), .B1(new_n598), .B2(new_n469), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n799), .A2(new_n804), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n220), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n876), .B1(G898), .B2(new_n220), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT124), .Z(new_n928));
  XNOR2_X1  g742(.A(new_n926), .B(new_n928), .ZN(G69));
  INV_X1    g743(.A(G227), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n925), .B1(new_n930), .B2(new_n648), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n328), .B(new_n545), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n925), .A2(new_n648), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT125), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n730), .B1(new_n701), .B2(new_n702), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n767), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n715), .A2(new_n673), .A3(new_n651), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n942), .A2(new_n734), .A3(new_n742), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n777), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n783), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n939), .B1(new_n945), .B2(new_n220), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n667), .A2(new_n942), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n667), .A2(KEYINPUT62), .A3(new_n942), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n375), .A2(new_n724), .A3(new_n800), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n654), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n777), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n220), .B(new_n935), .C1(new_n783), .C2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n933), .B(new_n934), .C1(new_n946), .C2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n783), .A2(new_n944), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n936), .B(new_n938), .C1(new_n958), .C2(new_n925), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n959), .A2(new_n932), .A3(new_n931), .A4(new_n955), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n957), .A2(new_n960), .ZN(G72));
  XNOR2_X1  g775(.A(new_n362), .B(KEYINPUT127), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n783), .A2(new_n954), .A3(new_n923), .ZN(new_n963));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT63), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n321), .B(new_n962), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n962), .A2(new_n321), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n783), .A2(new_n944), .A3(new_n923), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n965), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n871), .A3(new_n969), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n362), .A2(new_n321), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n965), .B1(new_n971), .B2(new_n659), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n830), .B2(new_n972), .ZN(G57));
endmodule


