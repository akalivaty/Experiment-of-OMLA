//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT81), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G15gat), .B(G22gat), .Z(new_n210));
  INV_X1    g009(.A(G1gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(G1gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n215), .A3(KEYINPUT86), .ZN(new_n216));
  INV_X1    g015(.A(G8gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT85), .ZN(new_n219));
  INV_X1    g018(.A(G43gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G50gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT84), .B(G43gat), .ZN(new_n223));
  INV_X1    g022(.A(G50gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n219), .B1(new_n225), .B2(KEYINPUT15), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n220), .A2(KEYINPUT84), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT84), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G43gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n229), .A3(new_n224), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n221), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT15), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(KEYINPUT85), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G29gat), .ZN(new_n234));
  INV_X1    g033(.A(G36gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT14), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT14), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(G29gat), .B2(G36gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(G29gat), .A2(G36gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT15), .B1(new_n224), .B2(G43gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n220), .A2(G50gat), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT83), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n224), .A2(G43gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT83), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n221), .A2(new_n244), .A3(new_n245), .A4(KEYINPUT15), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n240), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n226), .A2(new_n233), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n241), .A2(new_n242), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n240), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n240), .A2(new_n250), .A3(KEYINPUT82), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n248), .A2(new_n249), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n249), .B1(new_n248), .B2(new_n255), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n218), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G229gat), .A2(G233gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n216), .B(G8gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n248), .A2(new_n255), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT88), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n258), .A2(KEYINPUT18), .A3(new_n259), .A4(new_n262), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n267), .A2(KEYINPUT89), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(KEYINPUT89), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT88), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n263), .A2(new_n271), .A3(new_n264), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n218), .A2(new_n248), .A3(new_n255), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n262), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT13), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n209), .B1(new_n270), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n260), .A2(new_n261), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n261), .A2(KEYINPUT17), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n248), .A2(new_n249), .A3(new_n255), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n280), .B1(new_n283), .B2(new_n218), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT89), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT18), .A4(new_n259), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n267), .A2(KEYINPUT89), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n207), .B1(new_n274), .B2(new_n276), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n265), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n279), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G141gat), .B(G148gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT2), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n294), .B1(G155gat), .B2(G162gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT70), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G155gat), .B(G162gat), .Z(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n296), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT3), .ZN(new_n300));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(KEYINPUT1), .ZN(new_n302));
  XNOR2_X1  g101(.A(G127gat), .B(G134gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n296), .A2(new_n297), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n296), .A2(new_n297), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n300), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310));
  INV_X1    g109(.A(new_n304), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n296), .B(new_n297), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n299), .A2(new_n304), .A3(KEYINPUT4), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G225gat), .A2(G233gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n299), .B(new_n304), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n318), .B(KEYINPUT39), .C1(new_n317), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT39), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n315), .A2(new_n321), .A3(new_n317), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n323));
  XOR2_X1   g122(.A(G1gat), .B(G29gat), .Z(new_n324));
  XNOR2_X1  g123(.A(G57gat), .B(G85gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT71), .B(KEYINPUT0), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n326), .B(new_n327), .Z(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n322), .A2(new_n323), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n323), .B1(new_n322), .B2(new_n329), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n320), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT40), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT22), .ZN(new_n335));
  INV_X1    g134(.A(G211gat), .ZN(new_n336));
  INV_X1    g135(.A(G218gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G211gat), .B(G218gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n341), .B(KEYINPUT67), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n344));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n345), .A2(KEYINPUT24), .ZN(new_n346));
  INV_X1    g145(.A(G183gat), .ZN(new_n347));
  INV_X1    g146(.A(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n346), .A2(new_n349), .B1(G169gat), .B2(G176gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n350), .B(new_n353), .C1(KEYINPUT24), .C2(new_n345), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT27), .B1(new_n347), .B2(KEYINPUT64), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT27), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G183gat), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n357), .B(new_n348), .C1(KEYINPUT64), .C2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT27), .B(G183gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(KEYINPUT28), .A3(new_n348), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n362), .A2(new_n364), .B1(KEYINPUT26), .B2(new_n351), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n351), .A2(KEYINPUT26), .ZN(new_n366));
  INV_X1    g165(.A(G169gat), .ZN(new_n367));
  INV_X1    g166(.A(G176gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n345), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n356), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n344), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AOI211_X1 g173(.A(KEYINPUT68), .B(new_n372), .C1(new_n356), .C2(new_n370), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n354), .B(KEYINPUT25), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(KEYINPUT65), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT65), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n365), .A2(new_n379), .A3(new_n345), .A4(new_n369), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n377), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n372), .B1(new_n381), .B2(KEYINPUT29), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n343), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n373), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n371), .A2(new_n385), .A3(new_n372), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n341), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(KEYINPUT69), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(G8gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(new_n235), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OR4_X1    g191(.A1(KEYINPUT30), .A2(new_n383), .A3(new_n387), .A4(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n372), .B1(new_n356), .B2(new_n370), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(new_n344), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n356), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n373), .B1(new_n397), .B2(new_n385), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n342), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n387), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n391), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n392), .B1(new_n383), .B2(new_n387), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT30), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n319), .A2(new_n317), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n299), .A2(new_n304), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n405), .A2(new_n316), .ZN(new_n406));
  OAI211_X1 g205(.A(KEYINPUT5), .B(new_n404), .C1(new_n315), .C2(new_n406), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n317), .A2(KEYINPUT5), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n315), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n409), .A3(KEYINPUT78), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT78), .B1(new_n407), .B2(new_n409), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n328), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n333), .A2(new_n393), .A3(new_n403), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n308), .ZN(new_n415));
  OR3_X1    g214(.A1(new_n415), .A2(KEYINPUT74), .A3(KEYINPUT29), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT74), .B1(new_n415), .B2(KEYINPUT29), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n342), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n305), .B1(new_n341), .B2(KEYINPUT29), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n299), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n418), .A2(G228gat), .A3(G233gat), .A4(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT72), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(KEYINPUT72), .A3(new_n299), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n341), .B1(new_n415), .B2(KEYINPUT29), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT73), .ZN(new_n427));
  NAND2_X1  g226(.A1(G228gat), .A2(G233gat), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n426), .B2(new_n428), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n421), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT75), .B(G22gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n432), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n421), .B(new_n434), .C1(new_n429), .C2(new_n430), .ZN(new_n435));
  XOR2_X1   g234(.A(G78gat), .B(G106gat), .Z(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT31), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(new_n224), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT76), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n435), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n438), .A2(G22gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n431), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n435), .B2(new_n441), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT79), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n407), .A2(new_n409), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT78), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n329), .B1(new_n451), .B2(new_n410), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n449), .B2(new_n328), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n448), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n395), .A2(new_n398), .A3(new_n342), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n384), .A2(new_n341), .A3(new_n386), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT37), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT37), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n399), .A2(new_n459), .A3(new_n400), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT38), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n458), .A2(new_n460), .A3(new_n461), .A4(new_n392), .ZN(new_n462));
  INV_X1    g261(.A(new_n454), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n413), .A2(KEYINPUT79), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n328), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(new_n453), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n455), .A2(new_n462), .A3(new_n464), .A4(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT37), .B1(new_n383), .B2(new_n387), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n460), .A2(new_n469), .A3(new_n392), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n401), .B1(new_n470), .B2(new_n461), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n414), .B(new_n447), .C1(new_n468), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n397), .A2(new_n304), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n381), .A2(new_n311), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT34), .ZN(new_n476));
  INV_X1    g275(.A(G227gat), .ZN(new_n477));
  INV_X1    g276(.A(G233gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n473), .A2(new_n474), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT34), .B1(new_n482), .B2(new_n479), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT32), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n482), .A2(new_n479), .B1(new_n485), .B2(KEYINPUT33), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G43gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G71gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G99gat), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n489), .A2(KEYINPUT66), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(KEYINPUT66), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(KEYINPUT33), .A3(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(KEYINPUT32), .B(new_n493), .C1(new_n475), .C2(new_n480), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n484), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n494), .B1(new_n486), .B2(new_n489), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n483), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT36), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n466), .B1(new_n465), .B2(new_n463), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n393), .B2(new_n403), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n472), .B(new_n503), .C1(new_n505), .C2(new_n447), .ZN(new_n506));
  INV_X1    g305(.A(new_n446), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n495), .A2(new_n507), .A3(new_n498), .A4(new_n442), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n393), .A2(new_n403), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n463), .A2(new_n465), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n467), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT35), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n495), .A2(new_n498), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n455), .A2(new_n464), .A3(new_n467), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n514), .A2(new_n447), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n509), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n513), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n292), .B1(new_n506), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT9), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n521), .A2(G71gat), .A3(G78gat), .ZN(new_n522));
  AND2_X1   g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  INV_X1    g322(.A(G57gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(G64gat), .ZN(new_n525));
  INV_X1    g324(.A(G64gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(G57gat), .ZN(new_n527));
  OAI22_X1  g326(.A1(new_n522), .A2(new_n523), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT9), .B1(new_n525), .B2(new_n527), .ZN(new_n529));
  XNOR2_X1  g328(.A(G71gat), .B(G78gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT90), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(G57gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n524), .A2(G64gat), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n521), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n535), .A2(new_n536), .A3(new_n530), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n528), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT21), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n218), .B(new_n347), .C1(new_n544), .C2(new_n538), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n538), .A2(new_n544), .ZN(new_n546));
  OAI21_X1  g345(.A(G183gat), .B1(new_n260), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(KEYINPUT91), .ZN(new_n549));
  INV_X1    g348(.A(G231gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(new_n478), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(KEYINPUT91), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n551), .B1(new_n549), .B2(new_n552), .ZN(new_n555));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(new_n336), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n557), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n549), .A2(new_n552), .ZN(new_n560));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n559), .B1(new_n562), .B2(new_n553), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n543), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n557), .B1(new_n554), .B2(new_n555), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n553), .A3(new_n559), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n542), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT92), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT92), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(G99gat), .A3(G106gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n572), .A3(KEYINPUT8), .ZN(new_n573));
  OR2_X1    g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT7), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(G85gat), .A3(G92gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G99gat), .B(G106gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n573), .A2(new_n579), .A3(new_n581), .A4(new_n574), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n283), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n587));
  INV_X1    g386(.A(new_n585), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n261), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G190gat), .B(G218gat), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT93), .ZN(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(new_n592), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n594), .A2(new_n593), .A3(new_n599), .A4(new_n597), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G120gat), .B(G148gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(new_n368), .ZN(new_n605));
  INV_X1    g404(.A(G204gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n538), .A2(new_n585), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n529), .A2(new_n531), .A3(KEYINPUT90), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n536), .B1(new_n535), .B2(new_n530), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n612), .A2(new_n584), .A3(new_n583), .A4(new_n528), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT94), .B(KEYINPUT10), .Z(new_n614));
  NAND3_X1  g413(.A1(new_n609), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n539), .A2(new_n588), .A3(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n609), .A2(new_n613), .ZN(new_n620));
  INV_X1    g419(.A(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n608), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT96), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n615), .A2(new_n616), .A3(KEYINPUT95), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT95), .B1(new_n615), .B2(new_n616), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n618), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(new_n608), .A3(new_n622), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n568), .A2(new_n603), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n520), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n504), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g436(.A1(new_n635), .A2(new_n518), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n214), .A2(new_n217), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n641), .A2(KEYINPUT42), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(KEYINPUT42), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n642), .B(new_n643), .C1(new_n217), .C2(new_n638), .ZN(G1325gat));
  AOI21_X1  g443(.A(G15gat), .B1(new_n635), .B2(new_n514), .ZN(new_n645));
  INV_X1    g444(.A(new_n503), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n646), .A2(G15gat), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n645), .B1(new_n635), .B2(new_n647), .ZN(G1326gat));
  NAND2_X1  g447(.A1(new_n507), .A2(new_n442), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n635), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT43), .B(G22gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n653));
  INV_X1    g452(.A(new_n603), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT100), .B1(new_n505), .B2(new_n447), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n512), .A2(new_n656), .A3(new_n649), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n472), .A2(new_n655), .A3(new_n503), .A4(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n654), .B1(new_n658), .B2(new_n519), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n653), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n654), .B1(new_n506), .B2(new_n519), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n660), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n662), .A2(new_n653), .A3(new_n660), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n279), .A2(KEYINPUT98), .A3(new_n290), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n286), .A2(new_n287), .B1(new_n265), .B2(KEYINPUT88), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n272), .A2(new_n277), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n208), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n288), .A2(new_n265), .A3(new_n289), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n668), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n568), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n631), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n666), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G29gat), .B1(new_n677), .B2(new_n511), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n662), .A2(new_n291), .A3(new_n676), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n234), .A3(new_n504), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT45), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n678), .A2(new_n681), .A3(KEYINPUT101), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(G1328gat));
  OAI21_X1  g485(.A(G36gat), .B1(new_n677), .B2(new_n509), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n509), .B1(new_n688), .B2(KEYINPUT46), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n679), .A2(new_n235), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n688), .A2(KEYINPUT46), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT103), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n687), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(G1329gat));
  NAND4_X1  g496(.A1(new_n666), .A2(new_n646), .A3(new_n674), .A4(new_n676), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n223), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT47), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n223), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n679), .A2(new_n514), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n699), .B(new_n703), .C1(new_n700), .C2(KEYINPUT47), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1330gat));
  OAI21_X1  g506(.A(G50gat), .B1(new_n677), .B2(new_n447), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n679), .A2(new_n224), .A3(new_n649), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n708), .B2(new_n710), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(G1331gat));
  AOI211_X1 g512(.A(new_n603), .B(new_n568), .C1(new_n658), .C2(new_n519), .ZN(new_n714));
  INV_X1    g513(.A(new_n631), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n674), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n511), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(new_n524), .ZN(G1332gat));
  INV_X1    g518(.A(new_n717), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT49), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n518), .B1(new_n721), .B2(new_n526), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT105), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n526), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1333gat));
  NAND3_X1  g525(.A1(new_n720), .A2(G71gat), .A3(new_n646), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n717), .A2(new_n499), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(G71gat), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT106), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g530(.A1(new_n720), .A2(new_n649), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n568), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT107), .Z(new_n735));
  NAND4_X1  g534(.A1(new_n666), .A2(G85gat), .A3(new_n504), .A4(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(G85gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n658), .A2(new_n519), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n675), .A2(new_n674), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n603), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(KEYINPUT51), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n631), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n737), .B1(new_n745), .B2(new_n511), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n736), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1336gat));
  NOR2_X1   g548(.A1(new_n509), .A2(G92gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n659), .A2(new_n751), .A3(new_n739), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n659), .B2(new_n739), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT110), .B1(new_n754), .B2(new_n743), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT109), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n659), .A2(new_n751), .A3(new_n739), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n756), .A2(KEYINPUT110), .A3(new_n743), .A4(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n744), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n631), .B(new_n750), .C1(new_n755), .C2(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n518), .B(new_n735), .C1(new_n664), .C2(new_n665), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G92gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT52), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n631), .B(new_n750), .C1(new_n742), .C2(new_n744), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n763), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(KEYINPUT111), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n766), .B1(new_n761), .B2(new_n763), .ZN(new_n771));
  INV_X1    g570(.A(new_n768), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(G1337gat));
  XOR2_X1   g573(.A(KEYINPUT112), .B(G99gat), .Z(new_n775));
  NAND2_X1  g574(.A1(new_n666), .A2(new_n735), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n776), .B2(new_n503), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n745), .A2(new_n775), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n499), .B2(new_n778), .ZN(G1338gat));
  OAI21_X1  g578(.A(G106gat), .B1(new_n776), .B2(new_n447), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n447), .A2(G106gat), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n780), .B(new_n781), .C1(new_n745), .C2(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n631), .B(new_n782), .C1(new_n755), .C2(new_n760), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n786), .B2(new_n781), .ZN(G1339gat));
  NOR2_X1   g586(.A1(new_n617), .A2(new_n618), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n629), .A2(KEYINPUT54), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n607), .B1(new_n619), .B2(KEYINPUT54), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n790), .B2(new_n793), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n630), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n667), .B2(new_n673), .ZN(new_n797));
  INV_X1    g596(.A(new_n206), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n273), .A2(new_n262), .A3(new_n275), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT113), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n284), .A2(new_n259), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n631), .A2(new_n290), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n654), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n796), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n290), .A2(new_n802), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n603), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n568), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  INV_X1    g609(.A(new_n674), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n632), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n508), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n675), .B1(new_n804), .B2(new_n807), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n632), .A2(new_n811), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT114), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n813), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n509), .A2(new_n504), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n292), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n821), .A2(G113gat), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n811), .ZN(G1340gat));
  XNOR2_X1  g623(.A(KEYINPUT115), .B(G120gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(KEYINPUT115), .A2(G120gat), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n821), .A2(new_n715), .ZN(new_n827));
  MUX2_X1   g626(.A(new_n825), .B(new_n826), .S(new_n827), .Z(G1341gat));
  INV_X1    g627(.A(new_n821), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n675), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n603), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(G134gat), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT56), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(KEYINPUT116), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(G134gat), .ZN(new_n836));
  XNOR2_X1  g635(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n835), .B(new_n836), .C1(new_n833), .C2(new_n837), .ZN(G1343gat));
  NAND3_X1  g637(.A1(new_n813), .A2(new_n817), .A3(new_n649), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n503), .A2(new_n820), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(G141gat), .A3(new_n292), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(KEYINPUT58), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT95), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n617), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n626), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n788), .B1(new_n849), .B2(new_n618), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n792), .B1(new_n850), .B2(KEYINPUT54), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n791), .B1(new_n851), .B2(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n790), .A2(new_n793), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT55), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n291), .A3(new_n630), .ZN(new_n857));
  INV_X1    g656(.A(new_n803), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n603), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n807), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n846), .B(new_n568), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n812), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n852), .A2(new_n855), .B1(new_n279), .B2(new_n290), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n803), .B1(new_n863), .B2(new_n630), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n807), .B1(new_n864), .B2(new_n603), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n846), .B1(new_n865), .B2(new_n568), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n649), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n841), .B1(new_n867), .B2(KEYINPUT57), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n813), .A2(new_n817), .A3(new_n869), .A4(new_n649), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(new_n291), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G141gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n845), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n867), .A2(KEYINPUT57), .ZN(new_n875));
  AND4_X1   g674(.A1(new_n874), .A2(new_n875), .A3(new_n842), .A4(new_n870), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n868), .B2(new_n870), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n674), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n844), .B1(new_n878), .B2(G141gat), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n873), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g682(.A(KEYINPUT120), .B(new_n873), .C1(new_n879), .C2(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1344gat));
  NAND2_X1  g684(.A1(new_n634), .A2(new_n292), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n865), .A2(new_n568), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n447), .A2(KEYINPUT57), .ZN(new_n889));
  AOI22_X1  g688(.A1(KEYINPUT57), .A2(new_n839), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n890), .A2(KEYINPUT59), .A3(new_n631), .A4(new_n842), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n877), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n715), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n891), .B1(new_n893), .B2(KEYINPUT59), .ZN(new_n894));
  INV_X1    g693(.A(new_n843), .ZN(new_n895));
  AOI21_X1  g694(.A(G148gat), .B1(new_n895), .B2(new_n631), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n894), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n896), .ZN(G1345gat));
  AOI21_X1  g696(.A(G155gat), .B1(new_n895), .B2(new_n675), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n892), .A2(new_n568), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(G155gat), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n892), .B2(new_n654), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n654), .A2(G162gat), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n902), .B1(new_n843), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n895), .A2(KEYINPUT121), .A3(new_n903), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n509), .A2(new_n504), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n813), .A2(new_n817), .A3(new_n814), .A4(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n367), .A3(new_n674), .ZN(new_n911));
  OAI21_X1  g710(.A(G169gat), .B1(new_n909), .B2(new_n292), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1348gat));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n631), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n915), .A3(G176gat), .ZN(new_n916));
  XOR2_X1   g715(.A(KEYINPUT122), .B(G176gat), .Z(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n914), .B2(new_n917), .ZN(G1349gat));
  OAI21_X1  g717(.A(new_n347), .B1(new_n909), .B2(new_n568), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n910), .A2(new_n675), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n363), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT60), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(KEYINPUT123), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(KEYINPUT123), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n926), .B1(new_n921), .B2(new_n922), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n921), .A2(new_n926), .A3(new_n922), .ZN(new_n928));
  OAI22_X1  g727(.A1(new_n924), .A2(new_n925), .B1(new_n927), .B2(new_n928), .ZN(G1350gat));
  XNOR2_X1  g728(.A(KEYINPUT61), .B(G190gat), .ZN(new_n930));
  NAND2_X1  g729(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n909), .A2(new_n654), .ZN(new_n932));
  MUX2_X1   g731(.A(new_n930), .B(new_n931), .S(new_n932), .Z(G1351gat));
  NAND2_X1  g732(.A1(new_n503), .A2(new_n908), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n890), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n292), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n839), .A2(new_n934), .ZN(new_n938));
  INV_X1    g737(.A(G197gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n674), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT125), .ZN(G1352gat));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n936), .B2(new_n715), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n890), .A2(KEYINPUT126), .A3(new_n631), .A4(new_n935), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(G204gat), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n938), .A2(new_n606), .A3(new_n631), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(G1353gat));
  OAI21_X1  g749(.A(G211gat), .B1(new_n936), .B2(new_n568), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(KEYINPUT127), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n336), .A3(new_n675), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n951), .A2(new_n957), .A3(new_n952), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n936), .B2(new_n654), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n938), .A2(new_n337), .A3(new_n603), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1355gat));
endmodule


