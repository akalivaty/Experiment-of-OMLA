

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U550 ( .A1(n685), .A2(n913), .ZN(n684) );
  NOR2_X2 U551 ( .A1(n528), .A2(n527), .ZN(G160) );
  OR2_X1 U552 ( .A1(n792), .A2(n782), .ZN(n516) );
  NOR2_X1 U553 ( .A1(n912), .A2(n682), .ZN(n683) );
  XNOR2_X1 U554 ( .A(n684), .B(KEYINPUT102), .ZN(n692) );
  NOR2_X1 U555 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U556 ( .A1(n783), .A2(n516), .ZN(n784) );
  NOR2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  NOR2_X1 U558 ( .A1(G651), .A2(n635), .ZN(n646) );
  XOR2_X2 U559 ( .A(KEYINPUT17), .B(n517), .Z(n874) );
  NAND2_X1 U560 ( .A1(n874), .A2(G137), .ZN(n518) );
  XNOR2_X1 U561 ( .A(n518), .B(KEYINPUT68), .ZN(n522) );
  XOR2_X1 U562 ( .A(KEYINPUT23), .B(KEYINPUT66), .Z(n520) );
  INV_X1 U563 ( .A(G2105), .ZN(n523) );
  AND2_X1 U564 ( .A1(n523), .A2(G2104), .ZN(n873) );
  NAND2_X1 U565 ( .A1(G101), .A2(n873), .ZN(n519) );
  XNOR2_X1 U566 ( .A(n520), .B(n519), .ZN(n521) );
  NAND2_X1 U567 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n523), .ZN(n870) );
  NAND2_X1 U569 ( .A1(n870), .A2(G125), .ZN(n526) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n869) );
  NAND2_X1 U571 ( .A1(G113), .A2(n869), .ZN(n524) );
  XOR2_X1 U572 ( .A(KEYINPUT67), .B(n524), .Z(n525) );
  NAND2_X1 U573 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U574 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U575 ( .A1(G85), .A2(n638), .ZN(n530) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n635) );
  INV_X1 U577 ( .A(G651), .ZN(n531) );
  NOR2_X1 U578 ( .A1(n635), .A2(n531), .ZN(n642) );
  NAND2_X1 U579 ( .A1(G72), .A2(n642), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n536) );
  NOR2_X1 U581 ( .A1(G543), .A2(n531), .ZN(n532) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n532), .Z(n639) );
  NAND2_X1 U583 ( .A1(G60), .A2(n639), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G47), .A2(n646), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n535) );
  OR2_X1 U586 ( .A1(n536), .A2(n535), .ZN(G290) );
  NAND2_X1 U587 ( .A1(G64), .A2(n639), .ZN(n538) );
  NAND2_X1 U588 ( .A1(G52), .A2(n646), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n538), .A2(n537), .ZN(n543) );
  NAND2_X1 U590 ( .A1(G90), .A2(n638), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G77), .A2(n642), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U593 ( .A(KEYINPUT9), .B(n541), .Z(n542) );
  NOR2_X1 U594 ( .A1(n543), .A2(n542), .ZN(G171) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U596 ( .A1(G65), .A2(n639), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G53), .A2(n646), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U599 ( .A1(G91), .A2(n638), .ZN(n547) );
  NAND2_X1 U600 ( .A1(G78), .A2(n642), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n917) );
  INV_X1 U603 ( .A(n917), .ZN(G299) );
  INV_X1 U604 ( .A(G132), .ZN(G219) );
  INV_X1 U605 ( .A(G82), .ZN(G220) );
  INV_X1 U606 ( .A(G57), .ZN(G237) );
  NAND2_X1 U607 ( .A1(G63), .A2(n639), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G51), .A2(n646), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U610 ( .A(KEYINPUT6), .B(n552), .ZN(n560) );
  NAND2_X1 U611 ( .A1(G89), .A2(n638), .ZN(n553) );
  XNOR2_X1 U612 ( .A(n553), .B(KEYINPUT4), .ZN(n554) );
  XNOR2_X1 U613 ( .A(n554), .B(KEYINPUT74), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G76), .A2(n642), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U616 ( .A(KEYINPUT5), .B(n557), .ZN(n558) );
  XNOR2_X1 U617 ( .A(KEYINPUT75), .B(n558), .ZN(n559) );
  NOR2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U619 ( .A(KEYINPUT7), .B(n561), .Z(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(G102), .A2(n873), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G138), .A2(n874), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U624 ( .A1(G114), .A2(n869), .ZN(n565) );
  NAND2_X1 U625 ( .A1(G126), .A2(n870), .ZN(n564) );
  NAND2_X1 U626 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U627 ( .A1(n567), .A2(n566), .ZN(G164) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U629 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U630 ( .A(G223), .ZN(n817) );
  NAND2_X1 U631 ( .A1(n817), .A2(G567), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U633 ( .A1(n638), .A2(G81), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U635 ( .A1(G68), .A2(n642), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U637 ( .A(KEYINPUT13), .B(n573), .Z(n577) );
  NAND2_X1 U638 ( .A1(G56), .A2(n639), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(KEYINPUT14), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT69), .ZN(n576) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n646), .A2(G43), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n912) );
  INV_X1 U644 ( .A(G860), .ZN(n595) );
  OR2_X1 U645 ( .A1(n912), .A2(n595), .ZN(G153) );
  XOR2_X1 U646 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U648 ( .A1(n646), .A2(G54), .ZN(n580) );
  XOR2_X1 U649 ( .A(KEYINPUT71), .B(n580), .Z(n582) );
  NAND2_X1 U650 ( .A1(n642), .A2(G79), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U652 ( .A(KEYINPUT72), .B(n583), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G92), .A2(n638), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G66), .A2(n639), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U657 ( .A(KEYINPUT73), .B(KEYINPUT15), .ZN(n588) );
  XNOR2_X1 U658 ( .A(n589), .B(n588), .ZN(n913) );
  OR2_X1 U659 ( .A1(n913), .A2(G868), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(G284) );
  INV_X1 U661 ( .A(G868), .ZN(n660) );
  XNOR2_X1 U662 ( .A(KEYINPUT76), .B(n660), .ZN(n592) );
  NOR2_X1 U663 ( .A1(G286), .A2(n592), .ZN(n594) );
  NOR2_X1 U664 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U665 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U666 ( .A1(n595), .A2(G559), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n596), .A2(n913), .ZN(n597) );
  XNOR2_X1 U668 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n912), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G868), .A2(n913), .ZN(n598) );
  NOR2_X1 U671 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U672 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U673 ( .A1(G99), .A2(n873), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G111), .A2(n869), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n603), .B(KEYINPUT77), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G135), .A2(n874), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n870), .A2(G123), .ZN(n606) );
  XOR2_X1 U680 ( .A(KEYINPUT18), .B(n606), .Z(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n991) );
  XOR2_X1 U682 ( .A(G2096), .B(n991), .Z(n609) );
  NOR2_X1 U683 ( .A1(G2100), .A2(n609), .ZN(n610) );
  XOR2_X1 U684 ( .A(KEYINPUT78), .B(n610), .Z(G156) );
  NAND2_X1 U685 ( .A1(G67), .A2(n639), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G55), .A2(n646), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U688 ( .A(n613), .B(KEYINPUT81), .ZN(n615) );
  NAND2_X1 U689 ( .A1(G93), .A2(n638), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n642), .A2(G80), .ZN(n616) );
  XOR2_X1 U692 ( .A(KEYINPUT80), .B(n616), .Z(n617) );
  OR2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n659) );
  NAND2_X1 U694 ( .A1(n913), .A2(G559), .ZN(n657) );
  XOR2_X1 U695 ( .A(KEYINPUT79), .B(n912), .Z(n619) );
  XNOR2_X1 U696 ( .A(n657), .B(n619), .ZN(n620) );
  NOR2_X1 U697 ( .A1(G860), .A2(n620), .ZN(n621) );
  XOR2_X1 U698 ( .A(n659), .B(n621), .Z(G145) );
  NAND2_X1 U699 ( .A1(n646), .A2(G50), .ZN(n622) );
  XNOR2_X1 U700 ( .A(n622), .B(KEYINPUT82), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G62), .A2(n639), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(KEYINPUT83), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G88), .A2(n638), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n642), .A2(G75), .ZN(n628) );
  XOR2_X1 U707 ( .A(KEYINPUT84), .B(n628), .Z(n629) );
  NOR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U709 ( .A(KEYINPUT85), .B(n631), .Z(G166) );
  NAND2_X1 U710 ( .A1(G49), .A2(n646), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U713 ( .A1(n639), .A2(n634), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n635), .A2(G87), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U716 ( .A1(G86), .A2(n638), .ZN(n641) );
  NAND2_X1 U717 ( .A1(G61), .A2(n639), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n642), .A2(G73), .ZN(n643) );
  XOR2_X1 U720 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U722 ( .A1(n646), .A2(G48), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(G305) );
  XNOR2_X1 U724 ( .A(G166), .B(n912), .ZN(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n650) );
  XNOR2_X1 U726 ( .A(G288), .B(KEYINPUT87), .ZN(n649) );
  XNOR2_X1 U727 ( .A(n650), .B(n649), .ZN(n653) );
  XOR2_X1 U728 ( .A(n659), .B(G290), .Z(n651) );
  XNOR2_X1 U729 ( .A(n651), .B(G299), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n654), .B(G305), .ZN(n655) );
  XNOR2_X1 U732 ( .A(n656), .B(n655), .ZN(n889) );
  XNOR2_X1 U733 ( .A(n657), .B(n889), .ZN(n658) );
  NAND2_X1 U734 ( .A1(n658), .A2(G868), .ZN(n662) );
  NAND2_X1 U735 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U741 ( .A1(n666), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U743 ( .A1(G69), .A2(G120), .ZN(n667) );
  NOR2_X1 U744 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U745 ( .A1(G108), .A2(n668), .ZN(n821) );
  NAND2_X1 U746 ( .A1(n821), .A2(G567), .ZN(n674) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U749 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U750 ( .A1(G96), .A2(n671), .ZN(n822) );
  NAND2_X1 U751 ( .A1(G2106), .A2(n822), .ZN(n672) );
  XNOR2_X1 U752 ( .A(KEYINPUT88), .B(n672), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n674), .A2(n673), .ZN(n824) );
  NAND2_X1 U754 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U755 ( .A1(n824), .A2(n675), .ZN(n820) );
  NAND2_X1 U756 ( .A1(n820), .A2(G36), .ZN(G176) );
  XNOR2_X1 U757 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  NAND2_X1 U758 ( .A1(G160), .A2(G40), .ZN(n747) );
  INV_X1 U759 ( .A(n747), .ZN(n679) );
  AND2_X1 U760 ( .A1(n679), .A2(G1996), .ZN(n677) );
  NOR2_X1 U761 ( .A1(G1384), .A2(G164), .ZN(n676) );
  XNOR2_X1 U762 ( .A(n676), .B(KEYINPUT64), .ZN(n746) );
  NAND2_X1 U763 ( .A1(n677), .A2(n746), .ZN(n678) );
  XNOR2_X1 U764 ( .A(n678), .B(KEYINPUT26), .ZN(n681) );
  NAND2_X1 U765 ( .A1(n679), .A2(n746), .ZN(n724) );
  NAND2_X1 U766 ( .A1(n724), .A2(G1341), .ZN(n680) );
  NAND2_X1 U767 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U768 ( .A(KEYINPUT65), .B(n683), .Z(n685) );
  NAND2_X1 U769 ( .A1(n685), .A2(n913), .ZN(n690) );
  INV_X1 U770 ( .A(G2067), .ZN(n966) );
  NOR2_X1 U771 ( .A1(n724), .A2(n966), .ZN(n686) );
  XNOR2_X1 U772 ( .A(n686), .B(KEYINPUT101), .ZN(n688) );
  NAND2_X1 U773 ( .A1(n724), .A2(G1348), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U776 ( .A1(n692), .A2(n691), .ZN(n697) );
  INV_X1 U777 ( .A(n724), .ZN(n706) );
  NAND2_X1 U778 ( .A1(n706), .A2(G2072), .ZN(n693) );
  XNOR2_X1 U779 ( .A(n693), .B(KEYINPUT27), .ZN(n695) );
  INV_X1 U780 ( .A(G1956), .ZN(n844) );
  NOR2_X1 U781 ( .A1(n844), .A2(n706), .ZN(n694) );
  NOR2_X1 U782 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U783 ( .A1(n698), .A2(n917), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n697), .A2(n696), .ZN(n702) );
  NOR2_X1 U785 ( .A1(n698), .A2(n917), .ZN(n700) );
  XOR2_X1 U786 ( .A(KEYINPUT28), .B(KEYINPUT100), .Z(n699) );
  XNOR2_X1 U787 ( .A(n700), .B(n699), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n702), .A2(n701), .ZN(n704) );
  XNOR2_X1 U789 ( .A(KEYINPUT29), .B(KEYINPUT103), .ZN(n703) );
  XNOR2_X1 U790 ( .A(n704), .B(n703), .ZN(n710) );
  OR2_X1 U791 ( .A1(n706), .A2(G1961), .ZN(n708) );
  XOR2_X1 U792 ( .A(G2078), .B(KEYINPUT99), .Z(n705) );
  XNOR2_X1 U793 ( .A(KEYINPUT25), .B(n705), .ZN(n968) );
  NAND2_X1 U794 ( .A1(n706), .A2(n968), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n714) );
  NAND2_X1 U796 ( .A1(n714), .A2(G171), .ZN(n709) );
  NAND2_X1 U797 ( .A1(n710), .A2(n709), .ZN(n730) );
  NOR2_X1 U798 ( .A1(G2084), .A2(n724), .ZN(n721) );
  NAND2_X1 U799 ( .A1(G8), .A2(n724), .ZN(n792) );
  NOR2_X1 U800 ( .A1(G1966), .A2(n792), .ZN(n718) );
  NOR2_X1 U801 ( .A1(n721), .A2(n718), .ZN(n711) );
  NAND2_X1 U802 ( .A1(G8), .A2(n711), .ZN(n712) );
  XNOR2_X1 U803 ( .A(KEYINPUT30), .B(n712), .ZN(n713) );
  NOR2_X1 U804 ( .A1(G168), .A2(n713), .ZN(n716) );
  NOR2_X1 U805 ( .A1(G171), .A2(n714), .ZN(n715) );
  NOR2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U807 ( .A(KEYINPUT31), .B(n717), .Z(n728) );
  AND2_X1 U808 ( .A1(n730), .A2(n728), .ZN(n719) );
  XNOR2_X1 U809 ( .A(n720), .B(KEYINPUT104), .ZN(n723) );
  NAND2_X1 U810 ( .A1(n721), .A2(G8), .ZN(n722) );
  NAND2_X1 U811 ( .A1(n723), .A2(n722), .ZN(n739) );
  XOR2_X1 U812 ( .A(KEYINPUT32), .B(KEYINPUT105), .Z(n737) );
  NOR2_X1 U813 ( .A1(G1971), .A2(n792), .ZN(n726) );
  NOR2_X1 U814 ( .A1(G2090), .A2(n724), .ZN(n725) );
  NOR2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U816 ( .A1(n727), .A2(G303), .ZN(n731) );
  AND2_X1 U817 ( .A1(n728), .A2(n731), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n734) );
  INV_X1 U819 ( .A(n731), .ZN(n732) );
  OR2_X1 U820 ( .A1(n732), .A2(G286), .ZN(n733) );
  AND2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U822 ( .A1(G8), .A2(n735), .ZN(n736) );
  XNOR2_X1 U823 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U824 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U825 ( .A(n740), .B(KEYINPUT106), .ZN(n787) );
  NOR2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n781) );
  NOR2_X1 U827 ( .A1(G1971), .A2(G303), .ZN(n741) );
  NOR2_X1 U828 ( .A1(n781), .A2(n741), .ZN(n925) );
  NAND2_X1 U829 ( .A1(n787), .A2(n925), .ZN(n744) );
  INV_X1 U830 ( .A(n792), .ZN(n742) );
  NAND2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n918) );
  AND2_X1 U832 ( .A1(n742), .A2(n918), .ZN(n743) );
  AND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U834 ( .A1(KEYINPUT33), .A2(n745), .ZN(n785) );
  XOR2_X1 U835 ( .A(G1981), .B(G305), .Z(n932) );
  NOR2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n812) );
  XNOR2_X1 U837 ( .A(G2067), .B(KEYINPUT37), .ZN(n748) );
  XNOR2_X1 U838 ( .A(n748), .B(KEYINPUT90), .ZN(n810) );
  NAND2_X1 U839 ( .A1(G104), .A2(n873), .ZN(n750) );
  NAND2_X1 U840 ( .A1(G140), .A2(n874), .ZN(n749) );
  NAND2_X1 U841 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U842 ( .A(KEYINPUT34), .B(n751), .ZN(n756) );
  NAND2_X1 U843 ( .A1(G116), .A2(n869), .ZN(n753) );
  NAND2_X1 U844 ( .A1(G128), .A2(n870), .ZN(n752) );
  NAND2_X1 U845 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U846 ( .A(KEYINPUT35), .B(n754), .Z(n755) );
  NOR2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U848 ( .A(KEYINPUT36), .B(n757), .ZN(n886) );
  NOR2_X1 U849 ( .A1(n810), .A2(n886), .ZN(n985) );
  NAND2_X1 U850 ( .A1(n812), .A2(n985), .ZN(n808) );
  NAND2_X1 U851 ( .A1(n869), .A2(G107), .ZN(n758) );
  XNOR2_X1 U852 ( .A(KEYINPUT92), .B(n758), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n870), .A2(G119), .ZN(n759) );
  XOR2_X1 U854 ( .A(KEYINPUT91), .B(n759), .Z(n760) );
  NAND2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U856 ( .A(KEYINPUT93), .B(n762), .ZN(n767) );
  NAND2_X1 U857 ( .A1(G95), .A2(n873), .ZN(n764) );
  NAND2_X1 U858 ( .A1(G131), .A2(n874), .ZN(n763) );
  NAND2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U860 ( .A(KEYINPUT94), .B(n765), .Z(n766) );
  NAND2_X1 U861 ( .A1(n767), .A2(n766), .ZN(n866) );
  AND2_X1 U862 ( .A1(n866), .A2(G1991), .ZN(n778) );
  XOR2_X1 U863 ( .A(KEYINPUT96), .B(KEYINPUT38), .Z(n769) );
  NAND2_X1 U864 ( .A1(G105), .A2(n873), .ZN(n768) );
  XNOR2_X1 U865 ( .A(n769), .B(n768), .ZN(n774) );
  NAND2_X1 U866 ( .A1(G117), .A2(n869), .ZN(n771) );
  NAND2_X1 U867 ( .A1(G129), .A2(n870), .ZN(n770) );
  NAND2_X1 U868 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U869 ( .A(KEYINPUT95), .B(n772), .Z(n773) );
  NOR2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U871 ( .A1(n874), .A2(G141), .ZN(n775) );
  NAND2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n883) );
  AND2_X1 U873 ( .A1(n883), .A2(G1996), .ZN(n777) );
  OR2_X1 U874 ( .A1(n778), .A2(n777), .ZN(n984) );
  AND2_X1 U875 ( .A1(n984), .A2(n812), .ZN(n805) );
  XNOR2_X1 U876 ( .A(KEYINPUT97), .B(n805), .ZN(n779) );
  NAND2_X1 U877 ( .A1(n808), .A2(n779), .ZN(n797) );
  INV_X1 U878 ( .A(n797), .ZN(n780) );
  AND2_X1 U879 ( .A1(n932), .A2(n780), .ZN(n783) );
  NAND2_X1 U880 ( .A1(n781), .A2(KEYINPUT33), .ZN(n782) );
  OR2_X1 U881 ( .A1(n785), .A2(n784), .ZN(n799) );
  NOR2_X1 U882 ( .A1(G2090), .A2(G303), .ZN(n786) );
  NAND2_X1 U883 ( .A1(G8), .A2(n786), .ZN(n788) );
  NAND2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n789) );
  AND2_X1 U885 ( .A1(n789), .A2(n792), .ZN(n795) );
  NOR2_X1 U886 ( .A1(G1981), .A2(G305), .ZN(n790) );
  XOR2_X1 U887 ( .A(n790), .B(KEYINPUT24), .Z(n791) );
  NOR2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U889 ( .A(n793), .B(KEYINPUT98), .ZN(n794) );
  NOR2_X1 U890 ( .A1(n795), .A2(n794), .ZN(n796) );
  OR2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n801) );
  XNOR2_X1 U893 ( .A(G1986), .B(G290), .ZN(n921) );
  NAND2_X1 U894 ( .A1(n921), .A2(n812), .ZN(n800) );
  NAND2_X1 U895 ( .A1(n801), .A2(n800), .ZN(n815) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n883), .ZN(n802) );
  XOR2_X1 U897 ( .A(KEYINPUT107), .B(n802), .Z(n987) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n866), .ZN(n995) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n803) );
  NOR2_X1 U900 ( .A1(n995), .A2(n803), .ZN(n804) );
  NOR2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U902 ( .A1(n987), .A2(n806), .ZN(n807) );
  XNOR2_X1 U903 ( .A(n807), .B(KEYINPUT39), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n810), .A2(n886), .ZN(n992) );
  NAND2_X1 U906 ( .A1(n811), .A2(n992), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U909 ( .A(n816), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n817), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U912 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(G188) );
  INV_X1 U916 ( .A(G120), .ZN(G236) );
  INV_X1 U917 ( .A(G96), .ZN(G221) );
  INV_X1 U918 ( .A(G69), .ZN(G235) );
  NOR2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n823), .B(KEYINPUT110), .ZN(G325) );
  INV_X1 U921 ( .A(G325), .ZN(G261) );
  INV_X1 U922 ( .A(n824), .ZN(G319) );
  XOR2_X1 U923 ( .A(KEYINPUT42), .B(KEYINPUT111), .Z(n826) );
  XNOR2_X1 U924 ( .A(G2678), .B(KEYINPUT112), .ZN(n825) );
  XNOR2_X1 U925 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U926 ( .A(KEYINPUT43), .B(G2090), .Z(n828) );
  XNOR2_X1 U927 ( .A(G2067), .B(G2072), .ZN(n827) );
  XNOR2_X1 U928 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U929 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U930 ( .A(G2096), .B(G2100), .ZN(n831) );
  XNOR2_X1 U931 ( .A(n832), .B(n831), .ZN(n834) );
  XOR2_X1 U932 ( .A(G2084), .B(G2078), .Z(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(G227) );
  XOR2_X1 U934 ( .A(G1961), .B(G1966), .Z(n836) );
  XNOR2_X1 U935 ( .A(G1981), .B(G1976), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U937 ( .A(G1971), .B(G1986), .Z(n838) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U940 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U941 ( .A(KEYINPUT113), .B(G2474), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U943 ( .A(KEYINPUT41), .B(n843), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(G229) );
  NAND2_X1 U945 ( .A1(G124), .A2(n870), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n846), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U947 ( .A1(n869), .A2(G112), .ZN(n847) );
  NAND2_X1 U948 ( .A1(n848), .A2(n847), .ZN(n852) );
  NAND2_X1 U949 ( .A1(G100), .A2(n873), .ZN(n850) );
  NAND2_X1 U950 ( .A1(G136), .A2(n874), .ZN(n849) );
  NAND2_X1 U951 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U952 ( .A1(n852), .A2(n851), .ZN(G162) );
  XOR2_X1 U953 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n854) );
  XNOR2_X1 U954 ( .A(G164), .B(KEYINPUT117), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(n855), .B(KEYINPUT48), .Z(n857) );
  XNOR2_X1 U957 ( .A(G160), .B(KEYINPUT46), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(n858), .B(n991), .Z(n868) );
  NAND2_X1 U960 ( .A1(G103), .A2(n873), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G139), .A2(n874), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G115), .A2(n869), .ZN(n862) );
  NAND2_X1 U964 ( .A1(G127), .A2(n870), .ZN(n861) );
  NAND2_X1 U965 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U966 ( .A(KEYINPUT47), .B(n863), .Z(n864) );
  NOR2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n998) );
  XOR2_X1 U968 ( .A(n866), .B(n998), .Z(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n882) );
  NAND2_X1 U970 ( .A1(G118), .A2(n869), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G130), .A2(n870), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n880) );
  NAND2_X1 U973 ( .A1(G106), .A2(n873), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G142), .A2(n874), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U976 ( .A(KEYINPUT45), .B(n877), .Z(n878) );
  XNOR2_X1 U977 ( .A(KEYINPUT114), .B(n878), .ZN(n879) );
  NOR2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U979 ( .A(n882), .B(n881), .Z(n885) );
  XOR2_X1 U980 ( .A(n883), .B(G162), .Z(n884) );
  XNOR2_X1 U981 ( .A(n885), .B(n884), .ZN(n887) );
  XNOR2_X1 U982 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U983 ( .A1(G37), .A2(n888), .ZN(G395) );
  XOR2_X1 U984 ( .A(KEYINPUT118), .B(n889), .Z(n891) );
  XNOR2_X1 U985 ( .A(G171), .B(G286), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U987 ( .A(n913), .B(n892), .ZN(n893) );
  NOR2_X1 U988 ( .A1(G37), .A2(n893), .ZN(G397) );
  XNOR2_X1 U989 ( .A(G2451), .B(G2427), .ZN(n903) );
  XOR2_X1 U990 ( .A(G2430), .B(G2443), .Z(n895) );
  XNOR2_X1 U991 ( .A(G2435), .B(G2438), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U993 ( .A(G2454), .B(KEYINPUT109), .Z(n897) );
  XNOR2_X1 U994 ( .A(G1348), .B(G1341), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U996 ( .A(n899), .B(n898), .Z(n901) );
  XNOR2_X1 U997 ( .A(G2446), .B(KEYINPUT108), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(n904), .A2(G14), .ZN(n911) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n905) );
  XOR2_X1 U1003 ( .A(KEYINPUT119), .B(n905), .Z(n906) );
  XNOR2_X1 U1004 ( .A(n906), .B(KEYINPUT49), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  INV_X1 U1010 ( .A(n911), .ZN(G401) );
  XOR2_X1 U1011 ( .A(n912), .B(G1341), .Z(n930) );
  XNOR2_X1 U1012 ( .A(G171), .B(G1961), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(G1348), .B(n913), .ZN(n914) );
  NAND2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(KEYINPUT123), .B(n916), .ZN(n923) );
  XNOR2_X1 U1016 ( .A(G1956), .B(n917), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n927) );
  NAND2_X1 U1020 ( .A1(G1971), .A2(G303), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(KEYINPUT124), .B(n928), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1025 ( .A(KEYINPUT125), .B(n931), .Z(n936) );
  XNOR2_X1 U1026 ( .A(G1966), .B(G168), .ZN(n933) );
  NAND2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1028 ( .A(KEYINPUT57), .B(n934), .Z(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1030 ( .A(KEYINPUT126), .B(n937), .Z(n939) );
  XNOR2_X1 U1031 ( .A(G16), .B(KEYINPUT56), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n1014) );
  XNOR2_X1 U1033 ( .A(G1966), .B(G21), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(G5), .B(G1961), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n952) );
  XNOR2_X1 U1036 ( .A(KEYINPUT59), .B(G1348), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(n942), .B(G4), .ZN(n949) );
  XNOR2_X1 U1038 ( .A(G1956), .B(G20), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(G1981), .B(G6), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(G19), .B(G1341), .ZN(n943) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1042 ( .A(KEYINPUT127), .B(n945), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1045 ( .A(KEYINPUT60), .B(n950), .Z(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n959) );
  XNOR2_X1 U1047 ( .A(G1976), .B(G23), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G1971), .B(G22), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n956) );
  XOR2_X1 U1050 ( .A(G1986), .B(G24), .Z(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(KEYINPUT58), .B(n957), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(KEYINPUT61), .B(n960), .ZN(n962) );
  INV_X1 U1055 ( .A(G16), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n963), .A2(G11), .ZN(n1012) );
  XNOR2_X1 U1058 ( .A(G1996), .B(G32), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(G33), .B(G2072), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n974) );
  XNOR2_X1 U1061 ( .A(G26), .B(n966), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n967), .A2(G28), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(n968), .B(G27), .ZN(n970) );
  XOR2_X1 U1064 ( .A(G1991), .B(G25), .Z(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n975), .B(KEYINPUT53), .ZN(n978) );
  XOR2_X1 U1069 ( .A(G2084), .B(G34), .Z(n976) );
  XNOR2_X1 U1070 ( .A(KEYINPUT54), .B(n976), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(G35), .B(G2090), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(KEYINPUT122), .B(n981), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(G29), .A2(n982), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n983), .B(KEYINPUT55), .ZN(n1010) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n1006) );
  XOR2_X1 U1078 ( .A(G2090), .B(G162), .Z(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1080 ( .A(KEYINPUT51), .B(n988), .Z(n989) );
  XNOR2_X1 U1081 ( .A(KEYINPUT120), .B(n989), .ZN(n997) );
  XOR2_X1 U1082 ( .A(G2084), .B(G160), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1004) );
  XNOR2_X1 U1087 ( .A(G2072), .B(n998), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(G164), .B(G2078), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1090 ( .A(KEYINPUT50), .B(n1001), .Z(n1002) );
  XNOR2_X1 U1091 ( .A(KEYINPUT121), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(KEYINPUT52), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(G29), .A2(n1008), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(KEYINPUT62), .B(n1015), .Z(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

