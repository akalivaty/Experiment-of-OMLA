//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT88), .B(G224), .Z(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT7), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT64), .B1(new_n193), .B2(G143), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n193), .A2(KEYINPUT65), .A3(G143), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT65), .B1(new_n193), .B2(G143), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT66), .B1(new_n193), .B2(G143), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n196), .A3(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n207), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G125), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n204), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n200), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n207), .A2(new_n211), .A3(new_n217), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n214), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n192), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT89), .ZN(new_n224));
  INV_X1    g038(.A(new_n206), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n196), .A2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT65), .ZN(new_n227));
  AND4_X1   g041(.A1(new_n211), .A2(new_n225), .A3(new_n227), .A4(new_n217), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n194), .B2(new_n197), .ZN(new_n229));
  INV_X1    g043(.A(new_n219), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(G125), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n215), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT89), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n192), .ZN(new_n235));
  XNOR2_X1  g049(.A(G110), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT86), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G116), .B(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n240));
  INV_X1    g054(.A(G116), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n241), .A2(KEYINPUT5), .A3(G119), .ZN(new_n242));
  INV_X1    g056(.A(G113), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n240), .A2(new_n244), .B1(new_n246), .B2(new_n239), .ZN(new_n247));
  OR2_X1    g061(.A1(KEYINPUT82), .A2(G104), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT3), .A2(G107), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT82), .A2(G104), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT83), .B(G101), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT3), .A2(G107), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G104), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT3), .A2(G107), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n251), .A2(new_n252), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(G107), .B1(new_n248), .B2(new_n250), .ZN(new_n257));
  INV_X1    g071(.A(G107), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT84), .B1(new_n258), .B2(G104), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT84), .ZN(new_n260));
  INV_X1    g074(.A(G104), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G107), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(G101), .B1(new_n257), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n247), .A2(new_n256), .A3(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n255), .B1(new_n249), .B2(new_n261), .ZN(new_n267));
  OAI21_X1  g081(.A(G101), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n268), .A2(KEYINPUT4), .A3(new_n256), .ZN(new_n269));
  INV_X1    g083(.A(new_n239), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n245), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n246), .A2(new_n239), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n274), .B(G101), .C1(new_n266), .C2(new_n267), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n238), .B(new_n265), .C1(new_n269), .C2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n224), .A2(new_n235), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n238), .A2(KEYINPUT8), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n236), .B(KEYINPUT86), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT8), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n265), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n247), .B1(new_n256), .B2(new_n264), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n232), .A2(new_n215), .A3(KEYINPUT7), .A4(new_n191), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n188), .B1(new_n278), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G210), .B1(G237), .B2(G902), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT90), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n265), .B1(new_n269), .B2(new_n276), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n280), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT6), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(KEYINPUT87), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n277), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n191), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n233), .B(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n295), .B(new_n280), .C1(KEYINPUT87), .C2(new_n297), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n290), .A2(new_n294), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n293), .B(new_n292), .C1(new_n306), .C2(new_n289), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n187), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G110), .B(G140), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n190), .A2(G227), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  AND4_X1   g126(.A1(new_n211), .A2(new_n225), .A3(new_n227), .A4(new_n212), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n202), .B1(new_n207), .B2(new_n211), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n256), .B(new_n264), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n264), .A2(new_n256), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n213), .A3(new_n204), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT11), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n320));
  INV_X1    g134(.A(G134), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G137), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(G137), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT11), .ZN(new_n327));
  INV_X1    g141(.A(G137), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G134), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n325), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G131), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n326), .A2(KEYINPUT11), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n327), .B1(new_n332), .B2(new_n329), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n320), .A2(new_n322), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n325), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT70), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n331), .A2(KEYINPUT70), .A3(new_n336), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n318), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT12), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n331), .B2(new_n336), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n342), .A2(new_n343), .B1(new_n318), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n315), .A2(new_n346), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n331), .A2(KEYINPUT70), .A3(new_n336), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT70), .B1(new_n331), .B2(new_n336), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n204), .A2(new_n213), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n351), .A2(KEYINPUT10), .A3(new_n256), .A4(new_n264), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n268), .A2(new_n256), .A3(KEYINPUT4), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n228), .A2(new_n231), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n275), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n347), .A2(new_n350), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n312), .B1(new_n345), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n347), .A2(new_n352), .A3(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n341), .ZN(new_n360));
  INV_X1    g174(.A(new_n312), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G469), .B1(new_n363), .B2(G902), .ZN(new_n364));
  INV_X1    g178(.A(G469), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT85), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n356), .A2(new_n366), .A3(new_n361), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n366), .B1(new_n356), .B2(new_n361), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n368), .A2(new_n345), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n361), .B1(new_n360), .B2(new_n356), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n365), .B(new_n188), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n364), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT9), .B(G234), .ZN(new_n374));
  OAI21_X1  g188(.A(G221), .B1(new_n374), .B2(G902), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT16), .ZN(new_n377));
  INV_X1    g191(.A(G140), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G125), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT77), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(G125), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n214), .A2(G140), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT16), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT77), .A4(G125), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n381), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n193), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n381), .A2(new_n384), .A3(G146), .A4(new_n385), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(KEYINPUT78), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT78), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n390), .A3(new_n193), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G237), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n190), .A3(G214), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT91), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G143), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT91), .B(G143), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n397), .B1(new_n398), .B2(new_n394), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT17), .A3(G131), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT93), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT93), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n399), .A2(new_n402), .A3(KEYINPUT17), .A4(G131), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n399), .A2(G131), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT17), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n399), .A2(G131), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n392), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n382), .A2(new_n383), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(new_n193), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT18), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(new_n334), .ZN(new_n413));
  OAI221_X1 g227(.A(new_n411), .B1(new_n399), .B2(new_n413), .C1(new_n407), .C2(new_n412), .ZN(new_n414));
  XOR2_X1   g228(.A(KEYINPUT92), .B(G104), .Z(new_n415));
  XNOR2_X1  g229(.A(G113), .B(G122), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n409), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT94), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n409), .A2(new_n414), .A3(KEYINPUT94), .A4(new_n417), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n405), .A2(new_n407), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n410), .B(KEYINPUT19), .Z(new_n424));
  OAI211_X1 g238(.A(new_n388), .B(new_n423), .C1(new_n424), .C2(G146), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n414), .ZN(new_n426));
  INV_X1    g240(.A(new_n417), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n430));
  NOR2_X1   g244(.A1(G475), .A2(G902), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n420), .A2(new_n421), .B1(new_n426), .B2(new_n427), .ZN(new_n433));
  INV_X1    g247(.A(new_n431), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT20), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT97), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n417), .B1(new_n409), .B2(new_n414), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n420), .B2(new_n421), .ZN(new_n439));
  OAI21_X1  g253(.A(G475), .B1(new_n439), .B2(G902), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n241), .A2(KEYINPUT14), .A3(G122), .ZN(new_n441));
  XNOR2_X1  g255(.A(G116), .B(G122), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(G107), .B(new_n441), .C1(new_n443), .C2(KEYINPUT14), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n196), .A2(G128), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n196), .A2(G128), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n446), .A2(new_n447), .A3(G134), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n446), .A2(new_n447), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(new_n321), .ZN(new_n450));
  OAI221_X1 g264(.A(new_n444), .B1(G107), .B2(new_n443), .C1(new_n448), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n321), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n442), .B(new_n258), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n446), .A2(KEYINPUT13), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT13), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n445), .A2(new_n455), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n454), .A2(new_n456), .A3(new_n447), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n452), .B(new_n453), .C1(new_n457), .C2(new_n321), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n374), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT75), .B(G217), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n190), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n462), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n451), .A2(new_n458), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(G902), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G478), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n467), .A2(KEYINPUT15), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n468), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G234), .ZN(new_n472));
  OAI211_X1 g286(.A(G952), .B(new_n190), .C1(new_n472), .C2(new_n393), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT95), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(G902), .B(G953), .C1(new_n472), .C2(new_n393), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n476), .B(KEYINPUT96), .Z(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT21), .B(G898), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n436), .A2(new_n437), .A3(new_n440), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n436), .A2(new_n440), .A3(new_n481), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT97), .ZN(new_n484));
  AOI211_X1 g298(.A(new_n309), .B(new_n376), .C1(new_n482), .C2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT29), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT67), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n228), .B2(new_n231), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n220), .A2(KEYINPUT67), .A3(new_n221), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n337), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n325), .B1(new_n329), .B2(KEYINPUT69), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT69), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n322), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G131), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n351), .A2(new_n336), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n354), .B1(new_n348), .B2(new_n349), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(KEYINPUT30), .A3(new_n495), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n500), .A3(new_n273), .ZN(new_n501));
  NOR2_X1   g315(.A1(G237), .A2(G953), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G210), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT27), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT26), .B(G101), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n273), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n499), .A2(new_n495), .A3(new_n508), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n501), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT28), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n509), .A2(new_n511), .B1(new_n273), .B2(new_n496), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n499), .A2(KEYINPUT28), .A3(new_n495), .A4(new_n508), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n486), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n336), .A2(new_n494), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n213), .B2(new_n204), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(new_n341), .B2(new_n354), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT73), .A3(new_n508), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n509), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n519), .B(new_n521), .C1(new_n518), .C2(new_n508), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT28), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n509), .A2(new_n511), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n506), .A2(KEYINPUT29), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n188), .B(new_n515), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G472), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n509), .A2(new_n506), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n508), .B1(new_n496), .B2(new_n497), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n529), .B1(new_n500), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n496), .A2(new_n273), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n524), .A2(new_n513), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n531), .A2(new_n532), .B1(new_n534), .B2(new_n507), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n507), .B1(new_n518), .B2(new_n508), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n501), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT71), .B1(new_n537), .B2(KEYINPUT31), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT71), .ZN(new_n539));
  AOI211_X1 g353(.A(new_n539), .B(new_n532), .C1(new_n501), .C2(new_n536), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n535), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT32), .ZN(new_n542));
  NOR2_X1   g356(.A1(G472), .A2(G902), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT72), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n541), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n542), .B1(new_n541), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n528), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT74), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT74), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n528), .B(new_n550), .C1(new_n546), .C2(new_n547), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT23), .ZN(new_n552));
  INV_X1    g366(.A(G119), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(G128), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n554), .B(new_n555), .C1(G119), .C2(new_n201), .ZN(new_n556));
  XNOR2_X1  g370(.A(G119), .B(G128), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT24), .B(G110), .Z(new_n558));
  AOI22_X1  g372(.A1(new_n556), .A2(G110), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n389), .A2(new_n391), .A3(new_n559), .ZN(new_n560));
  OAI22_X1  g374(.A1(new_n556), .A2(G110), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n410), .A2(new_n193), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n388), .A3(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n560), .A2(KEYINPUT80), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT79), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT22), .B(G137), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT80), .B1(new_n560), .B2(new_n563), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n568), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT25), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n572), .B2(KEYINPUT81), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n572), .A2(KEYINPUT81), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n461), .B1(new_n472), .B2(G902), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n577), .B(KEYINPUT76), .Z(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n574), .B2(new_n575), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n569), .A2(new_n571), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n188), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n485), .A2(new_n549), .A3(new_n551), .A4(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n585), .B(new_n252), .Z(G3));
  OAI21_X1  g400(.A(new_n539), .B1(new_n531), .B2(new_n532), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n537), .A2(KEYINPUT71), .A3(KEYINPUT31), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n589), .B2(new_n535), .ZN(new_n590));
  INV_X1    g404(.A(G472), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n534), .A2(new_n507), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n501), .A2(new_n536), .A3(new_n532), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n587), .B2(new_n588), .ZN(new_n595));
  OAI22_X1  g409(.A1(new_n590), .A2(new_n591), .B1(new_n544), .B2(new_n595), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n596), .A2(new_n376), .A3(new_n583), .ZN(new_n597));
  INV_X1    g411(.A(new_n187), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n292), .A2(KEYINPUT98), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n306), .B2(new_n289), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n286), .A2(new_n287), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n601), .A2(new_n277), .A3(new_n235), .A4(new_n224), .ZN(new_n602));
  INV_X1    g416(.A(new_n599), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n303), .A2(new_n602), .A3(new_n188), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n292), .A2(KEYINPUT98), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n598), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n480), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n430), .B1(new_n429), .B2(new_n431), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n433), .A2(KEYINPUT20), .A3(new_n434), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n440), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n463), .A2(new_n465), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n467), .A2(G902), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n617));
  OAI211_X1 g431(.A(KEYINPUT33), .B(new_n463), .C1(new_n465), .C2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n465), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(KEYINPUT100), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n615), .B(new_n616), .C1(new_n618), .C2(new_n620), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n621), .A2(KEYINPUT101), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(KEYINPUT101), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n466), .A2(G478), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n612), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n609), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n597), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  OAI211_X1 g444(.A(KEYINPUT102), .B(KEYINPUT20), .C1(new_n433), .C2(new_n434), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n440), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n432), .A2(new_n435), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n471), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n609), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n597), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  INV_X1    g453(.A(new_n375), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n364), .B2(new_n372), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n560), .A2(new_n563), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT103), .ZN(new_n643));
  INV_X1    g457(.A(new_n568), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(KEYINPUT36), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n643), .B(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n582), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n576), .A2(new_n579), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n596), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n309), .B1(new_n484), .B2(new_n482), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n475), .B1(new_n478), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n635), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n607), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n549), .A2(new_n658), .A3(new_n551), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  XOR2_X1   g476(.A(new_n657), .B(KEYINPUT39), .Z(new_n663));
  NAND2_X1  g477(.A1(new_n641), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n188), .B1(new_n522), .B2(new_n506), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n507), .B1(new_n501), .B2(new_n509), .ZN(new_n668));
  OAI21_X1  g482(.A(G472), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(new_n546), .B2(new_n547), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT38), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(new_n305), .B2(new_n308), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n304), .A2(new_n307), .A3(KEYINPUT38), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n672), .A2(new_n187), .A3(new_n648), .A4(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n612), .ZN(new_n675));
  INV_X1    g489(.A(new_n471), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n666), .A2(new_n670), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  NOR2_X1   g493(.A1(new_n626), .A2(new_n657), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n549), .A2(new_n551), .A3(new_n660), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  INV_X1    g496(.A(new_n551), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT32), .B1(new_n595), .B2(new_n544), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n541), .A2(new_n542), .A3(new_n545), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n550), .B1(new_n686), .B2(new_n528), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n369), .A2(new_n345), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n371), .B1(new_n690), .B2(new_n367), .ZN(new_n691));
  OAI21_X1  g505(.A(G469), .B1(new_n691), .B2(G902), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n372), .A3(new_n375), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n583), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n688), .A2(new_n689), .A3(new_n627), .A4(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n549), .A2(new_n551), .A3(new_n627), .A4(new_n694), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT104), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n549), .A2(new_n636), .A3(new_n551), .A4(new_n694), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  NAND2_X1  g516(.A1(new_n484), .A2(new_n482), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n659), .A2(new_n693), .A3(new_n648), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n549), .A2(new_n703), .A3(new_n551), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  NAND3_X1  g520(.A1(new_n607), .A2(new_n612), .A3(new_n471), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT105), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n676), .B1(new_n436), .B2(new_n440), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n710), .A3(new_n607), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n591), .B1(new_n541), .B2(new_n188), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n525), .A2(new_n507), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n537), .B(new_n532), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n544), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n713), .A2(new_n716), .A3(new_n583), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n693), .A2(new_n480), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n712), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  NOR3_X1   g534(.A1(new_n716), .A2(new_n713), .A3(new_n648), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n659), .A2(new_n693), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n680), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  XNOR2_X1  g538(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n304), .A2(new_n307), .A3(new_n187), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n376), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n549), .A2(new_n551), .A3(new_n584), .A4(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n680), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n583), .B1(new_n686), .B2(new_n528), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(KEYINPUT42), .A3(new_n680), .A4(new_n727), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  INV_X1    g548(.A(new_n658), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n728), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n321), .ZN(G36));
  NAND2_X1  g551(.A1(new_n358), .A2(new_n362), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n365), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n358), .A2(new_n741), .A3(KEYINPUT45), .A4(new_n362), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n358), .A2(KEYINPUT45), .A3(new_n362), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT107), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n740), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(G469), .A2(G902), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n745), .A2(KEYINPUT46), .A3(new_n746), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n372), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n726), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n375), .A3(new_n663), .A4(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n754));
  INV_X1    g568(.A(new_n625), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n754), .B1(new_n755), .B2(new_n612), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n612), .A2(KEYINPUT108), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n436), .A2(new_n758), .A3(new_n440), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n625), .A2(KEYINPUT43), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n756), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n596), .B2(new_n649), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n544), .B1(new_n589), .B2(new_n535), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n763), .B(new_n649), .C1(new_n713), .C2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n762), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n753), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n762), .B(KEYINPUT44), .C1(new_n764), .C2(new_n767), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  INV_X1    g588(.A(new_n750), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT46), .B1(new_n745), .B2(new_n746), .ZN(new_n776));
  INV_X1    g590(.A(new_n372), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n774), .B1(new_n778), .B2(new_n640), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n777), .B1(new_n747), .B2(new_n748), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n640), .B1(new_n780), .B2(new_n750), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n680), .A2(new_n583), .A3(new_n752), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n549), .B2(new_n551), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n701), .A2(new_n705), .A3(new_n719), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n698), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n788), .B1(new_n698), .B2(new_n790), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n721), .A2(new_n727), .A3(new_n680), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n549), .A2(new_n551), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n471), .A2(new_n657), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n752), .A2(new_n634), .A3(new_n632), .A4(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(new_n650), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n793), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n736), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n608), .B(new_n187), .C1(new_n305), .C2(new_n308), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n675), .A2(new_n471), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n800), .B1(new_n801), .B2(new_n626), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n597), .A2(new_n802), .B1(new_n651), .B2(new_n652), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n585), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n733), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n791), .A2(new_n792), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  INV_X1    g621(.A(new_n657), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n641), .A2(new_n648), .A3(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n709), .A2(new_n710), .A3(new_n607), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n710), .B1(new_n709), .B2(new_n607), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n670), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n641), .A2(new_n648), .A3(new_n808), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n686), .B2(new_n669), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT111), .B1(new_n816), .B2(new_n712), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n661), .A2(new_n681), .A3(new_n723), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT112), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n661), .A2(new_n681), .A3(new_n723), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n812), .A2(new_n813), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n816), .A2(new_n712), .A3(KEYINPUT111), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n807), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT112), .B1(new_n818), .B2(new_n819), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n822), .A2(new_n821), .A3(new_n825), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n829), .A3(KEYINPUT52), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n806), .A2(KEYINPUT53), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n807), .B1(new_n822), .B2(new_n825), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n828), .A2(new_n829), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(new_n807), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT53), .B1(new_n806), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n831), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g651(.A(KEYINPUT113), .B(KEYINPUT53), .C1(new_n806), .C2(new_n834), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT54), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n696), .B(new_n689), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n805), .A2(new_n841), .A3(new_n842), .A4(new_n789), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n834), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT110), .B1(new_n842), .B2(new_n789), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n698), .A2(new_n790), .A3(new_n788), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n585), .A2(new_n803), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n847), .A2(new_n736), .A3(new_n798), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n845), .A2(new_n733), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n828), .A2(new_n829), .A3(KEYINPUT52), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(new_n828), .B2(new_n829), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n840), .B(new_n844), .C1(new_n852), .C2(KEYINPUT53), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n791), .A2(new_n792), .ZN(new_n856));
  INV_X1    g670(.A(new_n805), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n827), .A3(new_n857), .A4(new_n830), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n858), .A2(new_n841), .B1(new_n834), .B2(new_n843), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(KEYINPUT114), .A3(new_n840), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n190), .A2(G952), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT120), .ZN(new_n863));
  INV_X1    g677(.A(new_n722), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n713), .A2(new_n716), .A3(new_n583), .A4(new_n474), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n762), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n692), .A2(new_n372), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n375), .A3(new_n752), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n868), .A2(KEYINPUT117), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n474), .B1(new_n868), .B2(KEYINPUT117), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n670), .A2(new_n583), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI221_X1 g687(.A(new_n863), .B1(new_n864), .B2(new_n866), .C1(new_n873), .C2(new_n626), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n871), .A2(new_n731), .A3(new_n762), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT48), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI211_X1 g693(.A(new_n187), .B(new_n693), .C1(new_n673), .C2(new_n672), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n762), .A2(new_n865), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT116), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT50), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n867), .A2(new_n640), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n779), .A2(new_n782), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n866), .A2(new_n726), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n675), .A2(new_n755), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n869), .A2(new_n872), .A3(new_n870), .A4(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n871), .A2(KEYINPUT118), .A3(new_n721), .A4(new_n762), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n869), .A2(new_n870), .A3(new_n762), .A4(new_n721), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n892), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n884), .B(new_n889), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n879), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n884), .A2(new_n897), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n888), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n783), .A2(KEYINPUT115), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n783), .A2(KEYINPUT115), .B1(new_n640), .B2(new_n867), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT51), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n861), .B1(new_n902), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n897), .A2(new_n898), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(new_n884), .A3(new_n900), .A4(new_n889), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n885), .B1(new_n903), .B2(new_n908), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT121), .A4(new_n879), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n839), .A2(new_n855), .A3(new_n860), .A4(new_n916), .ZN(new_n917));
  OR2_X1    g731(.A1(G952), .A2(G953), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n867), .B(KEYINPUT49), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n672), .A2(new_n673), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n640), .A2(new_n598), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n921), .A2(new_n584), .A3(new_n625), .A4(new_n922), .ZN(new_n923));
  OR4_X1    g737(.A1(new_n670), .A2(new_n920), .A3(new_n760), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n924), .ZN(G75));
  NOR2_X1   g739(.A1(new_n190), .A2(G952), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n858), .A2(new_n841), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n844), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n929), .A2(G210), .A3(G902), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n299), .A2(new_n302), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n301), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n934), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n927), .B1(new_n930), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n929), .A2(G210), .A3(G902), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT122), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n859), .A2(new_n188), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n943), .A3(G210), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n941), .A2(new_n944), .A3(new_n936), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n939), .B1(new_n945), .B2(new_n933), .ZN(G51));
  INV_X1    g760(.A(new_n942), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(new_n745), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n746), .B(KEYINPUT57), .Z(new_n949));
  INV_X1    g763(.A(new_n853), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n840), .B1(new_n928), .B2(new_n844), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n691), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n926), .B1(new_n948), .B2(new_n954), .ZN(G54));
  NAND2_X1  g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n947), .A2(new_n433), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n956), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n429), .B1(new_n942), .B2(new_n958), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n957), .A2(new_n959), .A3(new_n926), .ZN(G60));
  OAI21_X1  g774(.A(new_n615), .B1(new_n618), .B2(new_n620), .ZN(new_n961));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT59), .Z(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n950), .B2(new_n951), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n927), .ZN(new_n966));
  INV_X1    g780(.A(new_n963), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n855), .A2(new_n860), .ZN(new_n968));
  INV_X1    g782(.A(new_n832), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n827), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n841), .B1(new_n970), .B2(new_n849), .ZN(new_n971));
  AOI22_X1  g785(.A1(new_n971), .A2(KEYINPUT113), .B1(new_n852), .B2(KEYINPUT53), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n835), .A2(new_n836), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n840), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n967), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n966), .B1(new_n975), .B2(new_n961), .ZN(G63));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT60), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n929), .A2(new_n646), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n581), .B1(new_n859), .B2(new_n978), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n980), .A2(new_n981), .A3(new_n927), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n980), .A2(new_n981), .A3(KEYINPUT61), .A4(new_n927), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(G66));
  INV_X1    g800(.A(new_n479), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n190), .B1(new_n987), .B2(new_n189), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n856), .A2(new_n804), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(new_n190), .ZN(new_n990));
  INV_X1    g804(.A(G898), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n931), .B1(new_n991), .B2(G953), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n990), .B(new_n992), .ZN(G69));
  NAND2_X1  g807(.A1(new_n498), .A2(new_n500), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(new_n424), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT62), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n822), .A2(new_n997), .A3(new_n678), .ZN(new_n998));
  AOI22_X1  g812(.A1(new_n770), .A2(new_n771), .B1(new_n783), .B2(new_n785), .ZN(new_n999));
  INV_X1    g813(.A(new_n678), .ZN(new_n1000));
  OAI21_X1  g814(.A(KEYINPUT62), .B1(new_n819), .B2(new_n1000), .ZN(new_n1001));
  AOI211_X1 g815(.A(new_n726), .B(new_n664), .C1(new_n626), .C2(new_n801), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n688), .A2(new_n1002), .A3(new_n584), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(KEYINPUT124), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n772), .A2(new_n1003), .A3(new_n786), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT124), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1006), .A2(new_n1007), .A3(new_n1001), .A4(new_n998), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n996), .B1(new_n1009), .B2(new_n190), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n781), .A2(new_n712), .A3(new_n663), .A4(new_n731), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1014), .B1(new_n728), .B2(new_n735), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1015), .A2(new_n819), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n999), .A2(new_n1016), .A3(new_n733), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n190), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n190), .A2(G900), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(KEYINPUT125), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT125), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n1022), .B(new_n1019), .C1(new_n1017), .C2(new_n190), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n996), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1011), .A2(new_n1013), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT126), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1010), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g841(.A(KEYINPUT126), .B(new_n996), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1028));
  AOI211_X1 g842(.A(KEYINPUT127), .B(new_n1013), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT127), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1031), .A2(new_n1028), .A3(new_n1011), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1030), .B1(new_n1032), .B2(new_n1012), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1025), .B1(new_n1029), .B2(new_n1033), .ZN(G72));
  NOR2_X1   g848(.A1(new_n1009), .A2(new_n989), .ZN(new_n1035));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n668), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1037), .B1(new_n989), .B2(new_n1017), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n926), .B1(new_n1040), .B2(new_n510), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n972), .A2(new_n973), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n510), .A2(new_n668), .A3(new_n1038), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(G57));
endmodule


