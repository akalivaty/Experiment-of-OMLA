

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U552 ( .A(n517), .B(KEYINPUT64), .ZN(n866) );
  NOR2_X1 U553 ( .A1(n713), .A2(n731), .ZN(n714) );
  INV_X1 U554 ( .A(KEYINPUT31), .ZN(n719) );
  NAND2_X1 U555 ( .A1(n737), .A2(n736), .ZN(n744) );
  NAND2_X1 U556 ( .A1(n676), .A2(n761), .ZN(n712) );
  BUF_X1 U557 ( .A(n712), .Z(n723) );
  NOR2_X1 U558 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X2 U559 ( .A1(G2105), .A2(n518), .ZN(n861) );
  NOR2_X1 U560 ( .A1(n632), .A2(G651), .ZN(n630) );
  NOR2_X1 U561 ( .A1(n530), .A2(n529), .ZN(n675) );
  BUF_X1 U562 ( .A(n675), .Z(G160) );
  INV_X1 U563 ( .A(G2104), .ZN(n518) );
  AND2_X1 U564 ( .A1(G2105), .A2(n518), .ZN(n517) );
  NAND2_X1 U565 ( .A1(G125), .A2(n866), .ZN(n522) );
  NAND2_X1 U566 ( .A1(G101), .A2(n861), .ZN(n519) );
  XNOR2_X1 U567 ( .A(n519), .B(KEYINPUT65), .ZN(n520) );
  XNOR2_X1 U568 ( .A(n520), .B(KEYINPUT23), .ZN(n521) );
  NAND2_X1 U569 ( .A1(n522), .A2(n521), .ZN(n524) );
  INV_X1 U570 ( .A(KEYINPUT66), .ZN(n523) );
  XNOR2_X1 U571 ( .A(n524), .B(n523), .ZN(n526) );
  AND2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n864) );
  NAND2_X1 U573 ( .A1(n864), .A2(G113), .ZN(n525) );
  NAND2_X1 U574 ( .A1(n526), .A2(n525), .ZN(n530) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XOR2_X1 U576 ( .A(KEYINPUT17), .B(n527), .Z(n860) );
  NAND2_X1 U577 ( .A1(G137), .A2(n860), .ZN(n528) );
  XNOR2_X1 U578 ( .A(KEYINPUT67), .B(n528), .ZN(n529) );
  NOR2_X1 U579 ( .A1(G543), .A2(G651), .ZN(n621) );
  NAND2_X1 U580 ( .A1(n621), .A2(G89), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n531), .B(KEYINPUT4), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n632) );
  INV_X1 U583 ( .A(G651), .ZN(n535) );
  NOR2_X1 U584 ( .A1(n632), .A2(n535), .ZN(n624) );
  NAND2_X1 U585 ( .A1(G76), .A2(n624), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U587 ( .A(n534), .B(KEYINPUT5), .ZN(n541) );
  NOR2_X1 U588 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n536), .Z(n636) );
  NAND2_X1 U590 ( .A1(G63), .A2(n636), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G51), .A2(n630), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT6), .B(n539), .Z(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U595 ( .A(n542), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U596 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U597 ( .A1(G85), .A2(n621), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G72), .A2(n624), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G60), .A2(n636), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G47), .A2(n630), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U603 ( .A1(n548), .A2(n547), .ZN(G290) );
  NAND2_X1 U604 ( .A1(G64), .A2(n636), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G52), .A2(n630), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n556) );
  NAND2_X1 U607 ( .A1(n621), .A2(G90), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n551), .B(KEYINPUT68), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G77), .A2(n624), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U612 ( .A1(n556), .A2(n555), .ZN(G171) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U614 ( .A1(n866), .A2(G123), .ZN(n557) );
  XNOR2_X1 U615 ( .A(n557), .B(KEYINPUT18), .ZN(n564) );
  NAND2_X1 U616 ( .A1(G135), .A2(n860), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G111), .A2(n864), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G99), .A2(n861), .ZN(n560) );
  XNOR2_X1 U620 ( .A(KEYINPUT75), .B(n560), .ZN(n561) );
  NOR2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U622 ( .A1(n564), .A2(n563), .ZN(n914) );
  XNOR2_X1 U623 ( .A(G2096), .B(n914), .ZN(n565) );
  OR2_X1 U624 ( .A1(G2100), .A2(n565), .ZN(G156) );
  INV_X1 U625 ( .A(G82), .ZN(G220) );
  INV_X1 U626 ( .A(G120), .ZN(G236) );
  INV_X1 U627 ( .A(G69), .ZN(G235) );
  INV_X1 U628 ( .A(G108), .ZN(G238) );
  NAND2_X1 U629 ( .A1(G88), .A2(n621), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G75), .A2(n624), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT79), .B(n568), .ZN(n572) );
  NAND2_X1 U633 ( .A1(G62), .A2(n636), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G50), .A2(n630), .ZN(n569) );
  AND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(G303) );
  NAND2_X1 U637 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT72), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT10), .B(n574), .ZN(G223) );
  INV_X1 U640 ( .A(G223), .ZN(n815) );
  NAND2_X1 U641 ( .A1(n815), .A2(G567), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  NAND2_X1 U643 ( .A1(G56), .A2(n636), .ZN(n576) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(n576), .Z(n582) );
  NAND2_X1 U645 ( .A1(n621), .A2(G81), .ZN(n577) );
  XNOR2_X1 U646 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U647 ( .A1(G68), .A2(n624), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U649 ( .A(KEYINPUT13), .B(n580), .Z(n581) );
  NOR2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n630), .A2(G43), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n935) );
  XNOR2_X1 U653 ( .A(G860), .B(KEYINPUT73), .ZN(n605) );
  OR2_X1 U654 ( .A1(n935), .A2(n605), .ZN(G153) );
  INV_X1 U655 ( .A(G171), .ZN(G301) );
  NAND2_X1 U656 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n630), .A2(G54), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G66), .A2(n636), .ZN(n586) );
  NAND2_X1 U659 ( .A1(G92), .A2(n621), .ZN(n585) );
  NAND2_X1 U660 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n624), .A2(G79), .ZN(n587) );
  XOR2_X1 U662 ( .A(KEYINPUT74), .B(n587), .Z(n588) );
  NOR2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U665 ( .A(KEYINPUT15), .B(n592), .Z(n945) );
  INV_X1 U666 ( .A(G868), .ZN(n639) );
  NAND2_X1 U667 ( .A1(n945), .A2(n639), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U669 ( .A1(G78), .A2(n624), .ZN(n595) );
  XNOR2_X1 U670 ( .A(n595), .B(KEYINPUT70), .ZN(n602) );
  NAND2_X1 U671 ( .A1(G65), .A2(n636), .ZN(n597) );
  NAND2_X1 U672 ( .A1(G53), .A2(n630), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U674 ( .A1(G91), .A2(n621), .ZN(n598) );
  XNOR2_X1 U675 ( .A(KEYINPUT69), .B(n598), .ZN(n599) );
  NOR2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(G299) );
  NOR2_X1 U678 ( .A1(G286), .A2(n639), .ZN(n604) );
  NOR2_X1 U679 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U680 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U681 ( .A1(n605), .A2(G559), .ZN(n606) );
  INV_X1 U682 ( .A(n945), .ZN(n886) );
  NAND2_X1 U683 ( .A1(n606), .A2(n886), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G868), .A2(n935), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n886), .A2(G868), .ZN(n608) );
  NOR2_X1 U687 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U689 ( .A1(G559), .A2(n886), .ZN(n611) );
  XNOR2_X1 U690 ( .A(n611), .B(KEYINPUT76), .ZN(n650) );
  XNOR2_X1 U691 ( .A(n650), .B(n935), .ZN(n612) );
  NOR2_X1 U692 ( .A1(n612), .A2(G860), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G93), .A2(n621), .ZN(n614) );
  NAND2_X1 U694 ( .A1(G80), .A2(n624), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U696 ( .A(KEYINPUT77), .B(n615), .ZN(n619) );
  NAND2_X1 U697 ( .A1(G67), .A2(n636), .ZN(n617) );
  NAND2_X1 U698 ( .A1(G55), .A2(n630), .ZN(n616) );
  AND2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n641) );
  XOR2_X1 U701 ( .A(n620), .B(n641), .Z(G145) );
  NAND2_X1 U702 ( .A1(G61), .A2(n636), .ZN(n623) );
  NAND2_X1 U703 ( .A1(G86), .A2(n621), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n624), .A2(G73), .ZN(n625) );
  XOR2_X1 U706 ( .A(KEYINPUT2), .B(n625), .Z(n626) );
  NOR2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(G48), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G49), .A2(n630), .ZN(n631) );
  XNOR2_X1 U711 ( .A(n631), .B(KEYINPUT78), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G74), .A2(G651), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G87), .A2(n632), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(G288) );
  NAND2_X1 U717 ( .A1(n639), .A2(n641), .ZN(n640) );
  XNOR2_X1 U718 ( .A(n640), .B(KEYINPUT82), .ZN(n653) );
  XNOR2_X1 U719 ( .A(G303), .B(n641), .ZN(n648) );
  XNOR2_X1 U720 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n643) );
  XNOR2_X1 U721 ( .A(G305), .B(KEYINPUT19), .ZN(n642) );
  XNOR2_X1 U722 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U723 ( .A(n644), .B(G290), .ZN(n646) );
  XNOR2_X1 U724 ( .A(G299), .B(G288), .ZN(n645) );
  XNOR2_X1 U725 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U726 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U727 ( .A(n649), .B(n935), .ZN(n885) );
  XNOR2_X1 U728 ( .A(n885), .B(n650), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G868), .A2(n651), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(G295) );
  NAND2_X1 U731 ( .A1(G2078), .A2(G2084), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(KEYINPUT83), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n655), .B(KEYINPUT20), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n656), .A2(G2090), .ZN(n657) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n658), .A2(G2072), .ZN(n659) );
  XNOR2_X1 U737 ( .A(KEYINPUT84), .B(n659), .ZN(G158) );
  XNOR2_X1 U738 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U739 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NOR2_X1 U740 ( .A1(G235), .A2(G236), .ZN(n660) );
  XNOR2_X1 U741 ( .A(n660), .B(KEYINPUT85), .ZN(n661) );
  NOR2_X1 U742 ( .A1(G238), .A2(n661), .ZN(n662) );
  NAND2_X1 U743 ( .A1(G57), .A2(n662), .ZN(n821) );
  NAND2_X1 U744 ( .A1(n821), .A2(G567), .ZN(n667) );
  NOR2_X1 U745 ( .A1(G220), .A2(G219), .ZN(n663) );
  XOR2_X1 U746 ( .A(KEYINPUT22), .B(n663), .Z(n664) );
  NOR2_X1 U747 ( .A1(G218), .A2(n664), .ZN(n665) );
  NAND2_X1 U748 ( .A1(G96), .A2(n665), .ZN(n822) );
  NAND2_X1 U749 ( .A1(n822), .A2(G2106), .ZN(n666) );
  NAND2_X1 U750 ( .A1(n667), .A2(n666), .ZN(n823) );
  NAND2_X1 U751 ( .A1(G483), .A2(G661), .ZN(n668) );
  NOR2_X1 U752 ( .A1(n823), .A2(n668), .ZN(n818) );
  NAND2_X1 U753 ( .A1(n818), .A2(G36), .ZN(G176) );
  NAND2_X1 U754 ( .A1(G138), .A2(n860), .ZN(n670) );
  NAND2_X1 U755 ( .A1(G102), .A2(n861), .ZN(n669) );
  NAND2_X1 U756 ( .A1(n670), .A2(n669), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n864), .A2(G114), .ZN(n672) );
  NAND2_X1 U758 ( .A1(G126), .A2(n866), .ZN(n671) );
  NAND2_X1 U759 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U760 ( .A1(n674), .A2(n673), .ZN(G164) );
  NAND2_X1 U761 ( .A1(n675), .A2(G40), .ZN(n760) );
  INV_X1 U762 ( .A(n760), .ZN(n676) );
  NOR2_X1 U763 ( .A1(G164), .A2(G1384), .ZN(n761) );
  NAND2_X1 U764 ( .A1(G8), .A2(n723), .ZN(n750) );
  NOR2_X1 U765 ( .A1(G1981), .A2(G305), .ZN(n677) );
  XOR2_X1 U766 ( .A(n677), .B(KEYINPUT24), .Z(n678) );
  NOR2_X1 U767 ( .A1(n750), .A2(n678), .ZN(n758) );
  INV_X1 U768 ( .A(n712), .ZN(n693) );
  OR2_X1 U769 ( .A1(n693), .A2(G1961), .ZN(n680) );
  XNOR2_X1 U770 ( .A(KEYINPUT25), .B(G2078), .ZN(n973) );
  NAND2_X1 U771 ( .A1(n693), .A2(n973), .ZN(n679) );
  NAND2_X1 U772 ( .A1(n680), .A2(n679), .ZN(n716) );
  NAND2_X1 U773 ( .A1(n716), .A2(G171), .ZN(n707) );
  INV_X1 U774 ( .A(n712), .ZN(n688) );
  NAND2_X1 U775 ( .A1(n688), .A2(G2072), .ZN(n681) );
  XNOR2_X1 U776 ( .A(n681), .B(KEYINPUT27), .ZN(n683) );
  INV_X1 U777 ( .A(G1956), .ZN(n993) );
  NOR2_X1 U778 ( .A1(n993), .A2(n693), .ZN(n682) );
  NOR2_X2 U779 ( .A1(n683), .A2(n682), .ZN(n687) );
  INV_X1 U780 ( .A(G299), .ZN(n686) );
  NOR2_X1 U781 ( .A1(n687), .A2(n686), .ZN(n685) );
  XOR2_X1 U782 ( .A(KEYINPUT92), .B(KEYINPUT28), .Z(n684) );
  XNOR2_X1 U783 ( .A(n685), .B(n684), .ZN(n704) );
  NAND2_X1 U784 ( .A1(n687), .A2(n686), .ZN(n702) );
  AND2_X1 U785 ( .A1(n688), .A2(G1996), .ZN(n689) );
  XOR2_X1 U786 ( .A(n689), .B(KEYINPUT26), .Z(n692) );
  AND2_X1 U787 ( .A1(n723), .A2(G1341), .ZN(n690) );
  NOR2_X1 U788 ( .A1(n690), .A2(n935), .ZN(n691) );
  NAND2_X1 U789 ( .A1(n692), .A2(n691), .ZN(n697) );
  NAND2_X1 U790 ( .A1(G1348), .A2(n723), .ZN(n695) );
  NAND2_X1 U791 ( .A1(G2067), .A2(n693), .ZN(n694) );
  NAND2_X1 U792 ( .A1(n695), .A2(n694), .ZN(n698) );
  OR2_X1 U793 ( .A1(n945), .A2(n698), .ZN(n696) );
  NAND2_X1 U794 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n945), .A2(n698), .ZN(n699) );
  NAND2_X1 U796 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U799 ( .A(n705), .B(KEYINPUT29), .Z(n706) );
  NAND2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n722) );
  INV_X1 U801 ( .A(G8), .ZN(n708) );
  NOR2_X1 U802 ( .A1(n708), .A2(G1966), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n709), .A2(n712), .ZN(n711) );
  INV_X1 U804 ( .A(KEYINPUT91), .ZN(n710) );
  XNOR2_X1 U805 ( .A(n711), .B(n710), .ZN(n733) );
  NAND2_X1 U806 ( .A1(n733), .A2(G8), .ZN(n713) );
  NOR2_X1 U807 ( .A1(G2084), .A2(n712), .ZN(n731) );
  XOR2_X1 U808 ( .A(KEYINPUT30), .B(n714), .Z(n715) );
  NOR2_X1 U809 ( .A1(G168), .A2(n715), .ZN(n718) );
  NOR2_X1 U810 ( .A1(G171), .A2(n716), .ZN(n717) );
  NOR2_X1 U811 ( .A1(n718), .A2(n717), .ZN(n720) );
  XNOR2_X1 U812 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n732) );
  NAND2_X1 U814 ( .A1(n732), .A2(G286), .ZN(n728) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n750), .ZN(n725) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n723), .ZN(n724) );
  NOR2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U818 ( .A1(n726), .A2(G303), .ZN(n727) );
  NAND2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U820 ( .A1(G8), .A2(n729), .ZN(n730) );
  XNOR2_X1 U821 ( .A(n730), .B(KEYINPUT32), .ZN(n737) );
  NAND2_X1 U822 ( .A1(G8), .A2(n731), .ZN(n735) );
  AND2_X1 U823 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U824 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U825 ( .A1(G2090), .A2(G303), .ZN(n738) );
  NAND2_X1 U826 ( .A1(G8), .A2(n738), .ZN(n739) );
  NAND2_X1 U827 ( .A1(n744), .A2(n739), .ZN(n740) );
  XNOR2_X1 U828 ( .A(n740), .B(KEYINPUT94), .ZN(n741) );
  NAND2_X1 U829 ( .A1(n741), .A2(n750), .ZN(n756) );
  XOR2_X1 U830 ( .A(G1981), .B(G305), .Z(n956) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n942) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n742) );
  NOR2_X1 U833 ( .A1(n942), .A2(n742), .ZN(n743) );
  NAND2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n748) );
  INV_X1 U835 ( .A(n750), .ZN(n746) );
  NAND2_X1 U836 ( .A1(G288), .A2(G1976), .ZN(n745) );
  XOR2_X1 U837 ( .A(KEYINPUT93), .B(n745), .Z(n943) );
  AND2_X1 U838 ( .A1(n746), .A2(n943), .ZN(n747) );
  AND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U840 ( .A1(KEYINPUT33), .A2(n749), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n942), .A2(KEYINPUT33), .ZN(n751) );
  NOR2_X1 U842 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U844 ( .A1(n956), .A2(n754), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U846 ( .A(n759), .B(KEYINPUT95), .ZN(n794) );
  NOR2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n810) );
  NAND2_X1 U848 ( .A1(G141), .A2(n860), .ZN(n763) );
  NAND2_X1 U849 ( .A1(G129), .A2(n866), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n766) );
  NAND2_X1 U851 ( .A1(n861), .A2(G105), .ZN(n764) );
  XOR2_X1 U852 ( .A(KEYINPUT38), .B(n764), .Z(n765) );
  NOR2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n864), .A2(G117), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n875) );
  NAND2_X1 U856 ( .A1(G1996), .A2(n875), .ZN(n769) );
  XOR2_X1 U857 ( .A(KEYINPUT89), .B(n769), .Z(n777) );
  NAND2_X1 U858 ( .A1(G131), .A2(n860), .ZN(n771) );
  NAND2_X1 U859 ( .A1(G119), .A2(n866), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G95), .A2(n861), .ZN(n773) );
  NAND2_X1 U862 ( .A1(G107), .A2(n864), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  OR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n876) );
  NAND2_X1 U865 ( .A1(G1991), .A2(n876), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U867 ( .A(KEYINPUT90), .B(n778), .ZN(n911) );
  NAND2_X1 U868 ( .A1(n810), .A2(n911), .ZN(n800) );
  INV_X1 U869 ( .A(n800), .ZN(n792) );
  XOR2_X1 U870 ( .A(G2067), .B(KEYINPUT37), .Z(n807) );
  XNOR2_X1 U871 ( .A(KEYINPUT87), .B(KEYINPUT35), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n864), .A2(G116), .ZN(n780) );
  NAND2_X1 U873 ( .A1(G128), .A2(n866), .ZN(n779) );
  NAND2_X1 U874 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U875 ( .A(n782), .B(n781), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n861), .A2(G104), .ZN(n783) );
  XNOR2_X1 U877 ( .A(n783), .B(KEYINPUT86), .ZN(n785) );
  NAND2_X1 U878 ( .A1(G140), .A2(n860), .ZN(n784) );
  NAND2_X1 U879 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U880 ( .A(KEYINPUT34), .B(n786), .ZN(n787) );
  NOR2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U882 ( .A(KEYINPUT36), .B(n789), .Z(n882) );
  AND2_X1 U883 ( .A1(n807), .A2(n882), .ZN(n916) );
  NAND2_X1 U884 ( .A1(n916), .A2(n810), .ZN(n790) );
  XNOR2_X1 U885 ( .A(n790), .B(KEYINPUT88), .ZN(n805) );
  INV_X1 U886 ( .A(n805), .ZN(n791) );
  NOR2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n793) );
  AND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n796) );
  XNOR2_X1 U889 ( .A(G1986), .B(G290), .ZN(n937) );
  NAND2_X1 U890 ( .A1(n937), .A2(n810), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n813) );
  NOR2_X1 U892 ( .A1(G1996), .A2(n875), .ZN(n908) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n798) );
  NOR2_X1 U894 ( .A1(G1991), .A2(n876), .ZN(n797) );
  XNOR2_X1 U895 ( .A(KEYINPUT96), .B(n797), .ZN(n913) );
  NOR2_X1 U896 ( .A1(n798), .A2(n913), .ZN(n799) );
  XNOR2_X1 U897 ( .A(n799), .B(KEYINPUT97), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U899 ( .A(KEYINPUT98), .B(n802), .Z(n803) );
  NOR2_X1 U900 ( .A1(n908), .A2(n803), .ZN(n804) );
  XNOR2_X1 U901 ( .A(n804), .B(KEYINPUT39), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n807), .A2(n882), .ZN(n808) );
  XNOR2_X1 U904 ( .A(KEYINPUT99), .B(n808), .ZN(n927) );
  NAND2_X1 U905 ( .A1(n809), .A2(n927), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U908 ( .A(KEYINPUT40), .B(n814), .ZN(G329) );
  NAND2_X1 U909 ( .A1(G2106), .A2(n815), .ZN(G217) );
  AND2_X1 U910 ( .A1(G15), .A2(G2), .ZN(n816) );
  NAND2_X1 U911 ( .A1(G661), .A2(n816), .ZN(G259) );
  NAND2_X1 U912 ( .A1(G3), .A2(G1), .ZN(n817) );
  XNOR2_X1 U913 ( .A(KEYINPUT102), .B(n817), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U915 ( .A(KEYINPUT103), .B(n820), .Z(G188) );
  INV_X1 U917 ( .A(G96), .ZN(G221) );
  NOR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(G325) );
  INV_X1 U919 ( .A(G325), .ZN(G261) );
  INV_X1 U920 ( .A(n823), .ZN(G319) );
  XOR2_X1 U921 ( .A(G2096), .B(G2678), .Z(n825) );
  XNOR2_X1 U922 ( .A(G2072), .B(KEYINPUT43), .ZN(n824) );
  XNOR2_X1 U923 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U924 ( .A(n826), .B(KEYINPUT42), .Z(n828) );
  XNOR2_X1 U925 ( .A(G2067), .B(G2090), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U927 ( .A(KEYINPUT104), .B(G2100), .Z(n830) );
  XNOR2_X1 U928 ( .A(G2078), .B(G2084), .ZN(n829) );
  XNOR2_X1 U929 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(G227) );
  XOR2_X1 U931 ( .A(G1981), .B(G1966), .Z(n834) );
  XNOR2_X1 U932 ( .A(G1991), .B(G1986), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U934 ( .A(G1976), .B(G1971), .Z(n836) );
  XNOR2_X1 U935 ( .A(G1961), .B(G1956), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U937 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U938 ( .A(G2474), .B(KEYINPUT41), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U940 ( .A(KEYINPUT105), .B(n841), .ZN(n842) );
  XOR2_X1 U941 ( .A(n842), .B(G1996), .Z(G229) );
  NAND2_X1 U942 ( .A1(G100), .A2(n861), .ZN(n844) );
  NAND2_X1 U943 ( .A1(G112), .A2(n864), .ZN(n843) );
  NAND2_X1 U944 ( .A1(n844), .A2(n843), .ZN(n851) );
  XOR2_X1 U945 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n846) );
  NAND2_X1 U946 ( .A1(G124), .A2(n866), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U948 ( .A(KEYINPUT106), .B(n847), .ZN(n849) );
  NAND2_X1 U949 ( .A1(n860), .A2(G136), .ZN(n848) );
  NAND2_X1 U950 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U951 ( .A1(n851), .A2(n850), .ZN(G162) );
  NAND2_X1 U952 ( .A1(n864), .A2(G118), .ZN(n853) );
  NAND2_X1 U953 ( .A1(G130), .A2(n866), .ZN(n852) );
  NAND2_X1 U954 ( .A1(n853), .A2(n852), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G142), .A2(n860), .ZN(n855) );
  NAND2_X1 U956 ( .A1(G106), .A2(n861), .ZN(n854) );
  NAND2_X1 U957 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U958 ( .A(KEYINPUT45), .B(n856), .Z(n857) );
  NOR2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U960 ( .A(G160), .B(n859), .ZN(n874) );
  NAND2_X1 U961 ( .A1(G139), .A2(n860), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G103), .A2(n861), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n871) );
  NAND2_X1 U964 ( .A1(n864), .A2(G115), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n865), .B(KEYINPUT108), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G127), .A2(n866), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n921) );
  XOR2_X1 U970 ( .A(n921), .B(G162), .Z(n872) );
  XNOR2_X1 U971 ( .A(n914), .B(n872), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n879) );
  XNOR2_X1 U973 ( .A(G164), .B(n875), .ZN(n877) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U975 ( .A(n879), .B(n878), .Z(n881) );
  XNOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n881), .B(n880), .ZN(n883) );
  XNOR2_X1 U978 ( .A(n883), .B(n882), .ZN(n884) );
  NOR2_X1 U979 ( .A1(G37), .A2(n884), .ZN(G395) );
  XOR2_X1 U980 ( .A(n885), .B(G286), .Z(n888) );
  XNOR2_X1 U981 ( .A(G171), .B(n886), .ZN(n887) );
  XNOR2_X1 U982 ( .A(n888), .B(n887), .ZN(n889) );
  NOR2_X1 U983 ( .A1(G37), .A2(n889), .ZN(G397) );
  XNOR2_X1 U984 ( .A(G2443), .B(G2427), .ZN(n899) );
  XOR2_X1 U985 ( .A(G2430), .B(KEYINPUT101), .Z(n891) );
  XNOR2_X1 U986 ( .A(G2454), .B(G2435), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n895) );
  XOR2_X1 U988 ( .A(G2438), .B(KEYINPUT100), .Z(n893) );
  XNOR2_X1 U989 ( .A(G1341), .B(G1348), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U991 ( .A(n895), .B(n894), .Z(n897) );
  XNOR2_X1 U992 ( .A(G2451), .B(G2446), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  NAND2_X1 U995 ( .A1(n900), .A2(G14), .ZN(n906) );
  NAND2_X1 U996 ( .A1(G319), .A2(n906), .ZN(n903) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n901) );
  XNOR2_X1 U998 ( .A(KEYINPUT49), .B(n901), .ZN(n902) );
  NOR2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(G57), .ZN(G237) );
  INV_X1 U1004 ( .A(n906), .ZN(G401) );
  INV_X1 U1005 ( .A(KEYINPUT55), .ZN(n932) );
  XOR2_X1 U1006 ( .A(KEYINPUT110), .B(KEYINPUT52), .Z(n930) );
  XOR2_X1 U1007 ( .A(G2090), .B(G162), .Z(n907) );
  NOR2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n909), .B(KEYINPUT51), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n920) );
  XOR2_X1 U1011 ( .A(G160), .B(G2084), .Z(n912) );
  NOR2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1015 ( .A(KEYINPUT109), .B(n918), .Z(n919) );
  NAND2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n926) );
  XOR2_X1 U1017 ( .A(G2072), .B(n921), .Z(n923) );
  XOR2_X1 U1018 ( .A(G164), .B(G2078), .Z(n922) );
  NOR2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1020 ( .A(KEYINPUT50), .B(n924), .Z(n925) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n928) );
  NAND2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1023 ( .A(n930), .B(n929), .ZN(n931) );
  NAND2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1025 ( .A1(n933), .A2(G29), .ZN(n965) );
  XOR2_X1 U1026 ( .A(G1341), .B(KEYINPUT120), .Z(n934) );
  XNOR2_X1 U1027 ( .A(n935), .B(n934), .ZN(n939) );
  XNOR2_X1 U1028 ( .A(G1956), .B(G299), .ZN(n936) );
  NOR2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(G1971), .B(G303), .ZN(n940) );
  NOR2_X1 U1032 ( .A1(n941), .A2(n940), .ZN(n952) );
  XNOR2_X1 U1033 ( .A(KEYINPUT119), .B(n942), .ZN(n944) );
  NAND2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n950) );
  XNOR2_X1 U1035 ( .A(G301), .B(G1961), .ZN(n947) );
  XNOR2_X1 U1036 ( .A(n945), .B(G1348), .ZN(n946) );
  NOR2_X1 U1037 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1038 ( .A(KEYINPUT118), .B(n948), .Z(n949) );
  NOR2_X1 U1039 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1040 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1041 ( .A(n953), .B(KEYINPUT121), .ZN(n960) );
  XNOR2_X1 U1042 ( .A(G1966), .B(G168), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(n954), .B(KEYINPUT116), .ZN(n955) );
  NAND2_X1 U1044 ( .A1(n956), .A2(n955), .ZN(n958) );
  XOR2_X1 U1045 ( .A(KEYINPUT57), .B(KEYINPUT117), .Z(n957) );
  XNOR2_X1 U1046 ( .A(n958), .B(n957), .ZN(n959) );
  NAND2_X1 U1047 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1048 ( .A(G16), .B(KEYINPUT56), .Z(n961) );
  XNOR2_X1 U1049 ( .A(KEYINPUT115), .B(n961), .ZN(n962) );
  NAND2_X1 U1050 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1051 ( .A1(n965), .A2(n964), .ZN(n1022) );
  XNOR2_X1 U1052 ( .A(G2084), .B(G34), .ZN(n966) );
  XNOR2_X1 U1053 ( .A(n966), .B(KEYINPUT54), .ZN(n985) );
  XNOR2_X1 U1054 ( .A(G2090), .B(G35), .ZN(n982) );
  XNOR2_X1 U1055 ( .A(KEYINPUT111), .B(G2067), .ZN(n967) );
  XNOR2_X1 U1056 ( .A(n967), .B(G26), .ZN(n972) );
  XOR2_X1 U1057 ( .A(G1991), .B(G25), .Z(n968) );
  NAND2_X1 U1058 ( .A1(n968), .A2(G28), .ZN(n970) );
  XNOR2_X1 U1059 ( .A(G33), .B(G2072), .ZN(n969) );
  NOR2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1061 ( .A1(n972), .A2(n971), .ZN(n978) );
  XOR2_X1 U1062 ( .A(n973), .B(G27), .Z(n975) );
  XNOR2_X1 U1063 ( .A(G1996), .B(G32), .ZN(n974) );
  NOR2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1065 ( .A(n976), .B(KEYINPUT112), .Z(n977) );
  NOR2_X1 U1066 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1067 ( .A(KEYINPUT53), .B(n979), .Z(n980) );
  XNOR2_X1 U1068 ( .A(n980), .B(KEYINPUT113), .ZN(n981) );
  NOR2_X1 U1069 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1070 ( .A(KEYINPUT114), .B(n983), .Z(n984) );
  NOR2_X1 U1071 ( .A1(n985), .A2(n984), .ZN(n1016) );
  NAND2_X1 U1072 ( .A1(KEYINPUT55), .A2(n1016), .ZN(n986) );
  NAND2_X1 U1073 ( .A1(G11), .A2(n986), .ZN(n1015) );
  XNOR2_X1 U1074 ( .A(KEYINPUT123), .B(G1341), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(n987), .B(G19), .ZN(n992) );
  XOR2_X1 U1076 ( .A(G1348), .B(KEYINPUT59), .Z(n988) );
  XNOR2_X1 U1077 ( .A(G4), .B(n988), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(G6), .B(G1981), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n996) );
  XOR2_X1 U1081 ( .A(G20), .B(n993), .Z(n994) );
  XNOR2_X1 U1082 ( .A(KEYINPUT122), .B(n994), .ZN(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(KEYINPUT124), .B(n997), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(n998), .B(KEYINPUT60), .ZN(n1002) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G21), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(G1961), .B(G5), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1010) );
  XNOR2_X1 U1090 ( .A(G1986), .B(G24), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G23), .B(G1976), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G1971), .B(KEYINPUT125), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(G22), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(KEYINPUT58), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(KEYINPUT61), .B(n1011), .Z(n1012) );
  NOR2_X1 U1099 ( .A1(G16), .A2(n1012), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(n1013), .B(KEYINPUT126), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1020) );
  INV_X1 U1102 ( .A(n1016), .ZN(n1018) );
  NOR2_X1 U1103 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n1023) );
  XNOR2_X1 U1108 ( .A(n1024), .B(n1023), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
  INV_X1 U1110 ( .A(G303), .ZN(G166) );
endmodule

