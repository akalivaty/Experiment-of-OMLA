

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591;

  INV_X1 U322 ( .A(n351), .ZN(n505) );
  XNOR2_X2 U323 ( .A(n391), .B(n390), .ZN(n576) );
  NOR2_X1 U324 ( .A1(n517), .A2(n421), .ZN(n560) );
  XNOR2_X1 U325 ( .A(n418), .B(KEYINPUT54), .ZN(n419) );
  XNOR2_X2 U326 ( .A(KEYINPUT119), .B(n565), .ZN(n577) );
  XNOR2_X1 U327 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U328 ( .A(n438), .B(n437), .ZN(n563) );
  XOR2_X1 U329 ( .A(KEYINPUT69), .B(KEYINPUT7), .Z(n290) );
  XOR2_X1 U330 ( .A(n344), .B(n343), .Z(n291) );
  XNOR2_X1 U331 ( .A(KEYINPUT107), .B(KEYINPUT46), .ZN(n369) );
  XNOR2_X1 U332 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U333 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n463) );
  XNOR2_X1 U334 ( .A(n464), .B(n463), .ZN(n466) );
  INV_X1 U335 ( .A(G71GAT), .ZN(n428) );
  INV_X1 U336 ( .A(KEYINPUT118), .ZN(n418) );
  NOR2_X1 U337 ( .A1(n483), .A2(n586), .ZN(n475) );
  XNOR2_X1 U338 ( .A(n431), .B(n430), .ZN(n434) );
  XNOR2_X1 U339 ( .A(n345), .B(n291), .ZN(n346) );
  XNOR2_X1 U340 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U341 ( .A(n347), .B(n346), .ZN(n348) );
  INV_X1 U342 ( .A(KEYINPUT59), .ZN(n458) );
  XNOR2_X1 U343 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U344 ( .A(n479), .B(G36GAT), .ZN(n480) );
  XNOR2_X1 U345 ( .A(n461), .B(n460), .ZN(G1352GAT) );
  XNOR2_X1 U346 ( .A(n481), .B(n480), .ZN(G1329GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n457) );
  XOR2_X1 U348 ( .A(G57GAT), .B(KEYINPUT5), .Z(n293) );
  XNOR2_X1 U349 ( .A(G1GAT), .B(KEYINPUT89), .ZN(n292) );
  XNOR2_X1 U350 ( .A(n293), .B(n292), .ZN(n310) );
  XOR2_X1 U351 ( .A(G155GAT), .B(G148GAT), .Z(n295) );
  XNOR2_X1 U352 ( .A(G127GAT), .B(G162GAT), .ZN(n294) );
  XNOR2_X1 U353 ( .A(n295), .B(n294), .ZN(n297) );
  XOR2_X1 U354 ( .A(G29GAT), .B(G85GAT), .Z(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n306) );
  XNOR2_X1 U356 ( .A(KEYINPUT1), .B(KEYINPUT90), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n298), .B(KEYINPUT6), .ZN(n299) );
  XOR2_X1 U358 ( .A(n299), .B(KEYINPUT4), .Z(n304) );
  XOR2_X1 U359 ( .A(G120GAT), .B(KEYINPUT0), .Z(n301) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(G134GAT), .ZN(n300) );
  XNOR2_X1 U361 ( .A(n301), .B(n300), .ZN(n432) );
  XNOR2_X1 U362 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n302) );
  XNOR2_X1 U363 ( .A(n302), .B(KEYINPUT2), .ZN(n439) );
  XNOR2_X1 U364 ( .A(n432), .B(n439), .ZN(n303) );
  XNOR2_X1 U365 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n306), .B(n305), .ZN(n308) );
  NAND2_X1 U367 ( .A1(G225GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n517) );
  XOR2_X1 U370 ( .A(G78GAT), .B(G211GAT), .Z(n312) );
  XNOR2_X1 U371 ( .A(G1GAT), .B(G183GAT), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n325) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G127GAT), .Z(n427) );
  XOR2_X1 U374 ( .A(G22GAT), .B(G155GAT), .Z(n440) );
  XNOR2_X1 U375 ( .A(n427), .B(n440), .ZN(n314) );
  XNOR2_X1 U376 ( .A(G71GAT), .B(G57GAT), .ZN(n313) );
  XNOR2_X1 U377 ( .A(n313), .B(KEYINPUT13), .ZN(n342) );
  XNOR2_X1 U378 ( .A(n314), .B(n342), .ZN(n318) );
  XOR2_X1 U379 ( .A(G64GAT), .B(KEYINPUT14), .Z(n316) );
  NAND2_X1 U380 ( .A1(G231GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U381 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U382 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U383 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n320) );
  XNOR2_X1 U384 ( .A(KEYINPUT15), .B(KEYINPUT80), .ZN(n319) );
  XNOR2_X1 U385 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U386 ( .A(G8GAT), .B(n321), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U388 ( .A(n325), .B(n324), .Z(n538) );
  INV_X1 U389 ( .A(n538), .ZN(n586) );
  XOR2_X1 U390 ( .A(KEYINPUT71), .B(KEYINPUT75), .Z(n327) );
  XNOR2_X1 U391 ( .A(G120GAT), .B(KEYINPUT72), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n349) );
  INV_X1 U393 ( .A(G92GAT), .ZN(n328) );
  NAND2_X1 U394 ( .A1(G64GAT), .A2(n328), .ZN(n331) );
  INV_X1 U395 ( .A(G64GAT), .ZN(n329) );
  NAND2_X1 U396 ( .A1(n329), .A2(G92GAT), .ZN(n330) );
  NAND2_X1 U397 ( .A1(n331), .A2(n330), .ZN(n333) );
  XNOR2_X1 U398 ( .A(G176GAT), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U399 ( .A(n333), .B(n332), .ZN(n410) );
  INV_X1 U400 ( .A(n410), .ZN(n334) );
  XOR2_X1 U401 ( .A(G99GAT), .B(G85GAT), .Z(n379) );
  NAND2_X1 U402 ( .A1(n334), .A2(n379), .ZN(n337) );
  INV_X1 U403 ( .A(n379), .ZN(n335) );
  NAND2_X1 U404 ( .A1(n335), .A2(n410), .ZN(n336) );
  NAND2_X1 U405 ( .A1(n337), .A2(n336), .ZN(n339) );
  NAND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n347) );
  XOR2_X1 U408 ( .A(G78GAT), .B(G148GAT), .Z(n341) );
  XNOR2_X1 U409 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n340) );
  XNOR2_X1 U410 ( .A(n341), .B(n340), .ZN(n448) );
  XNOR2_X1 U411 ( .A(n448), .B(n342), .ZN(n345) );
  XOR2_X1 U412 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n344) );
  XNOR2_X1 U413 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n343) );
  XOR2_X1 U414 ( .A(n349), .B(n348), .Z(n580) );
  INV_X1 U415 ( .A(KEYINPUT41), .ZN(n350) );
  XNOR2_X1 U416 ( .A(n580), .B(n350), .ZN(n351) );
  XOR2_X1 U417 ( .A(KEYINPUT70), .B(KEYINPUT67), .Z(n353) );
  XNOR2_X1 U418 ( .A(G141GAT), .B(G1GAT), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n353), .B(n352), .ZN(n368) );
  XOR2_X1 U420 ( .A(G197GAT), .B(G22GAT), .Z(n355) );
  XNOR2_X1 U421 ( .A(G15GAT), .B(G113GAT), .ZN(n354) );
  XNOR2_X1 U422 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U423 ( .A(n356), .B(G36GAT), .Z(n358) );
  XOR2_X1 U424 ( .A(G169GAT), .B(G8GAT), .Z(n414) );
  XNOR2_X1 U425 ( .A(n414), .B(G50GAT), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U427 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n360) );
  NAND2_X1 U428 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U429 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U430 ( .A(n362), .B(n361), .Z(n366) );
  XNOR2_X1 U431 ( .A(G43GAT), .B(G29GAT), .ZN(n363) );
  XNOR2_X1 U432 ( .A(n290), .B(n363), .ZN(n364) );
  XOR2_X1 U433 ( .A(KEYINPUT8), .B(n364), .Z(n384) );
  XNOR2_X1 U434 ( .A(n384), .B(KEYINPUT29), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U436 ( .A(n368), .B(n367), .ZN(n531) );
  INV_X1 U437 ( .A(n531), .ZN(n566) );
  NAND2_X1 U438 ( .A1(n505), .A2(n566), .ZN(n370) );
  NOR2_X1 U439 ( .A1(n586), .A2(n371), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n372), .B(KEYINPUT108), .ZN(n392) );
  XOR2_X1 U441 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n374) );
  XNOR2_X1 U442 ( .A(G106GAT), .B(KEYINPUT77), .ZN(n373) );
  XNOR2_X1 U443 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U444 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n376) );
  XNOR2_X1 U445 ( .A(G92GAT), .B(KEYINPUT78), .ZN(n375) );
  XNOR2_X1 U446 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U447 ( .A(n378), .B(n377), .Z(n391) );
  XOR2_X1 U448 ( .A(G36GAT), .B(G190GAT), .Z(n406) );
  XNOR2_X1 U449 ( .A(KEYINPUT64), .B(n406), .ZN(n381) );
  XNOR2_X1 U450 ( .A(G218GAT), .B(n379), .ZN(n380) );
  XNOR2_X1 U451 ( .A(n381), .B(n380), .ZN(n383) );
  NAND2_X1 U452 ( .A1(G232GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n383), .B(n382), .ZN(n385) );
  XNOR2_X1 U454 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U455 ( .A(KEYINPUT9), .B(n386), .Z(n389) );
  XNOR2_X1 U456 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n387), .B(G162GAT), .ZN(n449) );
  XNOR2_X1 U458 ( .A(G134GAT), .B(n449), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n389), .B(n388), .ZN(n390) );
  INV_X1 U460 ( .A(n576), .ZN(n541) );
  NAND2_X1 U461 ( .A1(n392), .A2(n541), .ZN(n393) );
  XNOR2_X1 U462 ( .A(n393), .B(KEYINPUT47), .ZN(n399) );
  XOR2_X1 U463 ( .A(n576), .B(KEYINPUT98), .Z(n394) );
  XNOR2_X1 U464 ( .A(n394), .B(KEYINPUT36), .ZN(n589) );
  NOR2_X1 U465 ( .A1(n589), .A2(n538), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n395), .B(KEYINPUT45), .ZN(n396) );
  NAND2_X1 U467 ( .A1(n396), .A2(n580), .ZN(n397) );
  NOR2_X1 U468 ( .A1(n397), .A2(n566), .ZN(n398) );
  NOR2_X1 U469 ( .A1(n399), .A2(n398), .ZN(n400) );
  XNOR2_X1 U470 ( .A(n400), .B(KEYINPUT48), .ZN(n528) );
  XOR2_X1 U471 ( .A(G183GAT), .B(KEYINPUT19), .Z(n402) );
  XNOR2_X1 U472 ( .A(KEYINPUT86), .B(KEYINPUT17), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n402), .B(n401), .ZN(n404) );
  XOR2_X1 U474 ( .A(KEYINPUT18), .B(KEYINPUT85), .Z(n403) );
  XOR2_X1 U475 ( .A(n404), .B(n403), .Z(n438) );
  INV_X1 U476 ( .A(n438), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n406), .B(n405), .ZN(n408) );
  NAND2_X1 U478 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U479 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U480 ( .A(n410), .B(n409), .Z(n416) );
  XOR2_X1 U481 ( .A(KEYINPUT87), .B(G218GAT), .Z(n412) );
  XNOR2_X1 U482 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n411) );
  XNOR2_X1 U483 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U484 ( .A(G197GAT), .B(n413), .Z(n444) );
  XNOR2_X1 U485 ( .A(n414), .B(n444), .ZN(n415) );
  XNOR2_X1 U486 ( .A(n416), .B(n415), .ZN(n520) );
  XNOR2_X1 U487 ( .A(n520), .B(KEYINPUT117), .ZN(n417) );
  NOR2_X1 U488 ( .A1(n528), .A2(n417), .ZN(n420) );
  XNOR2_X1 U489 ( .A(KEYINPUT92), .B(KEYINPUT26), .ZN(n455) );
  XOR2_X1 U490 ( .A(KEYINPUT84), .B(G176GAT), .Z(n423) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(KEYINPUT82), .ZN(n422) );
  XNOR2_X1 U492 ( .A(n423), .B(n422), .ZN(n436) );
  XOR2_X1 U493 ( .A(KEYINPUT83), .B(G190GAT), .Z(n425) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(G99GAT), .ZN(n424) );
  XNOR2_X1 U495 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U496 ( .A(n427), .B(n426), .Z(n431) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U498 ( .A(n432), .B(KEYINPUT20), .ZN(n433) );
  XNOR2_X1 U499 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U500 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U501 ( .A(n439), .B(KEYINPUT23), .Z(n442) );
  XNOR2_X1 U502 ( .A(n440), .B(KEYINPUT22), .ZN(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n453) );
  XOR2_X1 U505 ( .A(KEYINPUT88), .B(KEYINPUT24), .Z(n446) );
  NAND2_X1 U506 ( .A1(G228GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U508 ( .A(n447), .B(G204GAT), .Z(n451) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n453), .B(n452), .ZN(n561) );
  NOR2_X1 U512 ( .A1(n563), .A2(n561), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n455), .B(n454), .ZN(n548) );
  NAND2_X1 U514 ( .A1(n560), .A2(n548), .ZN(n588) );
  INV_X1 U515 ( .A(n588), .ZN(n585) );
  NAND2_X1 U516 ( .A1(n585), .A2(n566), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U518 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n459) );
  NAND2_X1 U519 ( .A1(n520), .A2(n563), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n462), .A2(n561), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n520), .B(KEYINPUT27), .ZN(n469) );
  NAND2_X1 U522 ( .A1(n548), .A2(n469), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U524 ( .A(KEYINPUT94), .B(n467), .Z(n468) );
  NOR2_X1 U525 ( .A1(n517), .A2(n468), .ZN(n474) );
  NAND2_X1 U526 ( .A1(n469), .A2(n517), .ZN(n470) );
  XNOR2_X1 U527 ( .A(n470), .B(KEYINPUT91), .ZN(n547) );
  XNOR2_X1 U528 ( .A(n561), .B(KEYINPUT66), .ZN(n471) );
  XOR2_X1 U529 ( .A(n471), .B(KEYINPUT28), .Z(n525) );
  INV_X1 U530 ( .A(n525), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n547), .A2(n472), .ZN(n529) );
  NOR2_X1 U532 ( .A1(n563), .A2(n529), .ZN(n473) );
  NOR2_X1 U533 ( .A1(n474), .A2(n473), .ZN(n483) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT99), .ZN(n476) );
  NOR2_X1 U535 ( .A1(n589), .A2(n476), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n477), .B(KEYINPUT37), .ZN(n516) );
  NAND2_X1 U537 ( .A1(n566), .A2(n580), .ZN(n486) );
  NOR2_X1 U538 ( .A1(n516), .A2(n486), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(KEYINPUT38), .ZN(n503) );
  NAND2_X1 U540 ( .A1(n520), .A2(n503), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n479) );
  NOR2_X1 U542 ( .A1(n538), .A2(n576), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(KEYINPUT16), .ZN(n485) );
  INV_X1 U544 ( .A(n483), .ZN(n484) );
  NAND2_X1 U545 ( .A1(n485), .A2(n484), .ZN(n506) );
  NOR2_X1 U546 ( .A1(n486), .A2(n506), .ZN(n495) );
  NAND2_X1 U547 ( .A1(n517), .A2(n495), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(KEYINPUT34), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n490) );
  NAND2_X1 U551 ( .A1(n495), .A2(n520), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U553 ( .A(G8GAT), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT35), .B(KEYINPUT97), .Z(n493) );
  NAND2_X1 U555 ( .A1(n495), .A2(n563), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U557 ( .A(G15GAT), .B(n494), .Z(G1326GAT) );
  NAND2_X1 U558 ( .A1(n525), .A2(n495), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  NAND2_X1 U561 ( .A1(n503), .A2(n517), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n502) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n500) );
  NAND2_X1 U565 ( .A1(n503), .A2(n563), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n503), .A2(n525), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n504), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n508) );
  NAND2_X1 U571 ( .A1(n531), .A2(n505), .ZN(n515) );
  NOR2_X1 U572 ( .A1(n515), .A2(n506), .ZN(n511) );
  NAND2_X1 U573 ( .A1(n511), .A2(n517), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n511), .A2(n520), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n511), .A2(n563), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT43), .B(KEYINPUT104), .Z(n513) );
  NAND2_X1 U580 ( .A1(n511), .A2(n525), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(n514), .ZN(G1335GAT) );
  XOR2_X1 U583 ( .A(G85GAT), .B(KEYINPUT105), .Z(n519) );
  NOR2_X1 U584 ( .A1(n516), .A2(n515), .ZN(n524) );
  NAND2_X1 U585 ( .A1(n524), .A2(n517), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n524), .A2(n520), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n524), .A2(n563), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n522), .B(KEYINPUT106), .ZN(n523) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n523), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n528), .A2(n529), .ZN(n530) );
  NAND2_X1 U596 ( .A1(n563), .A2(n530), .ZN(n542) );
  NOR2_X1 U597 ( .A1(n531), .A2(n542), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(KEYINPUT109), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  NOR2_X1 U600 ( .A1(n351), .A2(n542), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT110), .Z(n537) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(KEYINPUT111), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n540) );
  NOR2_X1 U606 ( .A1(n538), .A2(n542), .ZN(n539) );
  XOR2_X1 U607 ( .A(n540), .B(n539), .Z(G1342GAT) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n544) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT113), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U614 ( .A1(n549), .A2(n528), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(KEYINPUT114), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n558), .A2(n566), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT52), .B(KEYINPUT115), .Z(n553) );
  NAND2_X1 U619 ( .A1(n558), .A2(n505), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT53), .Z(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n586), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT116), .ZN(n557) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n558), .A2(n576), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT55), .B(n562), .ZN(n564) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n577), .A2(n566), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n569) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT56), .B(n570), .Z(n572) );
  NAND2_X1 U637 ( .A1(n577), .A2(n505), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1349GAT) );
  NAND2_X1 U639 ( .A1(n586), .A2(n577), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U641 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(KEYINPUT122), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT123), .B(n575), .Z(n579) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1351GAT) );
  NOR2_X1 U646 ( .A1(n588), .A2(n580), .ZN(n584) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n582) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

