//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n209), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(new_n203), .A3(new_n207), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT71), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n208), .A2(new_n209), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(KEYINPUT71), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n210), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G226gat), .A2(G233gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(KEYINPUT29), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  XOR2_X1   g021(.A(KEYINPUT66), .B(G190gat), .Z(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT27), .B(G183gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT28), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT28), .ZN(new_n230));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  AND4_X1   g035(.A1(new_n222), .A2(new_n229), .A3(new_n230), .A4(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(KEYINPUT23), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n222), .A2(KEYINPUT24), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(G183gat), .A3(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G183gat), .ZN(new_n245));
  INV_X1    g044(.A(G190gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI22_X1  g046(.A1(KEYINPUT65), .A2(new_n240), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n231), .B1(KEYINPUT23), .B2(new_n234), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n239), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n238), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n239), .A2(KEYINPUT25), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n223), .A2(new_n245), .ZN(new_n254));
  AOI211_X1 g053(.A(new_n249), .B(new_n253), .C1(new_n254), .C2(new_n244), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n237), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT73), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n237), .A2(new_n256), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT73), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n221), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n257), .A2(new_n218), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n217), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n219), .A3(new_n261), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n212), .A2(new_n213), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n215), .A2(KEYINPUT71), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n266), .A2(new_n267), .B1(new_n209), .B2(new_n208), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n257), .A2(new_n218), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n265), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G64gat), .B(G92gat), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n273), .B(new_n274), .Z(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n264), .A2(KEYINPUT30), .A3(new_n271), .A4(new_n275), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n271), .A3(new_n275), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT69), .B(G113gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G120gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n285), .A2(new_n286), .B1(G113gat), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n286), .B2(new_n285), .ZN(new_n289));
  XOR2_X1   g088(.A(G127gat), .B(G134gat), .Z(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(KEYINPUT1), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G113gat), .B(G120gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n290), .B1(KEYINPUT1), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT68), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n297), .B1(new_n300), .B2(KEYINPUT2), .ZN(new_n301));
  INV_X1    g100(.A(G148gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G141gat), .ZN(new_n303));
  INV_X1    g102(.A(G141gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G148gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT75), .B1(new_n304), .B2(G148gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n301), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n305), .A2(new_n303), .B1(KEYINPUT2), .B2(new_n297), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n300), .A2(new_n297), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(KEYINPUT74), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(KEYINPUT74), .B2(new_n313), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n296), .B(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n283), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n296), .A2(new_n316), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT4), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(new_n296), .B2(new_n316), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n321), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n328), .A3(new_n315), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n296), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n321), .A2(KEYINPUT4), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n330), .B(new_n318), .C1(new_n322), .C2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n320), .B1(new_n326), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n323), .A2(new_n325), .A3(new_n330), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n283), .A2(new_n318), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT0), .ZN(new_n338));
  XNOR2_X1  g137(.A(G57gat), .B(G85gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  NAND3_X1  g139(.A1(new_n333), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT6), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n340), .B1(new_n333), .B2(new_n336), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI211_X1 g144(.A(new_n342), .B(new_n340), .C1(new_n333), .C2(new_n336), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n279), .B(new_n282), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G22gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT84), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n268), .B2(KEYINPUT29), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT29), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n217), .A2(KEYINPUT84), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n352), .A3(new_n328), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n316), .ZN(new_n354));
  AND2_X1   g153(.A1(G228gat), .A2(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n329), .A2(new_n269), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(new_n268), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n354), .A2(KEYINPUT85), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT85), .B1(new_n354), .B2(new_n358), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n268), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n214), .B2(new_n216), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n266), .A2(KEYINPUT81), .A3(new_n267), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n210), .B(KEYINPUT82), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT3), .B1(new_n366), .B2(new_n269), .ZN(new_n367));
  INV_X1    g166(.A(new_n316), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n361), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n369), .A2(new_n370), .A3(new_n356), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n370), .B1(new_n369), .B2(new_n356), .ZN(new_n372));
  OAI221_X1 g171(.A(new_n348), .B1(new_n359), .B2(new_n360), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G78gat), .B(G106gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT79), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT31), .B(G50gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  OAI22_X1  g178(.A1(new_n371), .A2(new_n372), .B1(new_n360), .B2(new_n359), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G22gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT87), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(KEYINPUT87), .A3(G22gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n379), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n373), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n377), .B(KEYINPUT80), .Z(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT86), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT86), .ZN(new_n390));
  AOI211_X1 g189(.A(new_n390), .B(new_n387), .C1(new_n381), .C2(new_n373), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n347), .B(new_n385), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT88), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n260), .A2(new_n296), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n260), .A2(new_n296), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n394), .A2(G227gat), .A3(G233gat), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT32), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n395), .ZN(new_n399));
  NAND2_X1  g198(.A1(G227gat), .A2(G233gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT34), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT34), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n403), .A3(new_n400), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT33), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n396), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G15gat), .B(G43gat), .Z(new_n407));
  XNOR2_X1  g206(.A(G71gat), .B(G99gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n402), .B(new_n404), .C1(new_n406), .C2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(new_n396), .B2(new_n405), .ZN(new_n412));
  INV_X1    g211(.A(new_n404), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n403), .B1(new_n399), .B2(new_n400), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n398), .B1(new_n411), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n411), .A2(new_n415), .A3(new_n398), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(KEYINPUT36), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT36), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n411), .A2(new_n415), .A3(new_n398), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n420), .B1(new_n421), .B2(new_n416), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n392), .A2(new_n393), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT89), .ZN(new_n426));
  INV_X1    g225(.A(new_n340), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n334), .A2(new_n319), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT39), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n368), .B(new_n296), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n430), .B2(new_n318), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n334), .A2(new_n429), .A3(new_n319), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT40), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n426), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n432), .A2(KEYINPUT89), .A3(KEYINPUT40), .A4(new_n433), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n282), .A2(new_n277), .A3(new_n278), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n344), .B1(new_n434), .B2(new_n435), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT37), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n277), .B1(new_n442), .B2(new_n275), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT38), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n272), .B2(KEYINPUT37), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n268), .B1(new_n262), .B2(new_n263), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n265), .A2(new_n217), .A3(new_n270), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(KEYINPUT37), .A3(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n448), .B(new_n276), .C1(new_n272), .C2(KEYINPUT37), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n443), .A2(new_n445), .B1(new_n449), .B2(new_n444), .ZN(new_n450));
  INV_X1    g249(.A(new_n344), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n342), .A3(new_n341), .ZN(new_n452));
  INV_X1    g251(.A(new_n346), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n280), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n441), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n389), .ZN(new_n456));
  INV_X1    g255(.A(new_n391), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n458), .B2(new_n385), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n393), .B1(new_n392), .B2(new_n423), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n425), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n385), .B1(new_n389), .B2(new_n391), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n417), .A2(KEYINPUT90), .A3(new_n418), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT90), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n421), .B2(new_n416), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n347), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT35), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n439), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n421), .A2(new_n416), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n345), .A2(new_n346), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(new_n469), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n462), .A2(new_n471), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n202), .B1(new_n461), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n459), .ZN(new_n478));
  INV_X1    g277(.A(new_n460), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n424), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n470), .A2(new_n475), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT91), .ZN(new_n482));
  XNOR2_X1  g281(.A(G113gat), .B(G141gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(G197gat), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT11), .B(G169gat), .Z(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT12), .ZN(new_n487));
  XOR2_X1   g286(.A(G15gat), .B(G22gat), .Z(new_n488));
  INV_X1    g287(.A(G1gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT16), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(G1gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G8gat), .ZN(new_n495));
  INV_X1    g294(.A(G8gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500));
  INV_X1    g299(.A(G29gat), .ZN(new_n501));
  INV_X1    g300(.A(G36gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G43gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G50gat), .ZN(new_n507));
  INV_X1    g306(.A(G50gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G43gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT15), .ZN(new_n510));
  NAND2_X1  g309(.A1(G29gat), .A2(G36gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(KEYINPUT92), .A2(G29gat), .A3(G36gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n505), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n506), .A2(KEYINPUT94), .A3(G50gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT94), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(G43gat), .B2(new_n508), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n508), .A2(G43gat), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT93), .B(KEYINPUT15), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n524), .A3(KEYINPUT95), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT94), .B1(new_n506), .B2(G50gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n507), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n522), .B1(new_n528), .B2(new_n517), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n505), .A2(new_n510), .A3(new_n515), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n505), .A2(new_n515), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(KEYINPUT15), .A3(new_n507), .A4(new_n509), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n525), .A2(new_n531), .A3(KEYINPUT17), .A4(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n499), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n525), .A2(new_n531), .A3(new_n533), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n536), .A2(new_n498), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT97), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n536), .A2(new_n498), .A3(KEYINPUT97), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n541), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT18), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n541), .A2(KEYINPUT18), .A3(new_n547), .A4(new_n542), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n536), .A2(new_n498), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n542), .B(KEYINPUT13), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND4_X1   g354(.A1(new_n487), .A2(new_n550), .A3(new_n551), .A4(new_n555), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n548), .A2(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n487), .B1(new_n557), .B2(new_n551), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n477), .A2(new_n482), .A3(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(KEYINPUT41), .ZN(new_n563));
  NAND2_X1  g362(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n566), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G99gat), .ZN(new_n569));
  INV_X1    g368(.A(G106gat), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT104), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT104), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(G99gat), .A3(G106gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(KEYINPUT8), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G99gat), .B(G106gat), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n568), .A2(new_n578), .A3(new_n574), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n534), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n536), .A2(new_n538), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT96), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n580), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n536), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n562), .A2(KEYINPUT41), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(G190gat), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n539), .A2(new_n540), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n246), .B(new_n591), .C1(new_n592), .C2(new_n581), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n590), .A2(new_n593), .A3(G218gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT103), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(G218gat), .B1(new_n590), .B2(new_n593), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n563), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  INV_X1    g398(.A(new_n563), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(new_n595), .A3(new_n600), .A4(new_n594), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G134gat), .B(G162gat), .Z(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606));
  INV_X1    g405(.A(G231gat), .ZN(new_n607));
  INV_X1    g406(.A(G233gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(G64gat), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G64gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(G57gat), .ZN(new_n614));
  INV_X1    g413(.A(G71gat), .ZN(new_n615));
  INV_X1    g414(.A(G78gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT9), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n612), .A2(new_n614), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G57gat), .B(G64gat), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT9), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n618), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n619), .A2(KEYINPUT98), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(G71gat), .B2(G78gat), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n625), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(G57gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(G64gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n614), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n617), .B1(new_n634), .B2(KEYINPUT9), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n626), .A2(new_n628), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT99), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n622), .B1(new_n631), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n630), .B1(new_n625), .B2(new_n629), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n635), .A2(KEYINPUT99), .A3(new_n636), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(KEYINPUT101), .A3(new_n622), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n609), .B1(new_n645), .B2(KEYINPUT21), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT21), .ZN(new_n647));
  INV_X1    g446(.A(new_n609), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n640), .A2(new_n647), .A3(new_n644), .A4(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(G127gat), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n650), .B1(new_n646), .B2(new_n649), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n606), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  INV_X1    g454(.A(new_n606), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n651), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n645), .A2(KEYINPUT21), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n499), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n647), .B1(new_n640), .B2(new_n644), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT102), .B1(new_n662), .B2(new_n498), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(new_n298), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n658), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n654), .A2(new_n657), .A3(new_n667), .A4(new_n668), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n598), .A2(new_n601), .A3(new_n603), .ZN(new_n673));
  XNOR2_X1  g472(.A(G120gat), .B(G148gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(G176gat), .B(G204gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(G230gat), .A2(G233gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT106), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT10), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n586), .B1(new_n640), .B2(new_n644), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n586), .A2(new_n638), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n680), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n580), .A2(new_n680), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n645), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n679), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT101), .B1(new_n643), .B2(new_n622), .ZN(new_n688));
  AOI211_X1 g487(.A(new_n639), .B(new_n621), .C1(new_n641), .C2(new_n642), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n580), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n690), .A2(G230gat), .A3(G233gat), .A4(new_n682), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n677), .B1(new_n687), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g494(.A(KEYINPUT107), .B(new_n677), .C1(new_n687), .C2(new_n692), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n691), .B(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT10), .B1(new_n690), .B2(new_n682), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n645), .A2(new_n685), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n678), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(new_n676), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n695), .A2(new_n696), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n605), .A2(new_n672), .A3(new_n673), .A4(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n561), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n473), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT109), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n561), .A2(new_n709), .A3(new_n473), .A4(new_n705), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT108), .B(G1gat), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n708), .B2(new_n710), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(G1324gat));
  NOR2_X1   g513(.A1(new_n706), .A2(new_n471), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT16), .B(G8gat), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G8gat), .B1(new_n706), .B2(new_n471), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n715), .A2(KEYINPUT42), .A3(new_n716), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(G1325gat));
  OAI21_X1  g521(.A(G15gat), .B1(new_n706), .B2(new_n423), .ZN(new_n723));
  INV_X1    g522(.A(new_n466), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n724), .A2(G15gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n706), .B2(new_n725), .ZN(G1326gat));
  NOR2_X1   g525(.A1(new_n706), .A2(new_n462), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT43), .B(G22gat), .Z(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n605), .A2(new_n673), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n672), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n703), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n477), .A2(new_n482), .A3(new_n560), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n473), .A2(new_n501), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n730), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OR3_X1    g537(.A1(new_n736), .A2(new_n730), .A3(new_n737), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n732), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n477), .A2(new_n482), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n462), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n392), .B(new_n423), .C1(new_n743), .C2(new_n455), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n470), .A3(new_n475), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n731), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n740), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n734), .A2(new_n559), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n748), .A2(new_n473), .A3(new_n749), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n738), .B(new_n739), .C1(new_n750), .C2(new_n501), .ZN(G1328gat));
  NAND3_X1  g550(.A1(new_n748), .A2(new_n439), .A3(new_n749), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G36gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n439), .A2(new_n502), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n736), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n755), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n757));
  OAI221_X1 g556(.A(new_n753), .B1(KEYINPUT110), .B2(KEYINPUT46), .C1(new_n756), .C2(new_n757), .ZN(G1329gat));
  INV_X1    g557(.A(new_n736), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n724), .A2(G43gat), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n759), .A2(new_n760), .B1(KEYINPUT111), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n423), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n742), .A2(new_n763), .A3(new_n747), .A4(new_n749), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G43gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1330gat));
  NAND2_X1  g567(.A1(new_n743), .A2(new_n508), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT112), .Z(new_n770));
  NOR2_X1   g569(.A1(new_n736), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n742), .A2(new_n743), .A3(new_n747), .A4(new_n749), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(G50gat), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n772), .B2(G50gat), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT48), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AOI221_X4 g576(.A(new_n771), .B1(new_n774), .B2(KEYINPUT48), .C1(G50gat), .C2(new_n772), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(G1331gat));
  NOR4_X1   g578(.A1(new_n731), .A2(new_n560), .A3(new_n733), .A4(new_n703), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT114), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n745), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n473), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n610), .A2(new_n611), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1332gat));
  AOI21_X1  g585(.A(new_n471), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n788), .B(new_n789), .Z(G1333gat));
  OAI21_X1  g589(.A(G71gat), .B1(new_n782), .B2(new_n423), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n466), .A2(new_n615), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n782), .B2(new_n792), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g593(.A1(new_n782), .A2(new_n462), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(new_n616), .ZN(G1335gat));
  NOR2_X1   g595(.A1(new_n672), .A2(new_n560), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n745), .A2(new_n731), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT51), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n695), .A2(new_n696), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n702), .A2(new_n698), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n745), .A2(new_n803), .A3(new_n731), .A4(new_n797), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n799), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(G85gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n806), .A3(new_n473), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n797), .A2(new_n802), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(KEYINPUT115), .Z(new_n809));
  AND2_X1   g608(.A1(new_n748), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n473), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n811), .B2(new_n806), .ZN(G1336gat));
  NAND4_X1  g611(.A1(new_n742), .A2(new_n439), .A3(new_n747), .A4(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G92gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n805), .A2(new_n565), .A3(new_n439), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT52), .ZN(G1337gat));
  AOI21_X1  g616(.A(G99gat), .B1(new_n805), .B2(new_n466), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n423), .A2(new_n569), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n810), .B2(new_n819), .ZN(G1338gat));
  NOR2_X1   g619(.A1(KEYINPUT116), .A2(KEYINPUT53), .ZN(new_n821));
  AND2_X1   g620(.A1(KEYINPUT116), .A2(KEYINPUT53), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n742), .A2(new_n743), .A3(new_n747), .A4(new_n809), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G106gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n805), .A2(new_n570), .A3(new_n743), .ZN(new_n825));
  AOI211_X1 g624(.A(new_n821), .B(new_n822), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AND4_X1   g625(.A1(KEYINPUT116), .A2(new_n824), .A3(new_n825), .A4(KEYINPUT53), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(G1339gat));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n705), .A2(new_n829), .A3(new_n559), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT117), .B1(new_n704), .B2(new_n560), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n542), .B1(new_n541), .B2(new_n547), .ZN(new_n833));
  OAI22_X1  g632(.A1(new_n833), .A2(KEYINPUT118), .B1(new_n553), .B2(new_n554), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n833), .A2(KEYINPUT118), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n486), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n557), .A2(new_n487), .A3(new_n551), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n684), .A2(new_n686), .A3(new_n679), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n701), .A2(new_n839), .A3(KEYINPUT54), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  INV_X1    g640(.A(new_n679), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n841), .B(new_n842), .C1(new_n699), .C2(new_n700), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n677), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n801), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n676), .B1(new_n687), .B2(new_n841), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT55), .B1(new_n846), .B2(new_n840), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n838), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n731), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n801), .B(new_n844), .C1(new_n556), .C2(new_n558), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n847), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n703), .A2(new_n838), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n849), .B1(new_n853), .B2(new_n731), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n733), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n832), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n462), .A2(new_n472), .ZN(new_n858));
  NOR4_X1   g657(.A1(new_n857), .A2(new_n707), .A3(new_n439), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n284), .A3(new_n560), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n743), .A2(new_n724), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n707), .A2(new_n439), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n559), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n860), .A2(new_n865), .ZN(G1340gat));
  AOI21_X1  g665(.A(G120gat), .B1(new_n859), .B2(new_n802), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n864), .A2(new_n287), .A3(new_n703), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(G1341gat));
  NAND3_X1  g668(.A1(new_n859), .A2(new_n650), .A3(new_n672), .ZN(new_n870));
  OAI21_X1  g669(.A(G127gat), .B1(new_n864), .B2(new_n733), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1342gat));
  INV_X1    g671(.A(G134gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n859), .A2(new_n873), .A3(new_n731), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n864), .B2(new_n732), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1343gat));
  NAND2_X1  g677(.A1(new_n743), .A2(new_n423), .ZN(new_n879));
  NOR4_X1   g678(.A1(new_n857), .A2(new_n707), .A3(new_n439), .A4(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n560), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n423), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT119), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n885), .B1(new_n857), .B2(new_n462), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n830), .A2(new_n831), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n846), .A2(new_n840), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT55), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT120), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n891), .B(KEYINPUT55), .C1(new_n846), .C2(new_n840), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n850), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT121), .B1(new_n893), .B2(new_n852), .ZN(new_n894));
  INV_X1    g693(.A(new_n838), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n802), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n847), .B(KEYINPUT120), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n896), .B(new_n897), .C1(new_n898), .C2(new_n850), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n894), .A2(new_n732), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n672), .B1(new_n900), .B2(new_n849), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT57), .B(new_n743), .C1(new_n887), .C2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n884), .B1(new_n886), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n559), .A2(new_n304), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n881), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n302), .A2(KEYINPUT59), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n903), .B2(new_n802), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n743), .A2(KEYINPUT57), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n832), .B2(new_n855), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n704), .A2(new_n560), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n743), .B1(new_n901), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n911), .B1(new_n913), .B2(new_n885), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n883), .A2(new_n802), .ZN(new_n915));
  OAI21_X1  g714(.A(G148gat), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT59), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT122), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT59), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n909), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n880), .A2(new_n302), .A3(new_n802), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n907), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT59), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n919), .B1(new_n916), .B2(KEYINPUT59), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g726(.A(KEYINPUT123), .B(new_n922), .C1(new_n927), .C2(new_n909), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n924), .A2(new_n928), .ZN(G1345gat));
  AOI21_X1  g728(.A(G155gat), .B1(new_n880), .B2(new_n672), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n672), .A2(G155gat), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT124), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n903), .B2(new_n932), .ZN(G1346gat));
  AOI21_X1  g732(.A(G162gat), .B1(new_n880), .B2(new_n731), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n732), .A2(new_n299), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n903), .B2(new_n935), .ZN(G1347gat));
  NOR4_X1   g735(.A1(new_n857), .A2(new_n473), .A3(new_n471), .A4(new_n858), .ZN(new_n937));
  AOI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n560), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n473), .A2(new_n471), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n862), .A2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n560), .A2(G169gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1348gat));
  INV_X1    g741(.A(G176gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n937), .A2(new_n943), .A3(new_n802), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n940), .A2(new_n802), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n943), .ZN(G1349gat));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n856), .A2(new_n861), .A3(new_n672), .A4(new_n939), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n245), .B1(new_n948), .B2(KEYINPUT125), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n949), .B1(KEYINPUT125), .B2(new_n948), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n937), .A2(new_n224), .A3(new_n672), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(new_n951), .A3(new_n947), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  AOI22_X1  g754(.A1(new_n953), .A2(new_n954), .B1(new_n955), .B2(KEYINPUT60), .ZN(new_n956));
  INV_X1    g755(.A(new_n954), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(KEYINPUT60), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n957), .A2(new_n958), .A3(new_n952), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n956), .A2(new_n959), .ZN(G1350gat));
  AOI21_X1  g759(.A(new_n246), .B1(new_n940), .B2(new_n731), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT61), .Z(new_n962));
  NAND3_X1  g761(.A1(new_n937), .A2(new_n223), .A3(new_n731), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1351gat));
  NOR4_X1   g763(.A1(new_n857), .A2(new_n473), .A3(new_n471), .A4(new_n879), .ZN(new_n965));
  AOI21_X1  g764(.A(G197gat), .B1(new_n965), .B2(new_n560), .ZN(new_n966));
  NOR4_X1   g765(.A1(new_n914), .A2(new_n473), .A3(new_n471), .A4(new_n763), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n560), .A2(G197gat), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(G1352gat));
  INV_X1    g768(.A(G204gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n965), .A2(new_n970), .A3(new_n802), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT62), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n970), .B1(new_n967), .B2(new_n802), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n972), .A2(new_n973), .ZN(G1353gat));
  NAND3_X1  g773(.A1(new_n965), .A2(new_n205), .A3(new_n672), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n967), .A2(new_n672), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  NAND3_X1  g778(.A1(new_n965), .A2(new_n206), .A3(new_n731), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n967), .A2(new_n731), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n981), .B2(new_n206), .ZN(G1355gat));
endmodule


