//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n210));
  XNOR2_X1  g0010(.A(new_n209), .B(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n207), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  AND2_X1   g0022(.A1(KEYINPUT65), .A2(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(KEYINPUT65), .A2(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n202), .A2(new_n203), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n211), .B(new_n222), .C1(new_n227), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  OAI211_X1 g0049(.A(new_n249), .B(G274), .C1(G41), .C2(G45), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT67), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G226), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(G1), .B(G13), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n252), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n254), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(KEYINPUT68), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G222), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(G223), .A3(G1698), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n270), .B(new_n271), .C1(new_n213), .C2(new_n268), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n259), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G200), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT74), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT65), .ZN(new_n278));
  INV_X1    g0078(.A(G20), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT65), .A2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT71), .B1(new_n282), .B2(new_n254), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT71), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n225), .A2(new_n284), .A3(G33), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT8), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT70), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n202), .ZN(new_n288));
  NAND3_X1  g0088(.A1(KEYINPUT70), .A2(KEYINPUT8), .A3(G58), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n283), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n279), .A2(new_n254), .A3(KEYINPUT72), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT72), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(G20), .B2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n295), .A2(G150), .B1(G20), .B2(new_n204), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT69), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT69), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n300), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n226), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G50), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n302), .B1(new_n249), .B2(G20), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(G50), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT9), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n274), .A2(G190), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(KEYINPUT9), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n277), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(new_n277), .B2(new_n313), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n274), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n308), .B1(new_n274), .B2(G169), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT76), .ZN(new_n323));
  INV_X1    g0123(.A(new_n302), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n283), .A2(G77), .A3(new_n285), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n295), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT12), .B1(new_n304), .B2(G68), .ZN(new_n329));
  OR3_X1    g0129(.A1(new_n304), .A2(KEYINPUT12), .A3(G68), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n306), .A2(G68), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n325), .A2(new_n326), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n302), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT11), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n338), .A2(KEYINPUT76), .A3(new_n328), .A4(new_n331), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n263), .A2(new_n267), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n233), .A2(G1698), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(G226), .B2(G1698), .ZN(new_n344));
  INV_X1    g0144(.A(G97), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n342), .A2(new_n344), .B1(new_n254), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n273), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT75), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n256), .A2(G238), .A3(new_n257), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n252), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n348), .B1(new_n252), .B2(new_n349), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT13), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n347), .B(new_n354), .C1(new_n350), .C2(new_n351), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n357), .A3(G169), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(G179), .A3(new_n355), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n357), .B1(new_n356), .B2(G169), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n341), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n275), .B1(new_n353), .B2(new_n355), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n353), .A2(new_n355), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(G190), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT77), .B1(new_n365), .B2(new_n340), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n353), .A2(G190), .A3(new_n355), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n356), .A2(G200), .ZN(new_n368));
  AND4_X1   g0168(.A1(KEYINPUT77), .A2(new_n340), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n362), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n288), .B(new_n289), .C1(G1), .C2(new_n279), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n299), .A2(new_n301), .A3(new_n226), .A4(new_n304), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n372), .A2(new_n373), .B1(new_n290), .B2(new_n304), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n265), .A2(new_n266), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT7), .B1(new_n376), .B2(G20), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n261), .A2(new_n262), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n225), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n377), .A2(new_n380), .A3(G68), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n295), .A2(G159), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n279), .B1(new_n228), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT78), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G159), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n292), .B2(new_n294), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT78), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n388), .A2(new_n384), .A3(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT16), .B(new_n381), .C1(new_n386), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n302), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n280), .A2(new_n265), .A3(new_n281), .A4(new_n266), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT7), .ZN(new_n394));
  NOR2_X1   g0194(.A1(KEYINPUT7), .A2(G20), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(G68), .B(new_n394), .C1(new_n268), .C2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n388), .A2(new_n384), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT16), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n375), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n256), .A2(G232), .A3(new_n257), .ZN(new_n401));
  INV_X1    g0201(.A(G45), .ZN(new_n402));
  AOI21_X1  g0202(.A(G1), .B1(new_n255), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT67), .B1(new_n403), .B2(G274), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n250), .A2(new_n251), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(G226), .A2(G1698), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n261), .B2(new_n262), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT80), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  OAI211_X1 g0211(.A(G223), .B(new_n269), .C1(new_n261), .C2(new_n262), .ZN(new_n412));
  OAI211_X1 g0212(.A(KEYINPUT80), .B(new_n407), .C1(new_n261), .C2(new_n262), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n410), .A2(new_n411), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  AOI211_X1 g0214(.A(G179), .B(new_n406), .C1(new_n273), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n273), .ZN(new_n416));
  INV_X1    g0216(.A(new_n406), .ZN(new_n417));
  AOI21_X1  g0217(.A(G169), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT81), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n318), .A3(new_n417), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT81), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n406), .B1(new_n414), .B2(new_n273), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n420), .B(new_n421), .C1(G169), .C2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n400), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT18), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n400), .A2(new_n419), .A3(new_n426), .A4(new_n423), .ZN(new_n427));
  INV_X1    g0227(.A(new_n398), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n342), .A2(new_n395), .B1(KEYINPUT7), .B2(new_n393), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(G68), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n391), .B(new_n302), .C1(new_n430), .C2(KEYINPUT16), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n422), .A2(new_n275), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n422), .A2(G190), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n431), .A2(new_n433), .A3(new_n375), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT17), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n432), .B1(G190), .B2(new_n422), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n438), .A2(KEYINPUT17), .A3(new_n375), .A4(new_n431), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n425), .A2(new_n427), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n306), .A2(G77), .ZN(new_n442));
  INV_X1    g0242(.A(new_n304), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT73), .B1(new_n443), .B2(new_n213), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n443), .A2(KEYINPUT73), .A3(new_n213), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  XOR2_X1   g0246(.A(KEYINPUT8), .B(G58), .Z(new_n447));
  AOI22_X1  g0247(.A1(new_n447), .A2(new_n295), .B1(new_n282), .B2(G77), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT15), .B(G87), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(G33), .A3(new_n225), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n324), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n256), .B1(new_n342), .B2(new_n215), .ZN(new_n455));
  MUX2_X1   g0255(.A(G232), .B(G238), .S(G1698), .Z(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n342), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(new_n252), .C1(new_n214), .C2(new_n258), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n454), .B1(G200), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G190), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(new_n458), .ZN(new_n461));
  INV_X1    g0261(.A(G169), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n453), .B1(new_n462), .B2(new_n458), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(G179), .B2(new_n458), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n322), .A2(new_n371), .A3(new_n441), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n304), .A2(G116), .ZN(new_n468));
  INV_X1    g0268(.A(G116), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G20), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n254), .A2(G97), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G283), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n280), .A2(new_n471), .A3(new_n281), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n302), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT20), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n302), .A2(KEYINPUT20), .A3(new_n473), .A4(new_n470), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n468), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(G1), .A2(G13), .ZN(new_n479));
  AND3_X1   g0279(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(new_n300), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n254), .A2(G1), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n481), .A2(new_n299), .A3(new_n304), .A4(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT89), .B1(new_n484), .B2(new_n469), .ZN(new_n485));
  INV_X1    g0285(.A(new_n373), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT89), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(G116), .A4(new_n483), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT90), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n478), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n478), .B2(new_n489), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n216), .A2(G1698), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n376), .B(new_n494), .C1(G257), .C2(G1698), .ZN(new_n495));
  INV_X1    g0295(.A(G303), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n268), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G274), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n273), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT5), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(G41), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n501), .A2(KEYINPUT86), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n249), .A2(G45), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n500), .B2(G41), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(KEYINPUT86), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n497), .A2(new_n273), .B1(new_n499), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n402), .A2(G1), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(KEYINPUT5), .B2(new_n255), .ZN(new_n509));
  OAI211_X1 g0309(.A(G270), .B(new_n256), .C1(new_n509), .C2(new_n501), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT88), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G200), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n493), .B(new_n514), .C1(new_n460), .C2(new_n513), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n462), .B1(new_n507), .B2(new_n512), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n491), .B2(new_n492), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT21), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(KEYINPUT21), .B(new_n516), .C1(new_n491), .C2(new_n492), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n513), .A2(new_n318), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n491), .B2(new_n492), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n515), .A2(new_n519), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n503), .A2(G250), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n273), .A2(new_n524), .B1(new_n498), .B2(new_n503), .ZN(new_n525));
  OAI211_X1 g0325(.A(G244), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n526));
  OAI211_X1 g0326(.A(G238), .B(new_n269), .C1(new_n261), .C2(new_n262), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n526), .B(new_n527), .C1(new_n254), .C2(new_n469), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n525), .B1(new_n528), .B2(new_n273), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G179), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n462), .B2(new_n529), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n280), .A2(G33), .A3(G97), .A4(new_n281), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n376), .A2(new_n225), .A3(G68), .ZN(new_n535));
  NAND3_X1  g0335(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n280), .A2(new_n281), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G87), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(new_n345), .A3(new_n215), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n534), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n302), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n449), .A2(new_n443), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n373), .A2(new_n482), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n450), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT87), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n541), .A2(new_n302), .B1(new_n443), .B2(new_n449), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT87), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n549), .A3(new_n545), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n531), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n528), .A2(new_n273), .ZN(new_n552));
  INV_X1    g0352(.A(new_n525), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G200), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n529), .A2(G190), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n544), .A2(G87), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n548), .A4(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n443), .A2(new_n215), .ZN(new_n560));
  XOR2_X1   g0360(.A(new_n560), .B(KEYINPUT25), .Z(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n215), .B2(new_n484), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n282), .A2(new_n563), .B1(KEYINPUT23), .B2(G107), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n254), .A2(new_n469), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n279), .B1(new_n565), .B2(KEYINPUT23), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n342), .B2(new_n538), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n376), .A2(new_n225), .A3(KEYINPUT22), .A4(G87), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT24), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n567), .A2(new_n573), .A3(new_n569), .A4(new_n570), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n562), .B1(new_n575), .B2(new_n302), .ZN(new_n576));
  INV_X1    g0376(.A(G257), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G1698), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(G250), .B2(G1698), .ZN(new_n579));
  XNOR2_X1  g0379(.A(KEYINPUT91), .B(G294), .ZN(new_n580));
  OAI22_X1  g0380(.A1(new_n579), .A2(new_n378), .B1(new_n580), .B2(new_n254), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n273), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n499), .A2(new_n504), .A3(new_n505), .A4(new_n502), .ZN(new_n583));
  OAI211_X1 g0383(.A(G264), .B(new_n256), .C1(new_n509), .C2(new_n501), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n275), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT92), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT92), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n588), .A3(new_n275), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n587), .B(new_n589), .C1(G190), .C2(new_n585), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n576), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n585), .A2(G179), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n462), .B2(new_n585), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n324), .B1(new_n572), .B2(new_n574), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(new_n562), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n559), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT85), .B1(new_n429), .B2(G107), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n396), .B1(new_n263), .B2(new_n267), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n379), .B1(new_n225), .B2(new_n378), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT85), .ZN(new_n600));
  NOR4_X1   g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n215), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n215), .A2(G97), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT83), .ZN(new_n604));
  AND2_X1   g0404(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n605));
  NOR2_X1   g0405(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n345), .A2(G107), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OR2_X1    g0409(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n610));
  NAND2_X1  g0410(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n611));
  AND4_X1   g0411(.A1(new_n604), .A2(new_n610), .A3(new_n608), .A4(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n603), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n608), .A3(new_n611), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT83), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n607), .A2(new_n604), .A3(new_n608), .ZN(new_n616));
  INV_X1    g0416(.A(new_n603), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n613), .A2(new_n618), .A3(new_n282), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT84), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n295), .A2(G77), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n602), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n620), .B1(new_n619), .B2(new_n621), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n302), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n304), .A2(G97), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n544), .B2(G97), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n256), .B1(new_n509), .B2(new_n501), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n583), .B1(new_n577), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n376), .A2(G244), .A3(new_n269), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT4), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n263), .A2(new_n267), .A3(G250), .A4(G1698), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n632), .A2(new_n214), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n263), .A2(new_n267), .A3(new_n269), .A4(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n633), .A2(new_n634), .A3(new_n636), .A4(new_n472), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n273), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n630), .A2(new_n638), .A3(new_n460), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n629), .B1(new_n273), .B2(new_n637), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n639), .B1(new_n640), .B2(G200), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n625), .A2(new_n627), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n630), .A2(new_n638), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n462), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n630), .A2(new_n638), .A3(new_n318), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n625), .B2(new_n627), .ZN(new_n647));
  NOR4_X1   g0447(.A1(new_n523), .A2(new_n596), .A3(new_n642), .A4(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n467), .A2(new_n648), .ZN(G372));
  NAND2_X1  g0449(.A1(new_n437), .A2(new_n439), .ZN(new_n650));
  INV_X1    g0450(.A(new_n464), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n366), .B2(new_n369), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n650), .B1(new_n652), .B2(new_n362), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n425), .A2(new_n427), .ZN(new_n654));
  OAI22_X1  g0454(.A1(new_n653), .A2(new_n654), .B1(new_n316), .B2(new_n315), .ZN(new_n655));
  INV_X1    g0455(.A(new_n321), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n655), .A2(KEYINPUT93), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT93), .B1(new_n655), .B2(new_n656), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n647), .A2(new_n559), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(KEYINPUT26), .B1(new_n531), .B2(new_n546), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n519), .A2(new_n595), .A3(new_n520), .A4(new_n522), .ZN(new_n662));
  INV_X1    g0462(.A(new_n647), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n625), .A2(new_n627), .A3(new_n641), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n529), .A2(new_n462), .ZN(new_n665));
  AOI211_X1 g0465(.A(new_n318), .B(new_n525), .C1(new_n528), .C2(new_n273), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n546), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n558), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n576), .B2(new_n590), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n662), .A2(new_n663), .A3(new_n664), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n625), .A2(new_n627), .ZN(new_n671));
  INV_X1    g0471(.A(new_n646), .ZN(new_n672));
  INV_X1    g0472(.A(new_n668), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n671), .A2(new_n672), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n661), .A2(new_n670), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n467), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n659), .A2(new_n677), .ZN(G369));
  INV_X1    g0478(.A(KEYINPUT95), .ZN(new_n679));
  INV_X1    g0479(.A(new_n493), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n225), .A2(new_n249), .A3(G13), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT94), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n523), .B2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  INV_X1    g0493(.A(new_n595), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n686), .B1(new_n594), .B2(new_n562), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n591), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n595), .A2(new_n686), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n679), .B1(new_n693), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n692), .A2(KEYINPUT95), .A3(G330), .A4(new_n698), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n686), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n690), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n697), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n208), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n539), .A2(G116), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n229), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  INV_X1    g0516(.A(new_n627), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n619), .A2(new_n621), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT84), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(new_n622), .A3(new_n602), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n717), .B1(new_n720), .B2(new_n302), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n664), .B(new_n669), .C1(new_n721), .C2(new_n646), .ZN(new_n722));
  AND4_X1   g0522(.A1(new_n519), .A2(new_n520), .A3(new_n595), .A4(new_n522), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n551), .A2(new_n558), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n721), .A2(new_n646), .A3(new_n725), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n675), .B(new_n667), .C1(new_n726), .C2(new_n674), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n703), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT97), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT97), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n728), .A2(new_n732), .A3(new_n729), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n671), .A2(new_n559), .A3(new_n674), .A4(new_n672), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n667), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n674), .B1(new_n647), .B2(new_n673), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT98), .B1(new_n722), .B2(new_n723), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n642), .A2(new_n647), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT98), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n739), .A2(new_n740), .A3(new_n662), .A4(new_n669), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n737), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n742), .A2(KEYINPUT29), .A3(new_n703), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n731), .A2(new_n733), .B1(new_n743), .B2(KEYINPUT99), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n742), .A2(KEYINPUT29), .A3(new_n703), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT99), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n513), .A2(new_n318), .A3(new_n554), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT96), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n643), .A2(new_n585), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n529), .A2(new_n582), .A3(new_n584), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n521), .A2(new_n640), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT30), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT30), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n751), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n686), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT31), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n749), .A2(new_n750), .B1(new_n754), .B2(KEYINPUT30), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n703), .B1(new_n762), .B2(new_n757), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n648), .B2(new_n703), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n761), .B1(new_n764), .B2(new_n760), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n744), .A2(new_n747), .B1(G330), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n716), .B1(new_n766), .B2(G1), .ZN(G364));
  AND2_X1   g0567(.A1(new_n225), .A2(G13), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G45), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G1), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n711), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n692), .B2(G330), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G330), .B2(new_n692), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n226), .B1(G20), .B2(new_n462), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G179), .A2(G200), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n282), .A2(new_n460), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT102), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(KEYINPUT102), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G329), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n225), .A2(new_n318), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n786), .A2(new_n460), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n275), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT33), .B(G317), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G322), .A2(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n789), .A2(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n787), .A2(new_n275), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G311), .A2(new_n793), .B1(new_n794), .B2(G326), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n275), .A2(G179), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n282), .A2(new_n460), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n778), .A2(G190), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n282), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n342), .B1(new_n797), .B2(new_n798), .C1(new_n801), .C2(new_n580), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n796), .A2(G20), .A3(G190), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT101), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n802), .B1(G303), .B2(new_n804), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n785), .A2(new_n792), .A3(new_n795), .A4(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G50), .A2(new_n794), .B1(new_n788), .B2(G58), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G68), .A2(new_n790), .B1(new_n793), .B2(G77), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n800), .A2(G97), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n809), .B(new_n268), .C1(new_n538), .C2(new_n803), .ZN(new_n810));
  INV_X1    g0610(.A(new_n797), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n810), .B1(G107), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n779), .A2(new_n387), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT32), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n807), .A2(new_n808), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n777), .B1(new_n806), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n342), .A2(new_n710), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G355), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(G116), .B2(new_n208), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n244), .A2(G45), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n376), .B(new_n710), .C1(new_n230), .C2(new_n402), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G13), .A2(G33), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(G20), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n776), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n771), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n816), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n825), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n692), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n774), .A2(new_n775), .A3(new_n831), .ZN(G396));
  NOR2_X1   g0632(.A1(new_n464), .A2(new_n686), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n461), .B1(new_n453), .B2(new_n703), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n464), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n728), .B(new_n835), .Z(new_n836));
  NAND2_X1  g0636(.A1(new_n765), .A2(G330), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n771), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  INV_X1    g0639(.A(new_n771), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n776), .A2(new_n823), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n213), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n804), .A2(G107), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n811), .A2(G87), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(new_n342), .A3(new_n809), .A4(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G294), .A2(new_n788), .B1(new_n794), .B2(G303), .ZN(new_n846));
  INV_X1    g0646(.A(new_n793), .ZN(new_n847));
  INV_X1    g0647(.A(new_n790), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n846), .B1(new_n469), .B2(new_n847), .C1(new_n798), .C2(new_n848), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n845), .B(new_n849), .C1(G311), .C2(new_n784), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G143), .A2(new_n788), .B1(new_n793), .B2(G159), .ZN(new_n851));
  INV_X1    g0651(.A(G137), .ZN(new_n852));
  INV_X1    g0652(.A(new_n794), .ZN(new_n853));
  INV_X1    g0653(.A(G150), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n851), .B1(new_n852), .B2(new_n853), .C1(new_n854), .C2(new_n848), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT34), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(G132), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n783), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n804), .A2(G50), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n811), .A2(G68), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n378), .B1(new_n800), .B2(G58), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n859), .B(new_n863), .C1(new_n855), .C2(new_n856), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n850), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n842), .B1(new_n865), .B2(new_n777), .C1(new_n835), .C2(new_n824), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n839), .A2(new_n866), .ZN(G384));
  NAND2_X1  g0667(.A1(new_n613), .A2(new_n618), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT103), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT35), .ZN(new_n871));
  OAI211_X1 g0671(.A(G116), .B(new_n227), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n871), .B2(new_n870), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT36), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n230), .A2(G77), .A3(new_n383), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n201), .A2(G68), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n249), .B(G13), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n731), .A2(new_n733), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n742), .A2(KEYINPUT99), .A3(KEYINPUT29), .A4(new_n703), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n879), .A2(new_n467), .A3(new_n747), .A4(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT105), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n744), .A2(KEYINPUT105), .A3(new_n467), .A4(new_n747), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n883), .A2(new_n884), .A3(new_n659), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n382), .A2(new_n385), .A3(KEYINPUT78), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n389), .B1(new_n388), .B2(new_n384), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT16), .B1(new_n888), .B2(new_n381), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n375), .B1(new_n392), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n684), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n440), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n400), .A2(new_n891), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n424), .A2(new_n895), .A3(new_n896), .A4(new_n435), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n890), .A2(new_n419), .A3(new_n423), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n898), .A2(new_n435), .A3(new_n892), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n899), .B2(new_n896), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n894), .A2(new_n900), .A3(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT104), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n440), .A2(new_n400), .A3(new_n891), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n424), .A2(new_n435), .A3(new_n895), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n897), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n906), .B1(new_n911), .B2(new_n902), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT39), .B1(new_n905), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n902), .ZN(new_n914));
  NOR2_X1   g0714(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(new_n904), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n362), .A2(new_n686), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n835), .B(new_n703), .C1(new_n724), .C2(new_n727), .ZN(new_n921));
  INV_X1    g0721(.A(new_n833), .ZN(new_n922));
  OAI221_X1 g0722(.A(new_n362), .B1(new_n340), .B2(new_n703), .C1(new_n366), .C2(new_n369), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n340), .A2(new_n703), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n370), .A2(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n921), .A2(new_n922), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n905), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n654), .A2(new_n684), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n920), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n885), .B(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(G330), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n925), .A2(new_n923), .ZN(new_n933));
  INV_X1    g0733(.A(new_n523), .ZN(new_n934));
  INV_X1    g0734(.A(new_n596), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n934), .A2(new_n739), .A3(new_n935), .A4(new_n703), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n760), .B1(new_n936), .B2(new_n759), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n763), .A2(KEYINPUT31), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n933), .B(new_n835), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n914), .A2(new_n904), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT40), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT40), .B1(new_n903), .B2(new_n904), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n765), .A2(new_n835), .A3(new_n933), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n467), .A2(new_n765), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n932), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n945), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n931), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n249), .B2(new_n768), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n931), .A2(new_n948), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n878), .B1(new_n950), .B2(new_n951), .ZN(G367));
  NAND2_X1  g0752(.A1(new_n548), .A2(new_n557), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n686), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n673), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n954), .A2(new_n667), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n739), .B1(new_n721), .B2(new_n703), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n647), .A2(new_n686), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n707), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT42), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n957), .A2(new_n595), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n686), .B1(new_n962), .B2(new_n663), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n955), .B(new_n956), .C1(new_n964), .C2(KEYINPUT106), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT106), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n955), .A2(new_n956), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(new_n961), .C2(new_n963), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT43), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT43), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n964), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n965), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(KEYINPUT107), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n973), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT107), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n975), .A2(new_n969), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n959), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n974), .A2(new_n977), .B1(new_n702), .B2(new_n978), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n978), .A2(new_n707), .A3(new_n697), .ZN(new_n980));
  XNOR2_X1  g0780(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT110), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n978), .B1(new_n983), .B2(KEYINPUT44), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(new_n985), .B2(new_n708), .ZN(new_n986));
  OR3_X1    g0786(.A1(new_n985), .A2(new_n708), .A3(new_n984), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n982), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n988), .A2(new_n700), .A3(new_n701), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n982), .A2(new_n702), .A3(new_n986), .A4(new_n987), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT111), .B1(new_n699), .B2(new_n704), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n693), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n693), .A2(new_n992), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(new_n706), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n766), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n766), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n711), .B(new_n1000), .Z(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n770), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n976), .B1(new_n975), .B2(new_n969), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n970), .A2(KEYINPUT107), .A3(new_n973), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n702), .A2(new_n978), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n979), .A2(new_n1005), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n710), .A2(new_n376), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n239), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n827), .B1(new_n710), .B2(new_n450), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n840), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G150), .A2(new_n788), .B1(new_n790), .B2(G159), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G50), .A2(new_n793), .B1(new_n794), .B2(G143), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n268), .B1(new_n202), .B2(new_n803), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G68), .B2(new_n800), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G77), .A2(new_n811), .B1(new_n780), .B2(G137), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n793), .A2(G283), .B1(G107), .B2(new_n800), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT112), .Z(new_n1022));
  NAND2_X1  g0822(.A1(new_n811), .A2(G97), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n804), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n803), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(G116), .ZN(new_n1026));
  XOR2_X1   g0826(.A(KEYINPUT114), .B(KEYINPUT46), .Z(new_n1027));
  AOI21_X1  g0827(.A(new_n376), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n780), .A2(G317), .ZN(new_n1029));
  AND4_X1   g0829(.A1(new_n1023), .A2(new_n1024), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n580), .ZN(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT113), .B(G311), .Z(new_n1032));
  AOI22_X1  g0832(.A1(new_n1031), .A2(new_n790), .B1(new_n794), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n788), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1030), .B(new_n1033), .C1(new_n496), .C2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1020), .B1(new_n1022), .B2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT47), .Z(new_n1037));
  OAI221_X1 g0837(.A(new_n1014), .B1(new_n830), .B2(new_n967), .C1(new_n1037), .C2(new_n777), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1010), .A2(new_n1038), .ZN(G387));
  OR2_X1    g0839(.A1(new_n236), .A2(new_n402), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n713), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1040), .A2(new_n1011), .B1(new_n1041), .B2(new_n817), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n447), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1043), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n447), .B2(new_n201), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n713), .B(new_n402), .C1(new_n203), .C2(new_n213), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1042), .A2(new_n1048), .B1(G107), .B2(new_n208), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n840), .B1(new_n1049), .B2(new_n826), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n698), .B2(new_n830), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n800), .A2(new_n450), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n378), .B1(new_n1025), .B2(G77), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1023), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G150), .B2(new_n780), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G68), .A2(new_n793), .B1(new_n794), .B2(G159), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G50), .A2(new_n788), .B1(new_n790), .B2(new_n290), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n376), .B1(new_n780), .B2(G326), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n788), .A2(G317), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n790), .A2(new_n1032), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n794), .A2(G322), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n793), .A2(G303), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1065), .A2(KEYINPUT48), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(KEYINPUT48), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1031), .A2(new_n1025), .B1(new_n800), .B2(G283), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT49), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1059), .B1(new_n469), .B2(new_n797), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1058), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1051), .B1(new_n1073), .B2(new_n776), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT115), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n997), .B2(new_n770), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n998), .A2(new_n711), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n997), .A2(new_n766), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(G393));
  NAND3_X1  g0879(.A1(new_n989), .A2(new_n990), .A3(new_n770), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n826), .B1(new_n345), .B2(new_n208), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n247), .B2(new_n1011), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT116), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n800), .A2(G77), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n378), .B1(new_n1025), .B2(G68), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n844), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n201), .A2(new_n848), .B1(new_n847), .B2(new_n1043), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(G143), .C2(new_n780), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G150), .A2(new_n794), .B1(new_n788), .B2(G159), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT51), .Z(new_n1090));
  AOI22_X1  g0890(.A1(G311), .A2(new_n788), .B1(new_n794), .B2(G317), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT52), .Z(new_n1092));
  AOI22_X1  g0892(.A1(G294), .A2(new_n793), .B1(new_n790), .B2(G303), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n342), .B1(new_n798), .B2(new_n803), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G116), .B2(new_n800), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G107), .A2(new_n811), .B1(new_n780), .B2(G322), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1088), .A2(new_n1090), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n771), .B(new_n1083), .C1(new_n1098), .C2(new_n777), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT117), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n830), .B2(new_n959), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1080), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT118), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n991), .A2(new_n998), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n991), .A2(new_n998), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n711), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1103), .A2(new_n1106), .ZN(G390));
  NAND3_X1  g0907(.A1(new_n467), .A2(G330), .A3(new_n765), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n765), .A2(G330), .A3(new_n835), .A4(new_n933), .ZN(new_n1109));
  OAI211_X1 g0909(.A(G330), .B(new_n835), .C1(new_n937), .C2(new_n938), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n925), .A2(new_n923), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n834), .A2(new_n464), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n742), .A2(new_n703), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n922), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1109), .A2(new_n1112), .A3(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1109), .A2(new_n1112), .B1(new_n922), .B2(new_n921), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n885), .A2(new_n1108), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n921), .A2(new_n922), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n919), .B1(new_n1121), .B2(new_n933), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1111), .B1(new_n1114), .B2(new_n922), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n940), .A2(new_n918), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n917), .A2(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1109), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1115), .A2(new_n933), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1124), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n913), .B(new_n916), .C1(new_n926), .C2(new_n919), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1109), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1120), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1109), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n885), .A2(new_n1137), .A3(new_n1119), .A4(new_n1108), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1134), .A2(new_n711), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n841), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1034), .A2(new_n858), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n852), .A2(new_n848), .B1(new_n847), .B2(new_n1142), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1141), .B(new_n1143), .C1(G128), .C2(new_n794), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n803), .A2(new_n854), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n342), .B1(G159), .B2(new_n800), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n201), .C2(new_n797), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G125), .B2(new_n784), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n469), .A2(new_n1034), .B1(new_n853), .B2(new_n798), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n345), .A2(new_n847), .B1(new_n848), .B2(new_n215), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n804), .A2(G87), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1153), .A2(new_n342), .A3(new_n861), .A4(new_n1084), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G294), .B2(new_n784), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1144), .A2(new_n1149), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n771), .B1(new_n290), .B2(new_n1140), .C1(new_n1156), .C2(new_n777), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n917), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n823), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1137), .A2(KEYINPUT119), .A3(new_n770), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT119), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n1133), .B2(new_n1004), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1159), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1139), .A2(new_n1163), .ZN(G378));
  OAI211_X1 g0964(.A(new_n308), .B(new_n891), .C1(new_n317), .C2(new_n321), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n656), .B1(new_n309), .B2(new_n684), .C1(new_n315), .C2(new_n316), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1167), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n945), .A2(G330), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n945), .B2(G330), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n929), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n765), .A2(new_n835), .A3(new_n933), .A4(new_n940), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n939), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1175), .A2(KEYINPUT40), .B1(new_n1176), .B2(new_n943), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1170), .B1(new_n1177), .B2(new_n932), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n945), .A2(new_n1171), .A3(G330), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n930), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1174), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1170), .A2(new_n823), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n771), .B1(G50), .B2(new_n1140), .ZN(new_n1184));
  AOI21_X1  g0984(.A(G50), .B1(new_n266), .B2(new_n255), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n794), .A2(G116), .B1(G68), .B2(new_n800), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT120), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n345), .A2(new_n848), .B1(new_n1034), .B2(new_n215), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n811), .A2(G58), .ZN(new_n1189));
  AOI211_X1 g0989(.A(G41), .B(new_n376), .C1(new_n1025), .C2(G77), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n847), .C2(new_n449), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1187), .B(new_n1192), .C1(new_n798), .C2(new_n783), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT58), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1185), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n801), .A2(new_n854), .B1(new_n803), .B2(new_n1142), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G128), .A2(new_n788), .B1(new_n793), .B2(G137), .ZN(new_n1197));
  INV_X1    g0997(.A(G125), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n853), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1196), .B(new_n1199), .C1(G132), .C2(new_n790), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n811), .A2(G159), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n780), .C2(G124), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1195), .B1(new_n1194), .B2(new_n1193), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(KEYINPUT121), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n777), .B1(new_n1207), .B2(KEYINPUT121), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1184), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1182), .A2(new_n770), .B1(new_n1183), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT123), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n883), .A2(new_n884), .A3(new_n659), .A4(new_n1108), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT122), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n657), .A2(new_n658), .ZN(new_n1215));
  AOI211_X1 g1015(.A(KEYINPUT97), .B(KEYINPUT29), .C1(new_n676), .C2(new_n703), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n732), .B1(new_n728), .B2(new_n729), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n880), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n745), .A2(new_n746), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1218), .A2(new_n1219), .A3(new_n466), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1215), .B1(new_n1220), .B2(KEYINPUT105), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT122), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1221), .A2(new_n1222), .A3(new_n883), .A4(new_n1108), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1214), .A2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1213), .A2(new_n1133), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1212), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1138), .A2(KEYINPUT123), .A3(new_n1214), .A4(new_n1223), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT57), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT124), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n929), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT124), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1230), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1229), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n711), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1229), .B2(new_n1182), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1211), .B1(new_n1237), .B2(new_n1238), .ZN(G375));
  NAND2_X1  g1039(.A1(new_n1213), .A2(new_n1225), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1120), .A2(new_n1002), .A3(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n771), .B1(G68), .B2(new_n1140), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n784), .A2(G128), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n804), .A2(G159), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n378), .B1(new_n800), .B2(G50), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1243), .A2(new_n1189), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G132), .A2(new_n794), .B1(new_n793), .B2(G150), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n852), .B2(new_n1034), .C1(new_n848), .C2(new_n1142), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G283), .A2(new_n788), .B1(new_n794), .B2(G294), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n215), .B2(new_n847), .C1(new_n469), .C2(new_n848), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1052), .B(new_n342), .C1(new_n213), .C2(new_n797), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G97), .B2(new_n804), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n496), .B2(new_n783), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n1246), .A2(new_n1248), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1242), .B1(new_n1254), .B2(new_n776), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT125), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1111), .B2(new_n823), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1119), .B2(new_n770), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1241), .A2(new_n1258), .ZN(G381));
  OR2_X1    g1059(.A1(G390), .A2(G384), .ZN(new_n1260));
  OR2_X1    g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(new_n1260), .A2(G387), .A3(G381), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(G378), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1211), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1229), .A2(new_n1182), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1230), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n712), .B1(new_n1229), .B2(new_n1235), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1264), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1262), .A2(new_n1263), .A3(new_n1268), .ZN(G407));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1263), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G407), .B(G213), .C1(G343), .C2(new_n1270), .ZN(G409));
  AOI211_X1 g1071(.A(new_n1001), .B(new_n1181), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1178), .A2(new_n930), .A3(new_n1179), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1233), .B1(new_n1232), .B2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1180), .A2(KEYINPUT124), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n770), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1183), .A2(new_n1210), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1276), .A2(new_n1139), .A3(new_n1163), .A4(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(G213), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n1272), .A2(new_n1278), .B1(new_n1279), .B2(G343), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1268), .B2(new_n1263), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n839), .A2(KEYINPUT126), .A3(new_n866), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1258), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1213), .A2(KEYINPUT60), .A3(new_n1225), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1285), .A2(new_n711), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT60), .B1(new_n1213), .B2(new_n1225), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1240), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1284), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT126), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G384), .A2(new_n1290), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1279), .A2(G343), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(G2897), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1292), .A2(G2897), .A3(new_n1295), .A4(new_n1293), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1299), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1281), .B(new_n1294), .C1(new_n1268), .C2(new_n1263), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT63), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  XOR2_X1   g1103(.A(G393), .B(G396), .Z(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1010), .A2(new_n1038), .A3(G390), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G390), .B1(new_n1010), .B2(new_n1038), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1305), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(G390), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G387), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1010), .A2(new_n1038), .A3(G390), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n1304), .A3(new_n1311), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1308), .A2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1280), .B1(G375), .B2(G378), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(KEYINPUT63), .A3(new_n1294), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1300), .A2(new_n1303), .A3(new_n1313), .A4(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1314), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1301), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1314), .A2(KEYINPUT62), .A3(new_n1294), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1319), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1308), .A2(new_n1312), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT127), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1308), .A2(new_n1312), .A3(KEYINPUT127), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1316), .B1(new_n1323), .B2(new_n1328), .ZN(G405));
  NAND2_X1  g1129(.A1(G375), .A2(G378), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1270), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1294), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1330), .A2(new_n1270), .A3(new_n1294), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1324), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1333), .A2(new_n1313), .A3(new_n1334), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(G402));
endmodule


