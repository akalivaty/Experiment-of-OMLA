

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U548 ( .A1(n667), .A2(n653), .ZN(n661) );
  XNOR2_X1 U549 ( .A(n638), .B(KEYINPUT95), .ZN(n518) );
  AND2_X1 U550 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U551 ( .A(n519), .B(KEYINPUT29), .ZN(n687) );
  INV_X1 U552 ( .A(n735), .ZN(n527) );
  XNOR2_X1 U553 ( .A(n522), .B(n521), .ZN(n520) );
  INV_X1 U554 ( .A(KEYINPUT28), .ZN(n521) );
  NOR2_X1 U555 ( .A1(n680), .A2(n811), .ZN(n522) );
  INV_X1 U556 ( .A(KEYINPUT100), .ZN(n698) );
  OR2_X2 U557 ( .A1(n773), .A2(n625), .ZN(n638) );
  NAND2_X1 U558 ( .A1(n525), .A2(n526), .ZN(n729) );
  NOR2_X1 U559 ( .A1(n514), .A2(n512), .ZN(n526) );
  XOR2_X1 U560 ( .A(KEYINPUT15), .B(n660), .Z(n962) );
  NOR2_X1 U561 ( .A1(G651), .A2(n579), .ZN(n795) );
  AND2_X1 U562 ( .A1(n523), .A2(n513), .ZN(n511) );
  NOR2_X1 U563 ( .A1(n527), .A2(KEYINPUT33), .ZN(n512) );
  INV_X1 U564 ( .A(G2105), .ZN(n550) );
  XNOR2_X1 U565 ( .A(KEYINPUT104), .B(n752), .ZN(n513) );
  NAND2_X1 U566 ( .A1(n727), .A2(n934), .ZN(n514) );
  AND2_X1 U567 ( .A1(n751), .A2(n940), .ZN(n515) );
  NOR2_X1 U568 ( .A1(n740), .A2(n515), .ZN(n516) );
  XNOR2_X2 U569 ( .A(n517), .B(KEYINPUT64), .ZN(n700) );
  NAND2_X1 U570 ( .A1(n518), .A2(n639), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n681), .A2(n520), .ZN(n519) );
  NAND2_X1 U572 ( .A1(n524), .A2(n516), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n739), .A2(n529), .ZN(n524) );
  NAND2_X1 U574 ( .A1(n723), .A2(n724), .ZN(n525) );
  XNOR2_X1 U575 ( .A(n620), .B(KEYINPUT66), .ZN(n773) );
  XOR2_X1 U576 ( .A(n710), .B(KEYINPUT96), .Z(n528) );
  AND2_X1 U577 ( .A1(n738), .A2(n737), .ZN(n529) );
  INV_X1 U578 ( .A(KEYINPUT103), .ZN(n728) );
  NOR2_X1 U579 ( .A1(n579), .A2(n535), .ZN(n793) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n800) );
  XNOR2_X1 U581 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n753) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n579) );
  INV_X1 U583 ( .A(G651), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n793), .A2(G76), .ZN(n530) );
  XNOR2_X1 U585 ( .A(KEYINPUT76), .B(n530), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n800), .A2(G89), .ZN(n531) );
  XNOR2_X1 U587 ( .A(KEYINPUT4), .B(n531), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U589 ( .A(KEYINPUT5), .B(n534), .ZN(n544) );
  XNOR2_X1 U590 ( .A(KEYINPUT6), .B(KEYINPUT78), .ZN(n542) );
  NOR2_X1 U591 ( .A1(G543), .A2(n535), .ZN(n537) );
  XNOR2_X1 U592 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n536) );
  XNOR2_X1 U593 ( .A(n537), .B(n536), .ZN(n799) );
  NAND2_X1 U594 ( .A1(n799), .A2(G63), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n795), .A2(G51), .ZN(n538) );
  XOR2_X1 U596 ( .A(KEYINPUT77), .B(n538), .Z(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U598 ( .A(n542), .B(n541), .Z(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U600 ( .A(KEYINPUT7), .B(n545), .ZN(G168) );
  XOR2_X1 U601 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U602 ( .A1(G2105), .A2(G2104), .ZN(n546) );
  XOR2_X1 U603 ( .A(KEYINPUT17), .B(n546), .Z(n621) );
  NAND2_X1 U604 ( .A1(G138), .A2(n621), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n550), .A2(G2104), .ZN(n547) );
  XNOR2_X2 U606 ( .A(n547), .B(KEYINPUT65), .ZN(n614) );
  NAND2_X1 U607 ( .A1(G102), .A2(n614), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n554) );
  NOR2_X1 U609 ( .A1(G2104), .A2(n550), .ZN(n617) );
  NAND2_X1 U610 ( .A1(G126), .A2(n617), .ZN(n552) );
  AND2_X1 U611 ( .A1(G2105), .A2(G2104), .ZN(n990) );
  NAND2_X1 U612 ( .A1(G114), .A2(n990), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U614 ( .A1(n554), .A2(n553), .ZN(G164) );
  NAND2_X1 U615 ( .A1(G65), .A2(n799), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G78), .A2(n793), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n559) );
  NAND2_X1 U618 ( .A1(G91), .A2(n800), .ZN(n557) );
  XNOR2_X1 U619 ( .A(KEYINPUT71), .B(n557), .ZN(n558) );
  NOR2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n795), .A2(G53), .ZN(n560) );
  NAND2_X1 U622 ( .A1(n561), .A2(n560), .ZN(G299) );
  NAND2_X1 U623 ( .A1(n795), .A2(G52), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n799), .A2(G64), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G90), .A2(n800), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G77), .A2(n793), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT9), .B(n566), .Z(n567) );
  XNOR2_X1 U630 ( .A(KEYINPUT70), .B(n567), .ZN(n568) );
  NOR2_X1 U631 ( .A1(n569), .A2(n568), .ZN(G171) );
  INV_X1 U632 ( .A(G171), .ZN(G301) );
  NAND2_X1 U633 ( .A1(G88), .A2(n800), .ZN(n571) );
  NAND2_X1 U634 ( .A1(G75), .A2(n793), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G62), .A2(n799), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G50), .A2(n795), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U639 ( .A1(n575), .A2(n574), .ZN(G166) );
  INV_X1 U640 ( .A(G166), .ZN(G303) );
  NAND2_X1 U641 ( .A1(G49), .A2(n795), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G74), .A2(G651), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U644 ( .A1(n799), .A2(n578), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n579), .A2(G87), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(G288) );
  NAND2_X1 U647 ( .A1(G61), .A2(n799), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G86), .A2(n800), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n793), .A2(G73), .ZN(n584) );
  XOR2_X1 U651 ( .A(KEYINPUT2), .B(n584), .Z(n585) );
  NOR2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n795), .A2(G48), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(G305) );
  NAND2_X1 U655 ( .A1(G72), .A2(n793), .ZN(n589) );
  XNOR2_X1 U656 ( .A(n589), .B(KEYINPUT68), .ZN(n596) );
  NAND2_X1 U657 ( .A1(G60), .A2(n799), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G47), .A2(n795), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U660 ( .A1(G85), .A2(n800), .ZN(n592) );
  XNOR2_X1 U661 ( .A(KEYINPUT67), .B(n592), .ZN(n593) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n595), .ZN(G290) );
  BUF_X1 U664 ( .A(n621), .Z(n993) );
  NAND2_X1 U665 ( .A1(G131), .A2(n993), .ZN(n598) );
  NAND2_X1 U666 ( .A1(G107), .A2(n990), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n598), .A2(n597), .ZN(n601) );
  BUF_X1 U668 ( .A(n617), .Z(n989) );
  NAND2_X1 U669 ( .A1(n989), .A2(G119), .ZN(n599) );
  XOR2_X1 U670 ( .A(KEYINPUT92), .B(n599), .Z(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n614), .A2(G95), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n1006) );
  NAND2_X1 U674 ( .A1(G1991), .A2(n1006), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n604), .B(KEYINPUT93), .ZN(n613) );
  NAND2_X1 U676 ( .A1(G129), .A2(n989), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G117), .A2(n990), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n614), .A2(G105), .ZN(n607) );
  XOR2_X1 U680 ( .A(KEYINPUT38), .B(n607), .Z(n608) );
  NOR2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n993), .A2(G141), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n1003) );
  AND2_X1 U684 ( .A1(G1996), .A2(n1003), .ZN(n612) );
  NOR2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n854) );
  NOR2_X1 U686 ( .A1(G164), .A2(G1384), .ZN(n639) );
  NAND2_X1 U687 ( .A1(n614), .A2(G101), .ZN(n616) );
  INV_X1 U688 ( .A(KEYINPUT23), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n616), .B(n615), .ZN(n619) );
  NAND2_X1 U690 ( .A1(n617), .A2(G125), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U692 ( .A1(G137), .A2(n621), .ZN(n623) );
  NAND2_X1 U693 ( .A1(G113), .A2(n990), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n774) );
  INV_X1 U695 ( .A(G40), .ZN(n624) );
  OR2_X1 U696 ( .A1(n774), .A2(n624), .ZN(n625) );
  NOR2_X1 U697 ( .A1(n639), .A2(n638), .ZN(n751) );
  INV_X1 U698 ( .A(n751), .ZN(n626) );
  NOR2_X1 U699 ( .A1(n854), .A2(n626), .ZN(n743) );
  INV_X1 U700 ( .A(n743), .ZN(n636) );
  NAND2_X1 U701 ( .A1(G140), .A2(n993), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G104), .A2(n614), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U704 ( .A(KEYINPUT34), .B(n629), .ZN(n634) );
  NAND2_X1 U705 ( .A1(G128), .A2(n989), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G116), .A2(n990), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U708 ( .A(KEYINPUT35), .B(n632), .Z(n633) );
  NOR2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U710 ( .A(KEYINPUT36), .B(n635), .ZN(n1013) );
  XNOR2_X1 U711 ( .A(G2067), .B(KEYINPUT37), .ZN(n748) );
  NOR2_X1 U712 ( .A1(n1013), .A2(n748), .ZN(n857) );
  NAND2_X1 U713 ( .A1(n751), .A2(n857), .ZN(n746) );
  NAND2_X1 U714 ( .A1(n636), .A2(n746), .ZN(n637) );
  XNOR2_X1 U715 ( .A(KEYINPUT94), .B(n637), .ZN(n740) );
  INV_X1 U716 ( .A(KEYINPUT33), .ZN(n724) );
  NAND2_X1 U717 ( .A1(n700), .A2(G8), .ZN(n735) );
  INV_X1 U718 ( .A(G1996), .ZN(n640) );
  NOR2_X1 U719 ( .A1(n700), .A2(n640), .ZN(n642) );
  INV_X1 U720 ( .A(KEYINPUT26), .ZN(n641) );
  XNOR2_X1 U721 ( .A(n642), .B(n641), .ZN(n667) );
  NAND2_X1 U722 ( .A1(n700), .A2(G1341), .ZN(n665) );
  NAND2_X1 U723 ( .A1(n800), .A2(G81), .ZN(n643) );
  XNOR2_X1 U724 ( .A(n643), .B(KEYINPUT12), .ZN(n645) );
  NAND2_X1 U725 ( .A1(G68), .A2(n793), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U727 ( .A(KEYINPUT13), .B(n646), .ZN(n652) );
  NAND2_X1 U728 ( .A1(G56), .A2(n799), .ZN(n647) );
  XOR2_X1 U729 ( .A(KEYINPUT14), .B(n647), .Z(n650) );
  NAND2_X1 U730 ( .A1(G43), .A2(n795), .ZN(n648) );
  XNOR2_X1 U731 ( .A(KEYINPUT75), .B(n648), .ZN(n649) );
  NOR2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n943) );
  INV_X1 U734 ( .A(n943), .ZN(n663) );
  AND2_X1 U735 ( .A1(n665), .A2(n663), .ZN(n653) );
  NAND2_X1 U736 ( .A1(G92), .A2(n800), .ZN(n655) );
  NAND2_X1 U737 ( .A1(G79), .A2(n793), .ZN(n654) );
  NAND2_X1 U738 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U739 ( .A1(G66), .A2(n799), .ZN(n657) );
  NAND2_X1 U740 ( .A1(G54), .A2(n795), .ZN(n656) );
  NAND2_X1 U741 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U742 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U743 ( .A1(n661), .A2(n962), .ZN(n662) );
  XNOR2_X1 U744 ( .A(n662), .B(KEYINPUT99), .ZN(n674) );
  AND2_X1 U745 ( .A1(n663), .A2(n962), .ZN(n664) );
  AND2_X1 U746 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n668), .B(KEYINPUT98), .ZN(n672) );
  INV_X1 U749 ( .A(n700), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n683), .A2(G1348), .ZN(n670) );
  NOR2_X1 U751 ( .A1(n700), .A2(G2067), .ZN(n669) );
  NOR2_X1 U752 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n674), .A2(n673), .ZN(n679) );
  INV_X1 U755 ( .A(G299), .ZN(n811) );
  NAND2_X1 U756 ( .A1(G2072), .A2(n683), .ZN(n675) );
  XNOR2_X1 U757 ( .A(n675), .B(KEYINPUT27), .ZN(n677) );
  INV_X1 U758 ( .A(G1956), .ZN(n883) );
  NOR2_X1 U759 ( .A1(n683), .A2(n883), .ZN(n676) );
  NOR2_X1 U760 ( .A1(n677), .A2(n676), .ZN(n680) );
  NAND2_X1 U761 ( .A1(n811), .A2(n680), .ZN(n678) );
  NAND2_X1 U762 ( .A1(n679), .A2(n678), .ZN(n681) );
  XNOR2_X1 U763 ( .A(G2078), .B(KEYINPUT25), .ZN(n917) );
  NAND2_X1 U764 ( .A1(n683), .A2(n917), .ZN(n682) );
  XNOR2_X1 U765 ( .A(n682), .B(KEYINPUT97), .ZN(n685) );
  NOR2_X1 U766 ( .A1(n683), .A2(G1961), .ZN(n684) );
  NOR2_X1 U767 ( .A1(n685), .A2(n684), .ZN(n692) );
  NOR2_X1 U768 ( .A1(G301), .A2(n692), .ZN(n686) );
  NOR2_X1 U769 ( .A1(n687), .A2(n686), .ZN(n697) );
  NOR2_X1 U770 ( .A1(G1966), .A2(n735), .ZN(n711) );
  NOR2_X1 U771 ( .A1(n700), .A2(G2084), .ZN(n709) );
  INV_X1 U772 ( .A(n709), .ZN(n688) );
  NAND2_X1 U773 ( .A1(G8), .A2(n688), .ZN(n689) );
  OR2_X1 U774 ( .A1(n711), .A2(n689), .ZN(n690) );
  XNOR2_X1 U775 ( .A(KEYINPUT30), .B(n690), .ZN(n691) );
  NOR2_X1 U776 ( .A1(n691), .A2(G168), .ZN(n694) );
  AND2_X1 U777 ( .A1(G301), .A2(n692), .ZN(n693) );
  NOR2_X1 U778 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U779 ( .A(n695), .B(KEYINPUT31), .ZN(n696) );
  NOR2_X1 U780 ( .A1(n697), .A2(n696), .ZN(n699) );
  XNOR2_X1 U781 ( .A(n699), .B(n698), .ZN(n713) );
  NAND2_X1 U782 ( .A1(n713), .A2(G286), .ZN(n706) );
  NOR2_X1 U783 ( .A1(n700), .A2(G2090), .ZN(n701) );
  XNOR2_X1 U784 ( .A(n701), .B(KEYINPUT102), .ZN(n703) );
  NOR2_X1 U785 ( .A1(n735), .A2(G1971), .ZN(n702) );
  NOR2_X1 U786 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n704), .A2(G303), .ZN(n705) );
  NAND2_X1 U788 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U789 ( .A1(n707), .A2(G8), .ZN(n708) );
  XNOR2_X1 U790 ( .A(n708), .B(KEYINPUT32), .ZN(n720) );
  NAND2_X1 U791 ( .A1(n709), .A2(G8), .ZN(n710) );
  NOR2_X1 U792 ( .A1(n711), .A2(n528), .ZN(n712) );
  NAND2_X1 U793 ( .A1(KEYINPUT101), .A2(n714), .ZN(n718) );
  INV_X1 U794 ( .A(KEYINPUT101), .ZN(n716) );
  INV_X1 U795 ( .A(n714), .ZN(n715) );
  NAND2_X1 U796 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U797 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U798 ( .A1(n720), .A2(n719), .ZN(n732) );
  NOR2_X1 U799 ( .A1(G1976), .A2(G288), .ZN(n725) );
  NOR2_X1 U800 ( .A1(G1971), .A2(G303), .ZN(n721) );
  NOR2_X1 U801 ( .A1(n725), .A2(n721), .ZN(n950) );
  NAND2_X1 U802 ( .A1(n732), .A2(n950), .ZN(n722) );
  NAND2_X1 U803 ( .A1(G1976), .A2(G288), .ZN(n941) );
  NAND2_X1 U804 ( .A1(n722), .A2(n941), .ZN(n723) );
  NAND2_X1 U805 ( .A1(n725), .A2(KEYINPUT33), .ZN(n726) );
  OR2_X1 U806 ( .A1(n726), .A2(n735), .ZN(n727) );
  XOR2_X1 U807 ( .A(G1981), .B(G305), .Z(n934) );
  XNOR2_X1 U808 ( .A(n729), .B(n728), .ZN(n739) );
  NOR2_X1 U809 ( .A1(G1981), .A2(G305), .ZN(n730) );
  XOR2_X1 U810 ( .A(n730), .B(KEYINPUT24), .Z(n731) );
  OR2_X1 U811 ( .A1(n735), .A2(n731), .ZN(n738) );
  NOR2_X1 U812 ( .A1(G2090), .A2(G303), .ZN(n733) );
  NAND2_X1 U813 ( .A1(G8), .A2(n733), .ZN(n734) );
  NAND2_X1 U814 ( .A1(n732), .A2(n734), .ZN(n736) );
  NAND2_X1 U815 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U816 ( .A(G1986), .B(G290), .ZN(n940) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n1003), .ZN(n869) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n741) );
  NOR2_X1 U819 ( .A1(G1991), .A2(n1006), .ZN(n851) );
  NOR2_X1 U820 ( .A1(n741), .A2(n851), .ZN(n742) );
  NOR2_X1 U821 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U822 ( .A1(n869), .A2(n744), .ZN(n745) );
  XNOR2_X1 U823 ( .A(n745), .B(KEYINPUT39), .ZN(n747) );
  NAND2_X1 U824 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U825 ( .A1(n1013), .A2(n748), .ZN(n855) );
  NAND2_X1 U826 ( .A1(n749), .A2(n855), .ZN(n750) );
  NAND2_X1 U827 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U828 ( .A(n511), .B(n753), .ZN(G329) );
  XOR2_X1 U829 ( .A(G2427), .B(G2438), .Z(n755) );
  XNOR2_X1 U830 ( .A(G1341), .B(G2454), .ZN(n754) );
  XNOR2_X1 U831 ( .A(n755), .B(n754), .ZN(n756) );
  XOR2_X1 U832 ( .A(n756), .B(G2451), .Z(n758) );
  XNOR2_X1 U833 ( .A(G1348), .B(KEYINPUT106), .ZN(n757) );
  XNOR2_X1 U834 ( .A(n758), .B(n757), .ZN(n762) );
  XOR2_X1 U835 ( .A(G2430), .B(G2435), .Z(n760) );
  XNOR2_X1 U836 ( .A(G2446), .B(G2443), .ZN(n759) );
  XNOR2_X1 U837 ( .A(n760), .B(n759), .ZN(n761) );
  XOR2_X1 U838 ( .A(n762), .B(n761), .Z(n763) );
  AND2_X1 U839 ( .A1(G14), .A2(n763), .ZN(G401) );
  AND2_X1 U840 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U841 ( .A1(n989), .A2(G123), .ZN(n764) );
  XNOR2_X1 U842 ( .A(n764), .B(KEYINPUT18), .ZN(n766) );
  NAND2_X1 U843 ( .A1(G111), .A2(n990), .ZN(n765) );
  NAND2_X1 U844 ( .A1(n766), .A2(n765), .ZN(n770) );
  NAND2_X1 U845 ( .A1(G135), .A2(n993), .ZN(n768) );
  NAND2_X1 U846 ( .A1(G99), .A2(n614), .ZN(n767) );
  NAND2_X1 U847 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U848 ( .A1(n770), .A2(n769), .ZN(n1002) );
  XNOR2_X1 U849 ( .A(n1002), .B(G2096), .ZN(n771) );
  XNOR2_X1 U850 ( .A(n771), .B(KEYINPUT83), .ZN(n772) );
  OR2_X1 U851 ( .A1(G2100), .A2(n772), .ZN(G156) );
  INV_X1 U852 ( .A(G82), .ZN(G220) );
  NOR2_X1 U853 ( .A1(n773), .A2(n774), .ZN(G160) );
  NAND2_X1 U854 ( .A1(G7), .A2(G661), .ZN(n775) );
  XNOR2_X1 U855 ( .A(n775), .B(KEYINPUT10), .ZN(n776) );
  XNOR2_X1 U856 ( .A(KEYINPUT74), .B(n776), .ZN(G223) );
  INV_X1 U857 ( .A(G223), .ZN(n837) );
  NAND2_X1 U858 ( .A1(n837), .A2(G567), .ZN(n777) );
  XOR2_X1 U859 ( .A(KEYINPUT11), .B(n777), .Z(G234) );
  INV_X1 U860 ( .A(G860), .ZN(n783) );
  OR2_X1 U861 ( .A1(n943), .A2(n783), .ZN(G153) );
  NAND2_X1 U862 ( .A1(G868), .A2(G301), .ZN(n779) );
  OR2_X1 U863 ( .A1(n962), .A2(G868), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n779), .A2(n778), .ZN(G284) );
  INV_X1 U865 ( .A(G868), .ZN(n817) );
  NOR2_X1 U866 ( .A1(G286), .A2(n817), .ZN(n781) );
  NOR2_X1 U867 ( .A1(G868), .A2(G299), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U869 ( .A(KEYINPUT79), .B(n782), .Z(G297) );
  NAND2_X1 U870 ( .A1(G559), .A2(n783), .ZN(n784) );
  XNOR2_X1 U871 ( .A(KEYINPUT80), .B(n784), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n785), .A2(n962), .ZN(n787) );
  XOR2_X1 U873 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n786) );
  XNOR2_X1 U874 ( .A(n787), .B(n786), .ZN(G148) );
  NAND2_X1 U875 ( .A1(n962), .A2(G868), .ZN(n788) );
  NOR2_X1 U876 ( .A1(G559), .A2(n788), .ZN(n789) );
  XNOR2_X1 U877 ( .A(n789), .B(KEYINPUT82), .ZN(n791) );
  NOR2_X1 U878 ( .A1(n943), .A2(G868), .ZN(n790) );
  NOR2_X1 U879 ( .A1(n791), .A2(n790), .ZN(G282) );
  NAND2_X1 U880 ( .A1(n962), .A2(G559), .ZN(n814) );
  XNOR2_X1 U881 ( .A(n943), .B(n814), .ZN(n792) );
  NOR2_X1 U882 ( .A1(n792), .A2(G860), .ZN(n805) );
  NAND2_X1 U883 ( .A1(G80), .A2(n793), .ZN(n794) );
  XNOR2_X1 U884 ( .A(n794), .B(KEYINPUT84), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G55), .A2(n795), .ZN(n796) );
  XOR2_X1 U886 ( .A(KEYINPUT85), .B(n796), .Z(n797) );
  NAND2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n804) );
  NAND2_X1 U888 ( .A1(G67), .A2(n799), .ZN(n802) );
  NAND2_X1 U889 ( .A1(G93), .A2(n800), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n803) );
  OR2_X1 U891 ( .A1(n804), .A2(n803), .ZN(n816) );
  XOR2_X1 U892 ( .A(n805), .B(n816), .Z(G145) );
  XOR2_X1 U893 ( .A(n943), .B(G305), .Z(n806) );
  XNOR2_X1 U894 ( .A(G290), .B(n806), .ZN(n810) );
  XNOR2_X1 U895 ( .A(KEYINPUT86), .B(KEYINPUT19), .ZN(n808) );
  XOR2_X1 U896 ( .A(G288), .B(n816), .Z(n807) );
  XNOR2_X1 U897 ( .A(n808), .B(n807), .ZN(n809) );
  XOR2_X1 U898 ( .A(n810), .B(n809), .Z(n813) );
  XNOR2_X1 U899 ( .A(n811), .B(G166), .ZN(n812) );
  XNOR2_X1 U900 ( .A(n813), .B(n812), .ZN(n961) );
  XNOR2_X1 U901 ( .A(n814), .B(n961), .ZN(n815) );
  NAND2_X1 U902 ( .A1(n815), .A2(G868), .ZN(n819) );
  NAND2_X1 U903 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U904 ( .A1(n819), .A2(n818), .ZN(G295) );
  XOR2_X1 U905 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n823) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n820) );
  XOR2_X1 U907 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U908 ( .A1(n821), .A2(G2090), .ZN(n822) );
  XNOR2_X1 U909 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U910 ( .A1(G2072), .A2(n824), .ZN(G158) );
  XOR2_X1 U911 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U912 ( .A(KEYINPUT88), .B(G44), .ZN(n825) );
  XNOR2_X1 U913 ( .A(n825), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U914 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  NAND2_X1 U915 ( .A1(G120), .A2(G108), .ZN(n826) );
  NOR2_X1 U916 ( .A1(G237), .A2(n826), .ZN(n827) );
  NAND2_X1 U917 ( .A1(G69), .A2(n827), .ZN(n960) );
  NAND2_X1 U918 ( .A1(n960), .A2(G567), .ZN(n834) );
  NOR2_X1 U919 ( .A1(G220), .A2(G219), .ZN(n829) );
  XNOR2_X1 U920 ( .A(KEYINPUT22), .B(KEYINPUT89), .ZN(n828) );
  XNOR2_X1 U921 ( .A(n829), .B(n828), .ZN(n830) );
  NOR2_X1 U922 ( .A1(G218), .A2(n830), .ZN(n831) );
  NAND2_X1 U923 ( .A1(G96), .A2(n831), .ZN(n959) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n959), .ZN(n832) );
  XNOR2_X1 U925 ( .A(KEYINPUT90), .B(n832), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(n1023) );
  NAND2_X1 U927 ( .A1(G661), .A2(G483), .ZN(n835) );
  NOR2_X1 U928 ( .A1(n1023), .A2(n835), .ZN(n840) );
  NAND2_X1 U929 ( .A1(G36), .A2(n840), .ZN(n836) );
  XOR2_X1 U930 ( .A(KEYINPUT91), .B(n836), .Z(G176) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U933 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n839) );
  XOR2_X1 U935 ( .A(KEYINPUT107), .B(n839), .Z(n841) );
  NAND2_X1 U936 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n842), .B(KEYINPUT108), .ZN(G188) );
  XNOR2_X1 U938 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  NAND2_X1 U940 ( .A1(G124), .A2(n989), .ZN(n843) );
  XOR2_X1 U941 ( .A(KEYINPUT44), .B(n843), .Z(n844) );
  XNOR2_X1 U942 ( .A(n844), .B(KEYINPUT115), .ZN(n846) );
  NAND2_X1 U943 ( .A1(G112), .A2(n990), .ZN(n845) );
  NAND2_X1 U944 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U945 ( .A1(G136), .A2(n993), .ZN(n848) );
  NAND2_X1 U946 ( .A1(G100), .A2(n614), .ZN(n847) );
  NAND2_X1 U947 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U948 ( .A1(n850), .A2(n849), .ZN(G162) );
  NOR2_X1 U949 ( .A1(n851), .A2(n1002), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n852), .B(KEYINPUT120), .ZN(n853) );
  NAND2_X1 U951 ( .A1(n854), .A2(n853), .ZN(n878) );
  INV_X1 U952 ( .A(n855), .ZN(n856) );
  NOR2_X1 U953 ( .A1(n857), .A2(n856), .ZN(n876) );
  NAND2_X1 U954 ( .A1(G139), .A2(n993), .ZN(n859) );
  NAND2_X1 U955 ( .A1(G103), .A2(n614), .ZN(n858) );
  NAND2_X1 U956 ( .A1(n859), .A2(n858), .ZN(n864) );
  NAND2_X1 U957 ( .A1(G127), .A2(n989), .ZN(n861) );
  NAND2_X1 U958 ( .A1(G115), .A2(n990), .ZN(n860) );
  NAND2_X1 U959 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U960 ( .A(KEYINPUT47), .B(n862), .Z(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n1000) );
  XOR2_X1 U962 ( .A(G2072), .B(n1000), .Z(n866) );
  XOR2_X1 U963 ( .A(G164), .B(G2078), .Z(n865) );
  NOR2_X1 U964 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U965 ( .A(KEYINPUT50), .B(n867), .ZN(n872) );
  XOR2_X1 U966 ( .A(G2090), .B(G162), .Z(n868) );
  NOR2_X1 U967 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U968 ( .A(KEYINPUT51), .B(n870), .Z(n871) );
  NAND2_X1 U969 ( .A1(n872), .A2(n871), .ZN(n874) );
  XOR2_X1 U970 ( .A(G160), .B(G2084), .Z(n873) );
  NOR2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n875) );
  NAND2_X1 U972 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U973 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U974 ( .A(KEYINPUT52), .B(n879), .Z(n880) );
  NOR2_X1 U975 ( .A1(KEYINPUT55), .A2(n880), .ZN(n881) );
  XNOR2_X1 U976 ( .A(KEYINPUT121), .B(n881), .ZN(n882) );
  NAND2_X1 U977 ( .A1(n882), .A2(G29), .ZN(n933) );
  XNOR2_X1 U978 ( .A(G20), .B(n883), .ZN(n887) );
  XNOR2_X1 U979 ( .A(G1341), .B(G19), .ZN(n885) );
  XNOR2_X1 U980 ( .A(G6), .B(G1981), .ZN(n884) );
  NOR2_X1 U981 ( .A1(n885), .A2(n884), .ZN(n886) );
  NAND2_X1 U982 ( .A1(n887), .A2(n886), .ZN(n890) );
  XOR2_X1 U983 ( .A(KEYINPUT59), .B(G1348), .Z(n888) );
  XNOR2_X1 U984 ( .A(G4), .B(n888), .ZN(n889) );
  NOR2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U986 ( .A(KEYINPUT60), .B(n891), .ZN(n895) );
  XNOR2_X1 U987 ( .A(G1966), .B(G21), .ZN(n893) );
  XNOR2_X1 U988 ( .A(G1961), .B(G5), .ZN(n892) );
  NOR2_X1 U989 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U990 ( .A1(n895), .A2(n894), .ZN(n902) );
  XNOR2_X1 U991 ( .A(G1971), .B(G22), .ZN(n897) );
  XNOR2_X1 U992 ( .A(G24), .B(G1986), .ZN(n896) );
  NOR2_X1 U993 ( .A1(n897), .A2(n896), .ZN(n899) );
  XOR2_X1 U994 ( .A(G1976), .B(G23), .Z(n898) );
  NAND2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U996 ( .A(KEYINPUT58), .B(n900), .ZN(n901) );
  NOR2_X1 U997 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U998 ( .A(KEYINPUT61), .B(n903), .ZN(n905) );
  INV_X1 U999 ( .A(G16), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(n906) );
  NAND2_X1 U1001 ( .A1(n906), .A2(G11), .ZN(n931) );
  XNOR2_X1 U1002 ( .A(KEYINPUT126), .B(G2084), .ZN(n909) );
  XNOR2_X1 U1003 ( .A(KEYINPUT54), .B(G34), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n907), .B(KEYINPUT125), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n927) );
  XNOR2_X1 U1006 ( .A(G2090), .B(G35), .ZN(n925) );
  XNOR2_X1 U1007 ( .A(KEYINPUT123), .B(G2067), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n910), .B(G26), .ZN(n916) );
  XOR2_X1 U1009 ( .A(G2072), .B(G33), .Z(n911) );
  NAND2_X1 U1010 ( .A1(G28), .A2(n911), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(G25), .B(G1991), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT122), .B(n912), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n922) );
  XOR2_X1 U1015 ( .A(n917), .B(G27), .Z(n919) );
  XNOR2_X1 U1016 ( .A(G32), .B(G1996), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1018 ( .A(KEYINPUT124), .B(n920), .Z(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(KEYINPUT53), .B(n923), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(KEYINPUT55), .B(n928), .ZN(n929) );
  NOR2_X1 U1024 ( .A1(G29), .A2(n929), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n957) );
  XOR2_X1 U1027 ( .A(G16), .B(KEYINPUT56), .Z(n955) );
  XNOR2_X1 U1028 ( .A(G1966), .B(G168), .ZN(n935) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(n936), .B(KEYINPUT57), .ZN(n947) );
  XNOR2_X1 U1031 ( .A(G1348), .B(n962), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(G1971), .A2(G303), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(G1341), .B(n943), .ZN(n944) );
  NOR2_X1 U1037 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n953) );
  XNOR2_X1 U1039 ( .A(G301), .B(G1961), .ZN(n949) );
  XNOR2_X1 U1040 ( .A(G299), .B(G1956), .ZN(n948) );
  NOR2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1043 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1044 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1045 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1046 ( .A(n958), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1047 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1048 ( .A(G120), .ZN(G236) );
  INV_X1 U1049 ( .A(G96), .ZN(G221) );
  INV_X1 U1050 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(G325) );
  INV_X1 U1052 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1053 ( .A(n961), .B(G286), .Z(n964) );
  XNOR2_X1 U1054 ( .A(G171), .B(n962), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(n964), .B(n963), .ZN(n965) );
  NOR2_X1 U1056 ( .A1(G37), .A2(n965), .ZN(G397) );
  XNOR2_X1 U1057 ( .A(G2078), .B(G2072), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(n966), .B(G2100), .ZN(n976) );
  XOR2_X1 U1059 ( .A(KEYINPUT42), .B(KEYINPUT109), .Z(n968) );
  XNOR2_X1 U1060 ( .A(G2678), .B(KEYINPUT111), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(n968), .B(n967), .ZN(n972) );
  XOR2_X1 U1062 ( .A(KEYINPUT43), .B(G2096), .Z(n970) );
  XNOR2_X1 U1063 ( .A(G2090), .B(KEYINPUT110), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n970), .B(n969), .ZN(n971) );
  XOR2_X1 U1065 ( .A(n972), .B(n971), .Z(n974) );
  XNOR2_X1 U1066 ( .A(G2067), .B(G2084), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n974), .B(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(G227) );
  XOR2_X1 U1069 ( .A(KEYINPUT41), .B(KEYINPUT114), .Z(n978) );
  XNOR2_X1 U1070 ( .A(G1976), .B(G1991), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(n978), .B(n977), .ZN(n988) );
  XOR2_X1 U1072 ( .A(KEYINPUT112), .B(G2474), .Z(n980) );
  XNOR2_X1 U1073 ( .A(G1961), .B(G1971), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(n980), .B(n979), .ZN(n984) );
  XOR2_X1 U1075 ( .A(G1986), .B(G1981), .Z(n982) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G1956), .ZN(n981) );
  XNOR2_X1 U1077 ( .A(n982), .B(n981), .ZN(n983) );
  XOR2_X1 U1078 ( .A(n984), .B(n983), .Z(n986) );
  XNOR2_X1 U1079 ( .A(G1996), .B(KEYINPUT113), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(n986), .B(n985), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(n988), .B(n987), .ZN(G229) );
  NAND2_X1 U1082 ( .A1(G130), .A2(n989), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(G118), .A2(n990), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n999) );
  NAND2_X1 U1085 ( .A1(G142), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(G106), .A2(n614), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1088 ( .A(KEYINPUT116), .B(n996), .Z(n997) );
  XNOR2_X1 U1089 ( .A(KEYINPUT45), .B(n997), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XOR2_X1 U1091 ( .A(n1001), .B(n1000), .Z(n1005) );
  XOR2_X1 U1092 ( .A(n1003), .B(n1002), .Z(n1004) );
  XNOR2_X1 U1093 ( .A(n1005), .B(n1004), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(n1006), .B(G162), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1008), .B(n1007), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(n1010), .B(n1009), .Z(n1012) );
  XNOR2_X1 U1098 ( .A(G164), .B(G160), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1012), .B(n1011), .ZN(n1014) );
  XOR2_X1 U1100 ( .A(n1014), .B(n1013), .Z(n1015) );
  NOR2_X1 U1101 ( .A1(G37), .A2(n1015), .ZN(G395) );
  NOR2_X1 U1102 ( .A1(G401), .A2(n1023), .ZN(n1020) );
  NOR2_X1 U1103 ( .A1(G227), .A2(G229), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(KEYINPUT49), .B(n1016), .Z(n1017) );
  XNOR2_X1 U1105 ( .A(n1017), .B(KEYINPUT117), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(G397), .A2(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(G395), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(n1022), .B(KEYINPUT118), .ZN(G308) );
  INV_X1 U1110 ( .A(G308), .ZN(G225) );
  INV_X1 U1111 ( .A(n1023), .ZN(G319) );
endmodule

