

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593;

  XNOR2_X1 U323 ( .A(n411), .B(n410), .ZN(n536) );
  XOR2_X1 U324 ( .A(G134GAT), .B(G106GAT), .Z(n291) );
  XNOR2_X1 U325 ( .A(n382), .B(n291), .ZN(n341) );
  XNOR2_X1 U326 ( .A(KEYINPUT108), .B(KEYINPUT48), .ZN(n410) );
  XNOR2_X1 U327 ( .A(n342), .B(n341), .ZN(n344) );
  XNOR2_X1 U328 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U329 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U330 ( .A(n351), .B(n350), .Z(n564) );
  XNOR2_X1 U331 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U332 ( .A(n462), .B(n461), .ZN(G1351GAT) );
  XNOR2_X1 U333 ( .A(KEYINPUT81), .B(KEYINPUT17), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n292), .B(KEYINPUT19), .ZN(n293) );
  XOR2_X1 U335 ( .A(n293), .B(KEYINPUT80), .Z(n295) );
  XNOR2_X1 U336 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n325) );
  XOR2_X1 U338 ( .A(G127GAT), .B(G134GAT), .Z(n297) );
  XNOR2_X1 U339 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U341 ( .A(G113GAT), .B(n298), .Z(n426) );
  XNOR2_X1 U342 ( .A(n325), .B(n426), .ZN(n311) );
  XOR2_X1 U343 ( .A(G71GAT), .B(G190GAT), .Z(n300) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(G99GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U346 ( .A(KEYINPUT20), .B(G176GAT), .Z(n302) );
  XNOR2_X1 U347 ( .A(G15GAT), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U349 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U350 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n306) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U353 ( .A(KEYINPUT65), .B(n307), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n514) );
  XOR2_X1 U356 ( .A(G8GAT), .B(G183GAT), .Z(n364) );
  XOR2_X1 U357 ( .A(G36GAT), .B(G190GAT), .Z(n336) );
  XOR2_X1 U358 ( .A(n364), .B(n336), .Z(n313) );
  NAND2_X1 U359 ( .A1(G226GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U361 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n315) );
  XNOR2_X1 U362 ( .A(G64GAT), .B(G92GAT), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U364 ( .A(n317), .B(n316), .Z(n324) );
  XOR2_X1 U365 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n319) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(G211GAT), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n321) );
  XOR2_X1 U368 ( .A(G218GAT), .B(KEYINPUT84), .Z(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n448) );
  INV_X1 U370 ( .A(n448), .ZN(n322) );
  XOR2_X1 U371 ( .A(G176GAT), .B(G204GAT), .Z(n380) );
  XNOR2_X1 U372 ( .A(n322), .B(n380), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n327) );
  INV_X1 U374 ( .A(n325), .ZN(n326) );
  XOR2_X1 U375 ( .A(n327), .B(n326), .Z(n511) );
  INV_X1 U376 ( .A(n511), .ZN(n526) );
  INV_X1 U377 ( .A(KEYINPUT36), .ZN(n352) );
  XOR2_X1 U378 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n329) );
  XNOR2_X1 U379 ( .A(KEYINPUT66), .B(KEYINPUT11), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n351) );
  INV_X1 U381 ( .A(G43GAT), .ZN(n330) );
  NAND2_X1 U382 ( .A1(n330), .A2(G29GAT), .ZN(n333) );
  INV_X1 U383 ( .A(G29GAT), .ZN(n331) );
  NAND2_X1 U384 ( .A1(n331), .A2(G43GAT), .ZN(n332) );
  NAND2_X1 U385 ( .A1(n333), .A2(n332), .ZN(n335) );
  XNOR2_X1 U386 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n391) );
  XOR2_X1 U388 ( .A(n391), .B(n336), .Z(n338) );
  NAND2_X1 U389 ( .A1(G232GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U391 ( .A(G85GAT), .B(G92GAT), .Z(n340) );
  XNOR2_X1 U392 ( .A(G99GAT), .B(KEYINPUT72), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n382) );
  INV_X1 U394 ( .A(KEYINPUT75), .ZN(n343) );
  NAND2_X1 U395 ( .A1(n344), .A2(n343), .ZN(n347) );
  INV_X1 U396 ( .A(n344), .ZN(n345) );
  NAND2_X1 U397 ( .A1(n345), .A2(KEYINPUT75), .ZN(n346) );
  NAND2_X1 U398 ( .A1(n347), .A2(n346), .ZN(n349) );
  XOR2_X1 U399 ( .A(G50GAT), .B(G162GAT), .Z(n438) );
  XNOR2_X1 U400 ( .A(G218GAT), .B(n438), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n352), .B(n564), .ZN(n590) );
  XOR2_X1 U403 ( .A(G57GAT), .B(KEYINPUT69), .Z(n354) );
  XNOR2_X1 U404 ( .A(KEYINPUT70), .B(KEYINPUT13), .ZN(n353) );
  XOR2_X1 U405 ( .A(n354), .B(n353), .Z(n355) );
  XNOR2_X1 U406 ( .A(n355), .B(G64GAT), .ZN(n357) );
  XNOR2_X1 U407 ( .A(G71GAT), .B(G78GAT), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n377) );
  XOR2_X1 U409 ( .A(G22GAT), .B(G155GAT), .Z(n436) );
  XOR2_X1 U410 ( .A(n436), .B(KEYINPUT12), .Z(n359) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U413 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n361) );
  XNOR2_X1 U414 ( .A(KEYINPUT14), .B(KEYINPUT76), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U416 ( .A(n363), .B(n362), .Z(n368) );
  XOR2_X1 U417 ( .A(G15GAT), .B(G1GAT), .Z(n394) );
  XNOR2_X1 U418 ( .A(G127GAT), .B(G211GAT), .ZN(n365) );
  XNOR2_X1 U419 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n394), .B(n366), .ZN(n367) );
  XNOR2_X1 U421 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U422 ( .A(n377), .B(n369), .ZN(n479) );
  NOR2_X1 U423 ( .A1(n590), .A2(n479), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n370), .B(KEYINPUT45), .ZN(n401) );
  XOR2_X1 U425 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n372) );
  NAND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U428 ( .A(n373), .B(KEYINPUT31), .Z(n379) );
  XOR2_X1 U429 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n375) );
  XNOR2_X1 U430 ( .A(G120GAT), .B(KEYINPUT73), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n384) );
  XOR2_X1 U435 ( .A(G106GAT), .B(G148GAT), .Z(n442) );
  XOR2_X1 U436 ( .A(n442), .B(n382), .Z(n383) );
  XNOR2_X1 U437 ( .A(n384), .B(n383), .ZN(n403) );
  XOR2_X1 U438 ( .A(G22GAT), .B(G141GAT), .Z(n386) );
  XNOR2_X1 U439 ( .A(G169GAT), .B(G197GAT), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U441 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n388) );
  XNOR2_X1 U442 ( .A(G113GAT), .B(G8GAT), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n399) );
  XOR2_X1 U445 ( .A(n391), .B(KEYINPUT29), .Z(n393) );
  NAND2_X1 U446 ( .A1(G229GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n395) );
  XOR2_X1 U448 ( .A(n395), .B(n394), .Z(n397) );
  XNOR2_X1 U449 ( .A(G36GAT), .B(G50GAT), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n399), .B(n398), .ZN(n576) );
  INV_X1 U452 ( .A(n576), .ZN(n568) );
  NOR2_X1 U453 ( .A1(n403), .A2(n568), .ZN(n400) );
  NAND2_X1 U454 ( .A1(n401), .A2(n400), .ZN(n409) );
  XOR2_X1 U455 ( .A(KEYINPUT64), .B(KEYINPUT41), .Z(n402) );
  XNOR2_X1 U456 ( .A(n403), .B(n402), .ZN(n558) );
  NAND2_X1 U457 ( .A1(n568), .A2(n558), .ZN(n404) );
  XNOR2_X1 U458 ( .A(KEYINPUT46), .B(n404), .ZN(n405) );
  INV_X1 U459 ( .A(n479), .ZN(n585) );
  XNOR2_X1 U460 ( .A(n585), .B(KEYINPUT107), .ZN(n572) );
  NAND2_X1 U461 ( .A1(n405), .A2(n572), .ZN(n406) );
  NOR2_X1 U462 ( .A1(n564), .A2(n406), .ZN(n407) );
  XNOR2_X1 U463 ( .A(KEYINPUT47), .B(n407), .ZN(n408) );
  NAND2_X1 U464 ( .A1(n409), .A2(n408), .ZN(n411) );
  NAND2_X1 U465 ( .A1(n526), .A2(n536), .ZN(n413) );
  XOR2_X1 U466 ( .A(KEYINPUT54), .B(KEYINPUT117), .Z(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n431) );
  XOR2_X1 U468 ( .A(KEYINPUT88), .B(KEYINPUT5), .Z(n415) );
  XNOR2_X1 U469 ( .A(KEYINPUT4), .B(KEYINPUT87), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n430) );
  XOR2_X1 U471 ( .A(G85GAT), .B(G148GAT), .Z(n417) );
  XNOR2_X1 U472 ( .A(G29GAT), .B(G162GAT), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U474 ( .A(KEYINPUT1), .B(G57GAT), .Z(n419) );
  XNOR2_X1 U475 ( .A(G1GAT), .B(G155GAT), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U477 ( .A(n421), .B(n420), .Z(n428) );
  XNOR2_X1 U478 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n422), .B(KEYINPUT2), .ZN(n439) );
  XOR2_X1 U480 ( .A(n439), .B(KEYINPUT6), .Z(n424) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n524) );
  NOR2_X1 U486 ( .A1(n431), .A2(n524), .ZN(n575) );
  XOR2_X1 U487 ( .A(KEYINPUT82), .B(KEYINPUT24), .Z(n433) );
  XNOR2_X1 U488 ( .A(KEYINPUT86), .B(KEYINPUT83), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n447) );
  XOR2_X1 U490 ( .A(G78GAT), .B(G204GAT), .Z(n435) );
  XNOR2_X1 U491 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U493 ( .A(n437), .B(n436), .Z(n445) );
  XOR2_X1 U494 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U495 ( .A1(G228GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n473) );
  NAND2_X1 U501 ( .A1(n575), .A2(n473), .ZN(n453) );
  XOR2_X1 U502 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n451) );
  INV_X1 U503 ( .A(KEYINPUT55), .ZN(n450) );
  NOR2_X1 U504 ( .A1(n514), .A2(n454), .ZN(n570) );
  XOR2_X1 U505 ( .A(KEYINPUT99), .B(n558), .Z(n542) );
  NAND2_X1 U506 ( .A1(n570), .A2(n542), .ZN(n458) );
  XOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT56), .Z(n456) );
  XNOR2_X1 U508 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  NAND2_X1 U511 ( .A1(n570), .A2(n564), .ZN(n462) );
  XOR2_X1 U512 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n460) );
  XNOR2_X1 U513 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n459) );
  XOR2_X1 U514 ( .A(KEYINPUT95), .B(KEYINPUT34), .Z(n484) );
  NOR2_X1 U515 ( .A1(n576), .A2(n403), .ZN(n496) );
  INV_X1 U516 ( .A(n514), .ZN(n538) );
  NAND2_X1 U517 ( .A1(n526), .A2(n538), .ZN(n463) );
  NAND2_X1 U518 ( .A1(n473), .A2(n463), .ZN(n464) );
  XNOR2_X1 U519 ( .A(n464), .B(KEYINPUT25), .ZN(n470) );
  NOR2_X1 U520 ( .A1(n538), .A2(n473), .ZN(n466) );
  XNOR2_X1 U521 ( .A(KEYINPUT92), .B(KEYINPUT26), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U523 ( .A(KEYINPUT91), .B(n467), .Z(n574) );
  INV_X1 U524 ( .A(n574), .ZN(n468) );
  XOR2_X1 U525 ( .A(n526), .B(KEYINPUT27), .Z(n475) );
  NOR2_X1 U526 ( .A1(n468), .A2(n475), .ZN(n469) );
  NOR2_X1 U527 ( .A1(n470), .A2(n469), .ZN(n471) );
  NOR2_X1 U528 ( .A1(n471), .A2(n524), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n472), .B(KEYINPUT93), .ZN(n478) );
  XNOR2_X1 U530 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n474), .B(n473), .ZN(n540) );
  NOR2_X1 U532 ( .A1(n538), .A2(n540), .ZN(n476) );
  INV_X1 U533 ( .A(n524), .ZN(n507) );
  NOR2_X1 U534 ( .A1(n507), .A2(n475), .ZN(n535) );
  NAND2_X1 U535 ( .A1(n476), .A2(n535), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n494) );
  OR2_X1 U537 ( .A1(n479), .A2(n564), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n480), .Z(n481) );
  AND2_X1 U539 ( .A1(n494), .A2(n481), .ZN(n506) );
  NAND2_X1 U540 ( .A1(n496), .A2(n506), .ZN(n482) );
  XOR2_X1 U541 ( .A(KEYINPUT94), .B(n482), .Z(n490) );
  NAND2_X1 U542 ( .A1(n490), .A2(n524), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n490), .A2(n526), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(KEYINPUT96), .ZN(n487) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n487), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .Z(n489) );
  NAND2_X1 U549 ( .A1(n490), .A2(n538), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  XOR2_X1 U551 ( .A(G22GAT), .B(KEYINPUT97), .Z(n492) );
  NAND2_X1 U552 ( .A1(n490), .A2(n540), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(G1327GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT39), .B(KEYINPUT98), .Z(n499) );
  NOR2_X1 U555 ( .A1(n590), .A2(n585), .ZN(n493) );
  NAND2_X1 U556 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U557 ( .A(KEYINPUT37), .B(n495), .ZN(n521) );
  NAND2_X1 U558 ( .A1(n521), .A2(n496), .ZN(n497) );
  XOR2_X1 U559 ( .A(KEYINPUT38), .B(n497), .Z(n504) );
  NAND2_X1 U560 ( .A1(n504), .A2(n524), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U563 ( .A1(n504), .A2(n526), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n501), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U565 ( .A1(n504), .A2(n538), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n504), .A2(n540), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(G50GAT), .ZN(G1331GAT) );
  AND2_X1 U570 ( .A1(n542), .A2(n576), .ZN(n522) );
  NAND2_X1 U571 ( .A1(n522), .A2(n506), .ZN(n516) );
  NOR2_X1 U572 ( .A1(n507), .A2(n516), .ZN(n509) );
  XNOR2_X1 U573 ( .A(KEYINPUT100), .B(KEYINPUT42), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n510), .Z(G1332GAT) );
  NOR2_X1 U576 ( .A1(n511), .A2(n516), .ZN(n513) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(KEYINPUT101), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1333GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n516), .ZN(n515) );
  XOR2_X1 U580 ( .A(G71GAT), .B(n515), .Z(G1334GAT) );
  INV_X1 U581 ( .A(n540), .ZN(n517) );
  NOR2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n519) );
  XNOR2_X1 U583 ( .A(KEYINPUT102), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(KEYINPUT103), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n524), .A2(n530), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n530), .A2(n526), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n538), .A2(n530), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(KEYINPUT104), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(KEYINPUT105), .ZN(n534) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT106), .Z(n532) );
  NAND2_X1 U597 ( .A1(n530), .A2(n540), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(G1339GAT) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n537), .B(KEYINPUT109), .ZN(n554) );
  NAND2_X1 U602 ( .A1(n554), .A2(n538), .ZN(n539) );
  NOR2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n568), .A2(n550), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n541), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U607 ( .A1(n550), .A2(n542), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT110), .B(KEYINPUT50), .Z(n546) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(KEYINPUT111), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n549) );
  INV_X1 U612 ( .A(n550), .ZN(n547) );
  NOR2_X1 U613 ( .A1(n572), .A2(n547), .ZN(n548) );
  XOR2_X1 U614 ( .A(n549), .B(n548), .Z(G1342GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U616 ( .A1(n550), .A2(n564), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(n553), .ZN(G1343GAT) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT114), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n574), .A2(n554), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT113), .B(n555), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n565), .A2(n568), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT52), .B(KEYINPUT115), .Z(n560) );
  NAND2_X1 U625 ( .A1(n565), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT53), .Z(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1345GAT) );
  NAND2_X1 U629 ( .A1(n565), .A2(n585), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT116), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n570), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G169GAT), .ZN(G1348GAT) );
  INV_X1 U636 ( .A(n570), .ZN(n571) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G183GAT), .B(n573), .Z(G1350GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n589) );
  NOR2_X1 U640 ( .A1(n576), .A2(n589), .ZN(n581) );
  XOR2_X1 U641 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n578) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(KEYINPUT123), .B(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n583) );
  INV_X1 U647 ( .A(n589), .ZN(n586) );
  NAND2_X1 U648 ( .A1(n586), .A2(n403), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n584), .Z(G1353GAT) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(KEYINPUT126), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G211GAT), .B(n588), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U655 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

