//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055;
  XNOR2_X1  g000(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n194), .B(KEYINPUT1), .C1(new_n191), .C2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n194), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n189), .B2(G143), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n191), .A2(KEYINPUT65), .A3(G146), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n200), .A2(new_n201), .B1(G143), .B2(new_n189), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G137), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(G137), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n209), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n213), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n208), .A2(G137), .ZN(new_n216));
  OAI21_X1  g030(.A(G131), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n206), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G131), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT66), .A3(new_n214), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n222), .A3(G131), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n202), .A2(new_n224), .B1(new_n193), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n221), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n218), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g043(.A(KEYINPUT2), .B(G113), .Z(new_n230));
  XNOR2_X1  g044(.A(G116), .B(G119), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n230), .A2(new_n231), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n218), .A2(new_n234), .A3(new_n228), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT28), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n228), .A2(KEYINPUT69), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n221), .A2(new_n227), .A3(new_n241), .A4(new_n223), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n234), .A3(new_n218), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n236), .B(new_n239), .C1(new_n244), .C2(new_n238), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G101), .ZN(new_n246));
  NOR2_X1   g060(.A1(G237), .A2(G953), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G210), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n246), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n243), .A2(KEYINPUT30), .A3(new_n218), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT68), .B1(new_n229), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  AOI211_X1 g071(.A(new_n257), .B(new_n254), .C1(new_n218), .C2(new_n228), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n253), .B(new_n235), .C1(new_n256), .C2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n218), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n240), .B2(new_n242), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n251), .B1(new_n261), .B2(new_n234), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT31), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n259), .A2(KEYINPUT31), .A3(new_n262), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n252), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(G472), .A2(G902), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n188), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n245), .A2(new_n251), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n259), .A2(KEYINPUT31), .A3(new_n262), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT31), .B1(new_n259), .B2(new_n262), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT32), .A3(new_n268), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n245), .B2(new_n251), .ZN(new_n278));
  INV_X1    g092(.A(new_n251), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(new_n259), .B2(new_n244), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n276), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n239), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(KEYINPUT29), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n244), .A2(KEYINPUT72), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n243), .A2(new_n218), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n235), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n261), .A2(new_n287), .A3(new_n234), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n284), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  AOI211_X1 g103(.A(new_n282), .B(new_n283), .C1(new_n289), .C2(KEYINPUT28), .ZN(new_n290));
  OAI21_X1  g104(.A(G472), .B1(new_n281), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n270), .A2(new_n275), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT25), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT16), .ZN(new_n294));
  INV_X1    g108(.A(G140), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(G125), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(G125), .ZN(new_n297));
  INV_X1    g111(.A(G125), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G140), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n296), .B1(new_n300), .B2(new_n294), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n189), .ZN(new_n302));
  OAI211_X1 g116(.A(G146), .B(new_n296), .C1(new_n300), .C2(new_n294), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(KEYINPUT74), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(new_n305), .A3(new_n189), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n203), .A2(G119), .ZN(new_n307));
  INV_X1    g121(.A(G119), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G128), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT24), .B(G110), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n307), .B1(KEYINPUT73), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT73), .B(KEYINPUT23), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n314), .B(new_n309), .C1(new_n315), .C2(new_n307), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n312), .B1(new_n316), .B2(G110), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n304), .A2(new_n306), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n189), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n303), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n316), .A2(G110), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n310), .A2(new_n311), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT75), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n310), .A2(new_n311), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n321), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n318), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G953), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G221), .A3(G234), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G137), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n333), .A2(KEYINPUT76), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(KEYINPUT76), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n333), .A2(KEYINPUT76), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n210), .A2(KEYINPUT22), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT22), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G137), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT76), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n337), .A2(new_n341), .A3(KEYINPUT77), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n331), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n334), .A2(new_n332), .A3(new_n335), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT77), .B1(new_n337), .B2(new_n341), .ZN(new_n345));
  INV_X1    g159(.A(new_n331), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n329), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n318), .A2(new_n328), .A3(new_n347), .A4(new_n343), .ZN(new_n350));
  AOI21_X1  g164(.A(G902), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n293), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AND4_X1   g167(.A1(new_n318), .A2(new_n328), .A3(new_n347), .A4(new_n343), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n318), .A2(new_n328), .B1(new_n343), .B2(new_n347), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n276), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n357));
  INV_X1    g171(.A(G217), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(G234), .B2(new_n276), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n354), .A2(new_n355), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n359), .A2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n292), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(G234), .A2(G237), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n367), .A2(G952), .A3(new_n330), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n367), .A2(G902), .A3(G953), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT21), .B(G898), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G478), .ZN(new_n373));
  NOR2_X1   g187(.A1(KEYINPUT98), .A2(KEYINPUT15), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT98), .A2(KEYINPUT15), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  INV_X1    g193(.A(G122), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G116), .ZN(new_n381));
  INV_X1    g195(.A(G116), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G122), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n383), .A3(KEYINPUT95), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT95), .B1(new_n381), .B2(new_n383), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n379), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G128), .B(G143), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(new_n208), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n382), .A2(KEYINPUT14), .A3(G122), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n381), .A2(new_n383), .ZN(new_n391));
  OAI211_X1 g205(.A(G107), .B(new_n390), .C1(new_n391), .C2(KEYINPUT14), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n387), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  OR2_X1    g207(.A1(KEYINPUT96), .A2(KEYINPUT13), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT96), .A2(KEYINPUT13), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n394), .B(new_n395), .C1(G128), .C2(new_n191), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G134), .ZN(new_n397));
  INV_X1    g211(.A(new_n388), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(G134), .A3(new_n388), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT95), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n391), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n384), .A3(G107), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n387), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT97), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n406), .B1(new_n401), .B2(new_n405), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n393), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT9), .B(G234), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n411), .A2(new_n358), .A3(G953), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n385), .A2(new_n379), .A3(new_n386), .ZN(new_n415));
  AOI21_X1  g229(.A(G107), .B1(new_n403), .B2(new_n384), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n396), .A2(G134), .A3(new_n388), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n388), .B1(new_n396), .B2(G134), .ZN(new_n418));
  OAI22_X1  g232(.A1(new_n415), .A2(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT97), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n407), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n393), .A3(new_n412), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n378), .B1(new_n423), .B2(new_n276), .ZN(new_n424));
  AOI211_X1 g238(.A(G902), .B(new_n377), .C1(new_n414), .C2(new_n422), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(new_n191), .ZN(new_n428));
  NOR2_X1   g242(.A1(KEYINPUT90), .A2(G143), .ZN(new_n429));
  OAI211_X1 g243(.A(G214), .B(new_n247), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n247), .A2(G214), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n427), .B2(new_n191), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n432), .A3(new_n212), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT91), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n430), .A2(new_n432), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G131), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT17), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n430), .A2(new_n432), .A3(KEYINPUT91), .A4(new_n212), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n435), .A2(new_n437), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n304), .A2(new_n306), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n436), .A2(KEYINPUT17), .A3(G131), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  XOR2_X1   g257(.A(G113), .B(G122), .Z(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT93), .B(G104), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n300), .A2(G146), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n320), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT18), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(new_n212), .ZN(new_n450));
  OAI221_X1 g264(.A(new_n448), .B1(new_n436), .B2(new_n450), .C1(new_n437), .C2(new_n449), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n443), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n446), .B1(new_n443), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n276), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT94), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(KEYINPUT94), .B(new_n276), .C1(new_n452), .C2(new_n453), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(G475), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G475), .A2(G902), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n435), .A2(new_n437), .A3(new_n439), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n319), .B(KEYINPUT19), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n189), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT92), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(KEYINPUT92), .A3(new_n189), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n460), .A2(new_n464), .A3(new_n303), .A4(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n446), .B1(new_n466), .B2(new_n451), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n459), .B1(new_n452), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT20), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n470), .B(new_n459), .C1(new_n452), .C2(new_n467), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AND4_X1   g286(.A1(new_n372), .A2(new_n426), .A3(new_n458), .A4(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G221), .B1(new_n411), .B2(G902), .ZN(new_n474));
  XOR2_X1   g288(.A(new_n474), .B(KEYINPUT79), .Z(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G110), .B(G140), .ZN(new_n477));
  INV_X1    g291(.A(G227), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(G953), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n477), .B(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n221), .A2(new_n223), .ZN(new_n481));
  INV_X1    g295(.A(G101), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n379), .A2(G104), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT81), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n379), .A2(G104), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n484), .B1(new_n485), .B2(KEYINPUT3), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT3), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n487), .A2(new_n379), .A3(KEYINPUT81), .A4(G104), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n483), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT80), .ZN(new_n490));
  INV_X1    g304(.A(G104), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(G107), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n490), .B1(new_n492), .B2(new_n487), .ZN(new_n493));
  OAI211_X1 g307(.A(KEYINPUT80), .B(KEYINPUT3), .C1(new_n491), .C2(G107), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n482), .B1(new_n489), .B2(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT84), .B(KEYINPUT4), .Z(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n227), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI211_X1 g314(.A(KEYINPUT82), .B(new_n482), .C1(new_n489), .C2(new_n495), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n486), .A2(new_n488), .ZN(new_n502));
  INV_X1    g316(.A(new_n483), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n495), .A2(new_n502), .A3(new_n482), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT81), .B1(new_n492), .B2(new_n487), .ZN(new_n507));
  INV_X1    g321(.A(new_n488), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n494), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT80), .B1(new_n485), .B2(KEYINPUT3), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G101), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT82), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT83), .B1(new_n506), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT82), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n516), .B(G101), .C1(new_n509), .C2(new_n512), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(KEYINPUT4), .A3(new_n504), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT83), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n496), .A2(new_n516), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n500), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n198), .A2(new_n205), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT10), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G101), .B1(new_n492), .B2(new_n483), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n504), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n203), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n205), .B1(new_n202), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n531), .A2(new_n504), .A3(new_n526), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n529), .B1(KEYINPUT10), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n481), .B1(new_n522), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n519), .B1(new_n518), .B2(new_n520), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n537), .A2(new_n514), .A3(KEYINPUT83), .A4(new_n517), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n499), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n481), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n539), .A2(new_n540), .A3(new_n533), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n480), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n522), .A2(new_n481), .A3(new_n534), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT86), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n206), .B1(new_n504), .B2(new_n526), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n540), .B1(new_n532), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n481), .B2(KEYINPUT85), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n527), .A2(new_n523), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n531), .A2(new_n504), .A3(new_n526), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n481), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(new_n548), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n544), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n480), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n546), .A2(new_n549), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n548), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT86), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n543), .A2(new_n555), .A3(new_n556), .A4(new_n559), .ZN(new_n560));
  AOI211_X1 g374(.A(G469), .B(G902), .C1(new_n542), .C2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n550), .A2(new_n554), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n480), .B1(new_n541), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n540), .B1(new_n539), .B2(new_n533), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n543), .A2(new_n564), .A3(new_n556), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(G469), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(G469), .A2(G902), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n473), .B(new_n476), .C1(new_n561), .C2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G214), .B1(G237), .B2(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n498), .A2(new_n235), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n515), .B2(new_n521), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n231), .A2(KEYINPUT5), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n382), .A2(KEYINPUT5), .A3(G119), .ZN(new_n575));
  INV_X1    g389(.A(G113), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n232), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n528), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(G110), .B(G122), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n580), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n571), .B1(new_n536), .B2(new_n538), .ZN(new_n583));
  INV_X1    g397(.A(new_n579), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n581), .A2(new_n585), .A3(KEYINPUT6), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n206), .A2(new_n298), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n227), .A2(G125), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G224), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n589), .B1(new_n590), .B2(G953), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(G953), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n587), .A2(new_n592), .A3(new_n588), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT6), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n595), .B(new_n582), .C1(new_n583), .C2(new_n584), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n586), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n528), .A2(new_n578), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT87), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n580), .B(KEYINPUT8), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT87), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n579), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n599), .B(new_n600), .C1(new_n602), .C2(new_n598), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT88), .B(KEYINPUT7), .Z(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n587), .B(new_n588), .C1(new_n592), .C2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT89), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n589), .B(KEYINPUT7), .C1(new_n590), .C2(G953), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n603), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n610), .B2(new_n581), .ZN(new_n611));
  OAI21_X1  g425(.A(G210), .B1(G237), .B2(G902), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n597), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n612), .B1(new_n597), .B2(new_n611), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n570), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n366), .A2(new_n569), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(new_n482), .ZN(G3));
  AOI21_X1  g431(.A(G478), .B1(new_n423), .B2(new_n276), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n412), .B1(new_n421), .B2(new_n393), .ZN(new_n619));
  INV_X1    g433(.A(new_n393), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n620), .B(new_n413), .C1(new_n420), .C2(new_n407), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT99), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n423), .A2(KEYINPUT99), .A3(KEYINPUT33), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n373), .A2(G902), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n618), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(G475), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n454), .B2(new_n455), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n630), .A2(new_n457), .B1(new_n469), .B2(new_n471), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n628), .A2(new_n631), .A3(new_n371), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n615), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n365), .B(new_n476), .C1(new_n561), .C2(new_n568), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n274), .A2(new_n276), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n274), .A2(new_n268), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NAND2_X1  g457(.A1(new_n458), .A2(new_n472), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n644), .A2(new_n371), .A3(new_n426), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n645), .B(new_n570), .C1(new_n613), .C2(new_n614), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n569), .A2(new_n615), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n636), .A2(G472), .B1(new_n268), .B2(new_n274), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT36), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n336), .A2(new_n342), .A3(new_n331), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n346), .B1(new_n344), .B2(new_n345), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n329), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n348), .A2(new_n653), .A3(new_n318), .A4(new_n328), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n658), .A3(new_n363), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n360), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n652), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n651), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT101), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT37), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  AND2_X1   g482(.A1(new_n566), .A2(new_n567), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n542), .A2(new_n560), .ZN(new_n670));
  INV_X1    g484(.A(G469), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n671), .A3(new_n276), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n475), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n292), .A3(new_n662), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n424), .A2(new_n425), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n631), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n369), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n368), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n682), .B(new_n570), .C1(new_n614), .C2(new_n613), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n203), .ZN(G30));
  INV_X1    g499(.A(new_n570), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n631), .A2(new_n686), .A3(new_n426), .ZN(new_n687));
  INV_X1    g501(.A(new_n662), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n644), .A2(new_n570), .A3(new_n675), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n662), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT102), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n289), .A2(new_n251), .B1(new_n259), .B2(new_n262), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n695), .B2(G902), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n270), .A2(new_n275), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n691), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT38), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n613), .B2(new_n614), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n597), .A2(new_n611), .ZN(new_n702));
  INV_X1    g516(.A(new_n612), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n597), .A2(new_n611), .A3(new_n612), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n704), .A2(KEYINPUT38), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  OR3_X1    g521(.A1(new_n698), .A2(new_n699), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n680), .B(KEYINPUT39), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n673), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n710), .B(KEYINPUT40), .Z(new_n711));
  OAI21_X1  g525(.A(new_n699), .B1(new_n698), .B2(new_n707), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n708), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  NOR3_X1   g528(.A1(new_n628), .A2(new_n631), .A3(new_n681), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n715), .B(new_n570), .C1(new_n614), .C2(new_n613), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n674), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n189), .ZN(G48));
  NAND2_X1  g532(.A1(new_n543), .A2(new_n564), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT86), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT86), .B1(new_n557), .B2(new_n558), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n536), .A2(new_n538), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n533), .B1(new_n723), .B2(new_n500), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n480), .B1(new_n724), .B2(new_n481), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n719), .A2(new_n480), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(G469), .B1(new_n726), .B2(G902), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n476), .A3(new_n672), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n366), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n634), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  INV_X1    g546(.A(new_n366), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n727), .A2(new_n476), .A3(new_n672), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n647), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  AND3_X1   g550(.A1(new_n292), .A2(new_n473), .A3(new_n662), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n615), .A2(new_n728), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  NAND4_X1  g554(.A1(new_n727), .A2(new_n476), .A3(new_n672), .A4(new_n372), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n687), .B1(new_n613), .B2(new_n614), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g557(.A(KEYINPUT104), .B(G472), .Z(new_n744));
  NAND2_X1  g558(.A1(new_n636), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n289), .A2(KEYINPUT28), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n279), .B1(new_n746), .B2(new_n239), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n272), .A2(new_n273), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n268), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n745), .A2(new_n365), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  NAND4_X1  g567(.A1(new_n715), .A2(new_n662), .A3(new_n749), .A4(new_n745), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n738), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT32), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n267), .A2(new_n759), .A3(new_n269), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT32), .B1(new_n274), .B2(new_n268), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT105), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n759), .B1(new_n267), .B2(new_n269), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n275), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n291), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n365), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n613), .A2(new_n614), .A3(new_n686), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n673), .A3(KEYINPUT42), .A4(new_n715), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n758), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n365), .ZN(new_n771));
  INV_X1    g585(.A(new_n291), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n763), .A2(new_n275), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n772), .B1(new_n773), .B2(KEYINPUT105), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n771), .B1(new_n774), .B2(new_n765), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n715), .A2(KEYINPUT42), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n704), .A2(new_n570), .A3(new_n705), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n476), .B1(new_n561), .B2(new_n568), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(KEYINPUT106), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n777), .A2(new_n778), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n733), .A2(new_n782), .A3(new_n715), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n770), .A2(new_n780), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT107), .B(G131), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G33));
  NAND3_X1  g600(.A1(new_n733), .A2(new_n782), .A3(new_n682), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  AOI21_X1  g602(.A(KEYINPUT45), .B1(new_n563), .B2(new_n565), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n671), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n563), .A2(KEYINPUT45), .A3(new_n565), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n567), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(KEYINPUT46), .A3(new_n567), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n672), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n476), .A3(new_n709), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT108), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT108), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n797), .A2(new_n800), .A3(new_n476), .A4(new_n709), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT43), .B1(new_n628), .B2(new_n644), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT43), .ZN(new_n804));
  INV_X1    g618(.A(new_n627), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n624), .B2(new_n625), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n631), .B(new_n804), .C1(new_n618), .C2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n803), .A2(new_n662), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n808), .A2(new_n809), .A3(new_n652), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n809), .B1(new_n808), .B2(new_n652), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n768), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT109), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT109), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n810), .A2(new_n814), .A3(new_n768), .A4(new_n811), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n802), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g631(.A(KEYINPUT110), .B(G137), .Z(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(G39));
  NAND2_X1  g633(.A1(new_n797), .A2(new_n476), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT47), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n797), .A2(KEYINPUT47), .A3(new_n476), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n715), .A2(new_n771), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n777), .A3(new_n292), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT111), .Z(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  NAND2_X1  g643(.A1(new_n783), .A2(new_n781), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n767), .A2(new_n758), .A3(new_n769), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT106), .B1(new_n775), .B2(new_n779), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n730), .A2(new_n735), .A3(new_n739), .A4(new_n752), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n292), .A2(new_n662), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n631), .A2(new_n426), .A3(new_n680), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n754), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n782), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n787), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n686), .B1(new_n704), .B2(new_n705), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n673), .A3(new_n473), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n673), .A2(new_n365), .A3(new_n652), .ZN(new_n844));
  OAI22_X1  g658(.A1(new_n843), .A2(new_n663), .B1(new_n844), .B2(new_n646), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n733), .A2(new_n651), .B1(new_n634), .B2(new_n640), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n842), .A2(new_n632), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT114), .B1(new_n850), .B2(new_n616), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n848), .A2(KEYINPUT115), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n641), .B(new_n847), .C1(new_n366), .C2(new_n843), .ZN(new_n854));
  INV_X1    g668(.A(new_n845), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n851), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n841), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n692), .B1(new_n704), .B2(new_n705), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n360), .A2(new_n661), .A3(new_n680), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n360), .A2(new_n661), .A3(KEYINPUT116), .A4(new_n680), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n861), .A2(new_n673), .A3(new_n697), .A4(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n674), .B2(new_n716), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n835), .A2(new_n778), .ZN(new_n870));
  INV_X1    g684(.A(new_n683), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n870), .A2(new_n871), .B1(new_n755), .B2(new_n738), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n860), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n869), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n734), .A2(new_n842), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n876), .A2(new_n754), .B1(new_n674), .B2(new_n683), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT117), .B1(new_n877), .B2(new_n868), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n873), .B1(new_n879), .B2(new_n860), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT53), .B1(new_n859), .B2(new_n880), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n729), .A2(new_n647), .B1(new_n737), .B2(new_n738), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n729), .A2(new_n634), .B1(new_n743), .B2(new_n751), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n882), .A2(new_n883), .A3(new_n787), .A4(new_n838), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n784), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT115), .B1(new_n848), .B2(new_n851), .ZN(new_n886));
  AND4_X1   g700(.A1(KEYINPUT115), .A2(new_n851), .A3(new_n854), .A4(new_n855), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n874), .B1(new_n869), .B2(new_n872), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n877), .A2(new_n868), .A3(KEYINPUT117), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n860), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n875), .A2(KEYINPUT52), .A3(new_n878), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n888), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT54), .B1(new_n881), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n880), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n894), .B1(new_n888), .B2(new_n893), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n734), .A2(KEYINPUT118), .A3(new_n768), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n777), .B2(new_n728), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n803), .A2(new_n368), .A3(new_n807), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n901), .B1(new_n907), .B2(new_n767), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n901), .A3(new_n767), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT48), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n901), .B(KEYINPUT48), .C1(new_n907), .C2(new_n767), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n905), .A2(new_n750), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(G952), .B(new_n330), .C1(new_n915), .C2(new_n876), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n697), .A2(new_n771), .A3(new_n679), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n902), .A2(new_n904), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n628), .A2(new_n631), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n644), .A2(new_n618), .A3(new_n806), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n902), .A2(new_n904), .A3(new_n917), .A4(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n745), .A2(new_n662), .A3(new_n749), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n902), .A2(new_n904), .A3(new_n923), .A4(new_n906), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n914), .A2(new_n686), .A3(new_n707), .A4(new_n734), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT50), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n922), .B(new_n924), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n727), .A2(new_n672), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT112), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n475), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n822), .A2(new_n823), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n915), .A2(new_n777), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n913), .B(new_n920), .C1(new_n935), .C2(KEYINPUT51), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n925), .B(new_n926), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n922), .A2(new_n924), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n922), .B2(new_n924), .ZN(new_n941));
  OAI211_X1 g755(.A(KEYINPUT120), .B(new_n937), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n933), .A2(new_n934), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(KEYINPUT51), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n941), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n939), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT120), .B1(new_n946), .B2(new_n937), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n936), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n896), .A2(new_n900), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT122), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT122), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n896), .A2(new_n949), .A3(new_n952), .A4(new_n900), .ZN(new_n953));
  INV_X1    g767(.A(G952), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n330), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n931), .B(KEYINPUT49), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n697), .A2(new_n771), .ZN(new_n958));
  NOR4_X1   g772(.A1(new_n628), .A2(new_n644), .A3(new_n686), .A4(new_n475), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n957), .A2(new_n707), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT113), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n956), .A2(new_n961), .ZN(G75));
  NOR2_X1   g776(.A1(new_n330), .A2(G952), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n276), .B1(new_n897), .B2(new_n898), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT56), .B1(new_n965), .B2(G210), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n586), .A2(new_n596), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(new_n594), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT55), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n964), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n966), .B2(new_n970), .ZN(G51));
  XOR2_X1   g786(.A(new_n567), .B(KEYINPUT57), .Z(new_n973));
  INV_X1    g787(.A(new_n900), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n670), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n965), .A2(new_n791), .A3(new_n790), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n963), .B1(new_n977), .B2(new_n978), .ZN(G54));
  NAND3_X1  g793(.A1(new_n965), .A2(KEYINPUT58), .A3(G475), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n452), .A2(new_n467), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n982), .A2(new_n983), .A3(new_n963), .ZN(G60));
  NAND2_X1  g798(.A1(G478), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT59), .Z(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n626), .B(new_n987), .C1(new_n974), .C2(new_n975), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n964), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n896), .A2(new_n900), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n626), .B1(new_n990), .B2(new_n987), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n989), .A2(new_n991), .ZN(G63));
  INV_X1    g806(.A(KEYINPUT61), .ZN(new_n993));
  XNOR2_X1  g807(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n994));
  NAND2_X1  g808(.A1(G217), .A2(G902), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n897), .B2(new_n898), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(new_n657), .A3(new_n658), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n964), .B1(new_n997), .B2(new_n362), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n993), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n997), .A2(new_n362), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1002), .A2(KEYINPUT61), .A3(new_n964), .A4(new_n998), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(G66));
  OAI21_X1  g818(.A(G953), .B1(new_n370), .B2(new_n590), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n883), .B(new_n882), .C1(new_n886), .C2(new_n887), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1005), .B1(new_n1007), .B2(G953), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n967), .B1(G898), .B2(new_n330), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(G69));
  INV_X1    g824(.A(KEYINPUT62), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n877), .A2(new_n717), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n713), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n676), .B1(new_n631), .B2(new_n628), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n733), .A2(new_n782), .A3(new_n709), .A4(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n817), .A2(new_n1013), .A3(new_n828), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT125), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n713), .A2(new_n1012), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1017), .B1(new_n1018), .B2(KEYINPUT62), .ZN(new_n1019));
  AOI211_X1 g833(.A(KEYINPUT125), .B(new_n1011), .C1(new_n713), .C2(new_n1012), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n253), .B1(new_n256), .B2(new_n258), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT124), .Z(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(new_n461), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n767), .A2(new_n742), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n802), .B1(new_n816), .B2(new_n1027), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n1012), .A2(new_n787), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1028), .A2(new_n833), .A3(new_n828), .A4(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1030), .A2(new_n1025), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1031), .A2(G953), .ZN(new_n1032));
  OR2_X1    g846(.A1(new_n1025), .A2(new_n478), .ZN(new_n1033));
  AOI211_X1 g847(.A(new_n677), .B(new_n330), .C1(new_n1025), .C2(new_n478), .ZN(new_n1034));
  AOI22_X1  g848(.A1(new_n1026), .A2(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(G72));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1038), .B1(new_n1021), .B2(new_n1007), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n259), .A2(new_n244), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT126), .Z(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n279), .ZN(new_n1042));
  OR2_X1    g856(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n881), .A2(new_n895), .ZN(new_n1044));
  INV_X1    g858(.A(new_n263), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1037), .B1(new_n1045), .B2(new_n280), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1037), .B1(new_n1030), .B2(new_n1006), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n1041), .A2(new_n279), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n963), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g865(.A1(new_n1043), .A2(new_n1048), .A3(KEYINPUT127), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT127), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1051), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1053), .B1(new_n1054), .B2(new_n1047), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1052), .A2(new_n1055), .ZN(G57));
endmodule


