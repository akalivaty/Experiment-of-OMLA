//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT65), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n193), .A3(new_n194), .A4(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n190), .A2(KEYINPUT64), .A3(G143), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(new_n192), .B2(G146), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n192), .A2(G146), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n200), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n194), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n189), .B1(new_n199), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT88), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n211), .A2(new_n191), .A3(new_n193), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n212), .B1(new_n204), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n208), .A2(new_n209), .B1(new_n189), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n196), .A2(new_n198), .B1(new_n204), .B2(new_n206), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT88), .B1(new_n221), .B2(new_n189), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G953), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G224), .ZN(new_n225));
  XOR2_X1   g039(.A(new_n225), .B(KEYINPUT89), .Z(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n223), .B(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n231));
  INV_X1    g045(.A(G107), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(G104), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(G107), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G101), .ZN(new_n236));
  INV_X1    g050(.A(G101), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n230), .A2(new_n233), .A3(new_n237), .A4(new_n234), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(KEYINPUT4), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G119), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(KEYINPUT68), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT2), .B(G113), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n236), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(new_n238), .ZN(new_n246));
  OR2_X1    g060(.A1(new_n236), .A2(KEYINPUT4), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n245), .A3(new_n246), .A4(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G119), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G116), .ZN(new_n250));
  INV_X1    g064(.A(G116), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G119), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT5), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT5), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n249), .A3(G116), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n253), .A2(KEYINPUT87), .A3(G113), .A4(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT2), .B(G113), .Z(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n242), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n255), .A2(G113), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT87), .B1(new_n260), .B2(new_n253), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n229), .A2(G107), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n232), .A2(G104), .ZN(new_n263));
  OAI21_X1  g077(.A(G101), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n238), .A2(new_n264), .ZN(new_n265));
  OR3_X1    g079(.A1(new_n259), .A2(new_n261), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n248), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G122), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n270), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n248), .A2(new_n266), .A3(new_n269), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(KEYINPUT6), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n228), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n226), .A2(KEYINPUT7), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n199), .A2(new_n207), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n209), .A3(G125), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n219), .A2(new_n189), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n208), .A2(new_n209), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT7), .A4(new_n226), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n260), .A2(new_n253), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n258), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT91), .B1(new_n285), .B2(new_n265), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n265), .B1(new_n259), .B2(new_n261), .ZN(new_n287));
  INV_X1    g101(.A(new_n265), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT91), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n284), .A4(new_n258), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n286), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT90), .B(KEYINPUT8), .Z(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(new_n269), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n282), .A2(new_n283), .A3(new_n273), .A4(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT92), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n275), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G210), .B1(G237), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n301), .B(new_n275), .C1(new_n298), .C2(new_n299), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n188), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT96), .ZN(new_n306));
  XNOR2_X1  g120(.A(G113), .B(G122), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(new_n229), .ZN(new_n308));
  INV_X1    g122(.A(G140), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n189), .A2(G140), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT19), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT19), .B1(new_n310), .B2(new_n311), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n190), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT16), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n309), .A3(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(new_n311), .ZN(new_n317));
  OAI211_X1 g131(.A(G146), .B(new_n316), .C1(new_n317), .C2(new_n315), .ZN(new_n318));
  NOR2_X1   g132(.A1(G237), .A2(G953), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G214), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT93), .A2(G143), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n319), .B(G214), .C1(KEYINPUT93), .C2(G143), .ZN(new_n323));
  INV_X1    g137(.A(G131), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n324), .B1(new_n322), .B2(new_n323), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n314), .B(new_n318), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(KEYINPUT18), .A2(G131), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n322), .B2(new_n323), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n310), .A2(new_n311), .A3(new_n190), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n190), .B1(new_n310), .B2(new_n311), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n322), .A2(new_n323), .A3(new_n329), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n331), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n308), .B1(new_n328), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n336), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n333), .A2(new_n334), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n339), .A2(new_n340), .A3(new_n330), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n322), .A2(new_n323), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT17), .A3(G131), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n316), .B1(new_n317), .B2(new_n315), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n190), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n343), .A2(new_n345), .A3(new_n318), .ZN(new_n346));
  INV_X1    g160(.A(new_n327), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT17), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(new_n325), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n341), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n338), .B1(new_n350), .B2(new_n308), .ZN(new_n351));
  INV_X1    g165(.A(G475), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n297), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT20), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n355));
  NOR2_X1   g169(.A1(G475), .A2(G902), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT17), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n343), .A2(new_n345), .A3(new_n318), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n308), .B(new_n337), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n355), .B(new_n356), .C1(new_n360), .C2(new_n338), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n350), .A2(new_n308), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n297), .B1(new_n363), .B2(new_n360), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT94), .B(G475), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT9), .B(G234), .ZN(new_n367));
  INV_X1    g181(.A(G217), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n367), .A2(new_n368), .A3(G953), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G122), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G116), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n251), .A2(G122), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n372), .B(new_n373), .C1(KEYINPUT14), .C2(new_n232), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n232), .B1(new_n372), .B2(KEYINPUT14), .ZN(new_n375));
  INV_X1    g189(.A(new_n372), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n371), .A2(G116), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n213), .A2(new_n215), .A3(G143), .ZN(new_n379));
  INV_X1    g193(.A(G134), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n192), .A2(G128), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n380), .B1(new_n379), .B2(new_n381), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n374), .B(new_n378), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT13), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n192), .A2(KEYINPUT13), .A3(G128), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n379), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G134), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n372), .A2(new_n373), .A3(G107), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n232), .B1(new_n376), .B2(new_n377), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n390), .A2(new_n382), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT95), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n385), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n385), .B2(new_n393), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n370), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n385), .A2(new_n393), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT95), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n385), .A2(new_n393), .A3(new_n394), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n369), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n401), .A3(new_n297), .ZN(new_n402));
  INV_X1    g216(.A(G478), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT15), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n404), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n397), .A2(new_n401), .A3(new_n297), .A4(new_n406), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n362), .A2(new_n366), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(G234), .A2(G237), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n409), .A2(G952), .A3(new_n224), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n409), .A2(G902), .A3(G953), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT21), .B(G898), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n306), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n405), .A2(new_n407), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n413), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n354), .A2(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n416), .A2(KEYINPUT96), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n305), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n224), .A2(G227), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT82), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n204), .A2(new_n218), .ZN(new_n427));
  INV_X1    g241(.A(new_n212), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n265), .A3(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n217), .A2(G128), .B1(new_n191), .B2(new_n193), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n238), .B(new_n264), .C1(new_n430), .C2(new_n212), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT11), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n380), .B2(G137), .ZN(new_n434));
  INV_X1    g248(.A(G137), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT11), .A3(G134), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n380), .A2(G137), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G131), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n434), .A2(new_n436), .A3(new_n324), .A4(new_n437), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n432), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n429), .A2(KEYINPUT85), .A3(new_n431), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT85), .B1(new_n429), .B2(new_n431), .ZN(new_n447));
  INV_X1    g261(.A(new_n441), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n445), .B1(new_n449), .B2(KEYINPUT12), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n432), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n429), .A2(KEYINPUT85), .A3(new_n431), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n441), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT12), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(KEYINPUT86), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n444), .B1(new_n450), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT10), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n219), .A2(new_n458), .A3(new_n265), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n458), .B2(new_n431), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n241), .A2(new_n221), .A3(new_n246), .A4(new_n247), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(new_n448), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n426), .B1(new_n457), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n425), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n448), .B1(new_n460), .B2(new_n461), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n464), .A2(G469), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n450), .A2(new_n456), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n465), .B1(new_n471), .B2(new_n443), .ZN(new_n472));
  INV_X1    g286(.A(new_n466), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n425), .B1(new_n473), .B2(new_n462), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n470), .B(new_n297), .C1(new_n472), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(G469), .A2(G902), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n469), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G221), .B1(new_n367), .B2(G902), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(KEYINPUT81), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n421), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n368), .B1(G234), .B2(new_n297), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT25), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT24), .B(G110), .Z(new_n486));
  NAND3_X1  g300(.A1(new_n213), .A2(new_n215), .A3(G119), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n249), .A2(G128), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT78), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT78), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n486), .A2(new_n487), .A3(new_n491), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n345), .A2(new_n318), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT23), .B1(new_n210), .B2(G119), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(new_n249), .B2(G128), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT23), .A4(G119), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G110), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G110), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n496), .A2(new_n501), .A3(new_n497), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n318), .B(new_n332), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n224), .A2(G221), .A3(G234), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT79), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT22), .B(G137), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n500), .A2(new_n504), .A3(new_n509), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n485), .B1(new_n513), .B2(G902), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n511), .A2(KEYINPUT25), .A3(new_n297), .A4(new_n512), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n484), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n513), .A2(G902), .A3(new_n483), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT80), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n319), .A2(G210), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT27), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT26), .B(G101), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n527));
  NOR2_X1   g341(.A1(new_n380), .A2(G137), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n435), .A2(G134), .ZN(new_n529));
  OAI21_X1  g343(.A(G131), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n440), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n427), .B2(new_n428), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n532), .A2(new_n533), .B1(new_n221), .B2(new_n441), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT70), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n243), .B(new_n257), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT69), .B1(new_n219), .B2(new_n531), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n440), .A2(new_n530), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT64), .B1(new_n190), .B2(G143), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n191), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n541), .A2(new_n200), .B1(new_n216), .B2(new_n217), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n539), .B(new_n533), .C1(new_n542), .C2(new_n212), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n441), .A2(new_n207), .A3(new_n199), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n537), .A2(new_n543), .A3(new_n536), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT70), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n440), .B(new_n530), .C1(new_n542), .C2(new_n212), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n245), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n527), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n548), .A3(new_n536), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT28), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n526), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n534), .A2(KEYINPUT30), .A3(new_n537), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT67), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n549), .B2(new_n559), .ZN(new_n560));
  AOI211_X1 g374(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n544), .C2(new_n548), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n245), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n525), .A3(new_n547), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT31), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n565));
  NAND4_X1  g379(.A1(new_n562), .A2(new_n525), .A3(new_n547), .A4(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n556), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(G472), .A2(G902), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT73), .B(KEYINPUT32), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n521), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n564), .A2(new_n566), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n545), .A2(KEYINPUT70), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n545), .A2(KEYINPUT70), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n550), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n527), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n525), .B1(new_n577), .B2(new_n554), .ZN(new_n578));
  OAI211_X1 g392(.A(KEYINPUT32), .B(new_n568), .C1(new_n572), .C2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n570), .B1(new_n567), .B2(new_n568), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT74), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G472), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT75), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n555), .A2(new_n526), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n584), .B1(new_n551), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n538), .A2(new_n546), .B1(new_n245), .B2(new_n549), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n585), .B(KEYINPUT75), .C1(new_n588), .C2(new_n527), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT29), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n562), .A2(new_n547), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n526), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n587), .A2(new_n589), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n538), .A2(new_n546), .A3(KEYINPUT76), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n534), .A2(new_n537), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n245), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT76), .B1(new_n538), .B2(new_n546), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT28), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n586), .A2(new_n590), .ZN(new_n600));
  AOI21_X1  g414(.A(G902), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n583), .B1(new_n593), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(KEYINPUT77), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT77), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n604), .B(new_n583), .C1(new_n593), .C2(new_n601), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n482), .B(new_n520), .C1(new_n582), .C2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT97), .B(G101), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G3));
  NAND2_X1  g423(.A1(new_n397), .A2(new_n401), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n397), .A2(new_n401), .A3(KEYINPUT33), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n403), .A2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n402), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n616), .B1(G478), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n418), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(new_n305), .A3(new_n417), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n620), .A2(new_n305), .A3(KEYINPUT98), .A4(new_n417), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n567), .A2(new_n297), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(G472), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n567), .A2(new_n568), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n519), .ZN(new_n631));
  INV_X1    g445(.A(new_n481), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(new_n305), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n413), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n361), .A2(KEYINPUT99), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n354), .A2(new_n361), .A3(KEYINPUT99), .ZN(new_n640));
  AND4_X1   g454(.A1(new_n366), .A2(new_n415), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n633), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT35), .B(G107), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NOR2_X1   g460(.A1(new_n421), .A2(new_n630), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n483), .A2(G902), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n510), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n505), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n516), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n477), .A2(new_n480), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  AOI211_X1 g471(.A(new_n521), .B(new_n570), .C1(new_n567), .C2(new_n568), .ZN(new_n658));
  INV_X1    g472(.A(new_n579), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n660), .B(new_n571), .C1(new_n603), .C2(new_n605), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n411), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n410), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n364), .B2(new_n365), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n415), .A2(new_n639), .A3(new_n640), .A4(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n637), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n661), .A2(new_n654), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  NAND2_X1  g487(.A1(new_n591), .A2(new_n525), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n297), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n597), .A2(new_n525), .A3(new_n598), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n660), .A2(new_n571), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT101), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n303), .A2(new_n304), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT38), .Z(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n416), .A2(new_n188), .A3(new_n418), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n651), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n665), .B(KEYINPUT39), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n632), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n688));
  OR4_X1    g502(.A1(new_n679), .A2(new_n684), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT102), .B(G143), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G45));
  INV_X1    g505(.A(new_n418), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n618), .A2(new_n692), .A3(new_n665), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n637), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n661), .A2(new_n654), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  AND3_X1   g510(.A1(new_n454), .A2(KEYINPUT86), .A3(new_n455), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT86), .B1(new_n454), .B2(new_n455), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n443), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n465), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n474), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n701), .B2(G902), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n702), .A2(new_n480), .A3(new_n475), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n661), .A2(new_n520), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n626), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT41), .B(G113), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NOR2_X1   g521(.A1(new_n704), .A2(new_n643), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n251), .ZN(G18));
  AOI21_X1  g523(.A(new_n651), .B1(new_n414), .B2(new_n419), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n703), .A2(new_n305), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(new_n582), .B2(new_n606), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  XOR2_X1   g527(.A(new_n568), .B(KEYINPUT103), .Z(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n599), .A2(new_n554), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n526), .ZN(new_n717));
  INV_X1    g531(.A(new_n572), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n514), .A2(new_n515), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n483), .ZN(new_n722));
  INV_X1    g536(.A(new_n517), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n720), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n516), .A2(KEYINPUT105), .A3(new_n517), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT104), .B(G472), .Z(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n567), .B2(new_n297), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n719), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n299), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n301), .B1(new_n732), .B2(new_n275), .ZN(new_n733));
  INV_X1    g547(.A(new_n304), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n683), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n702), .A2(new_n475), .A3(new_n480), .A4(new_n417), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n729), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  NOR2_X1   g553(.A1(new_n719), .A2(new_n728), .ZN(new_n740));
  INV_X1    g554(.A(new_n693), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n652), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n703), .A2(new_n305), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n189), .ZN(G27));
  NAND4_X1  g559(.A1(new_n464), .A2(KEYINPUT106), .A3(G469), .A4(new_n468), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n475), .A3(new_n476), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n699), .A2(new_n462), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n467), .B1(new_n748), .B2(new_n426), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT106), .B1(new_n749), .B2(G469), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n480), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g567(.A(KEYINPUT107), .B(new_n480), .C1(new_n747), .C2(new_n750), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n303), .A2(new_n187), .A3(new_n304), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT32), .B1(new_n567), .B2(new_n568), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n759), .B2(new_n579), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT32), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n629), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n602), .B(KEYINPUT77), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n726), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n693), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n757), .A2(KEYINPUT109), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n579), .A2(new_n759), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n629), .A2(new_n761), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n773), .B(new_n762), .C1(new_n603), .C2(new_n605), .ZN(new_n774));
  INV_X1    g588(.A(new_n726), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n775), .A3(new_n768), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n770), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n580), .A2(KEYINPUT74), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n779), .A2(new_n658), .A3(new_n659), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n519), .B1(new_n780), .B2(new_n765), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n755), .B1(new_n751), .B2(new_n752), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n741), .A3(new_n754), .A4(new_n782), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n769), .A2(new_n778), .B1(new_n783), .B2(new_n767), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n324), .ZN(G33));
  INV_X1    g599(.A(new_n670), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n757), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  NAND2_X1  g602(.A1(new_n464), .A2(new_n468), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n470), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT46), .B1(new_n792), .B2(new_n476), .ZN(new_n793));
  INV_X1    g607(.A(new_n475), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(KEYINPUT46), .A3(new_n476), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n479), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n685), .ZN(new_n798));
  XNOR2_X1  g612(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n619), .B2(new_n692), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n692), .A2(KEYINPUT111), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n692), .A2(KEYINPUT111), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(KEYINPUT43), .A3(new_n618), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n630), .A3(new_n652), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT44), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n755), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n806), .B2(new_n805), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n798), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n435), .ZN(G39));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n797), .B(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n520), .A2(new_n693), .A3(new_n755), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n765), .A3(new_n780), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT112), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n811), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n797), .B(KEYINPUT47), .ZN(new_n818));
  INV_X1    g632(.A(new_n816), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(KEYINPUT113), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G140), .ZN(G42));
  NOR3_X1   g636(.A1(new_n726), .A2(new_n479), .A3(new_n188), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n801), .A2(new_n618), .A3(new_n802), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n702), .A2(new_n475), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n823), .B(new_n824), .C1(KEYINPUT49), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(KEYINPUT49), .B2(new_n825), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n679), .A2(new_n681), .A3(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT114), .Z(new_n829));
  AOI21_X1  g643(.A(new_n664), .B1(new_n800), .B2(new_n803), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n755), .A2(new_n825), .A3(new_n479), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n766), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT48), .Z(new_n833));
  AND3_X1   g647(.A1(new_n831), .A2(new_n520), .A3(new_n410), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n679), .A2(new_n620), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n830), .A2(new_n729), .ZN(new_n836));
  OAI211_X1 g650(.A(G952), .B(new_n224), .C1(new_n836), .C2(new_n743), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n833), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n702), .A2(new_n479), .A3(new_n475), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n813), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n836), .A2(new_n755), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n681), .A2(new_n188), .A3(new_n703), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT116), .B1(new_n845), .B2(new_n836), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT50), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n679), .A2(new_n418), .A3(new_n619), .A4(new_n834), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n830), .A2(new_n652), .A3(new_n740), .A4(new_n831), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT117), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  OR3_X1    g666(.A1(new_n848), .A2(new_n851), .A3(KEYINPUT117), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n844), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n851), .B(KEYINPUT118), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n848), .B1(new_n840), .B2(new_n841), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n843), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n838), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n661), .A2(new_n782), .A3(new_n520), .A4(new_n754), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n767), .B1(new_n860), .B2(new_n693), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n774), .A2(new_n775), .A3(new_n768), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT109), .B1(new_n862), .B2(new_n757), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n776), .A2(new_n777), .A3(new_n770), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n704), .B1(new_n626), .B2(new_n643), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n647), .A2(new_n654), .B1(new_n729), .B2(new_n737), .ZN(new_n867));
  INV_X1    g681(.A(new_n408), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n619), .B2(new_n692), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n631), .A2(new_n638), .A3(new_n632), .A4(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n607), .A2(new_n867), .A3(new_n712), .A4(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n742), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n757), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n653), .B1(new_n780), .B2(new_n765), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n416), .A2(new_n640), .A3(new_n639), .A4(new_n667), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n303), .A3(new_n187), .A4(new_n304), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n787), .A2(new_n874), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n865), .A2(new_n872), .A3(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n742), .A2(new_n743), .ZN(new_n883));
  INV_X1    g697(.A(new_n751), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n735), .A2(new_n652), .A3(new_n666), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n678), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n672), .A2(new_n695), .A3(new_n883), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT52), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n744), .B1(new_n875), .B2(new_n671), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT52), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n695), .A4(new_n886), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n859), .B1(new_n882), .B2(new_n892), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n607), .A2(new_n867), .A3(new_n712), .A4(new_n870), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n757), .A2(new_n873), .B1(new_n875), .B2(new_n879), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n781), .B(new_n703), .C1(new_n625), .C2(new_n642), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n787), .A4(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n784), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n888), .A2(new_n891), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(KEYINPUT53), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n893), .A2(new_n900), .A3(KEYINPUT54), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n858), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n829), .B1(new_n905), .B2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n224), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n297), .B1(new_n893), .B2(new_n900), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT56), .B1(new_n910), .B2(G210), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n274), .A2(new_n271), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n228), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n909), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n911), .A2(new_n914), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n911), .A2(KEYINPUT119), .A3(new_n914), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G51));
  XOR2_X1   g734(.A(new_n476), .B(KEYINPUT57), .Z(new_n921));
  NAND3_X1  g735(.A1(new_n903), .A2(new_n904), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n474), .B2(new_n472), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n910), .B(new_n791), .C1(new_n790), .C2(new_n789), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n908), .B1(new_n923), .B2(new_n924), .ZN(G54));
  NAND3_X1  g739(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n926), .A2(new_n351), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n351), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n927), .A2(new_n928), .A3(new_n908), .ZN(G60));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT59), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n903), .A2(new_n904), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n613), .A3(new_n612), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n903), .A2(new_n614), .A3(new_n904), .A4(new_n931), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n933), .A2(new_n909), .A3(new_n934), .ZN(G63));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT61), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n909), .B1(new_n936), .B2(KEYINPUT61), .ZN(new_n938));
  XNOR2_X1  g752(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n368), .A2(new_n297), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT53), .B1(new_n898), .B2(new_n899), .ZN(new_n942));
  NOR4_X1   g756(.A1(new_n892), .A2(new_n897), .A3(new_n784), .A4(new_n859), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n938), .B1(new_n944), .B2(new_n513), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n946));
  AND4_X1   g760(.A1(new_n946), .A2(new_n901), .A3(new_n650), .A4(new_n941), .ZN(new_n947));
  INV_X1    g761(.A(new_n941), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n893), .B2(new_n900), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n949), .B2(new_n650), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n937), .B(new_n945), .C1(new_n947), .C2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n650), .B(new_n941), .C1(new_n942), .C2(new_n943), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT121), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n949), .A2(new_n946), .A3(new_n650), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n937), .B1(new_n956), .B2(new_n945), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n952), .A2(new_n957), .ZN(G66));
  INV_X1    g772(.A(G224), .ZN(new_n959));
  OAI21_X1  g773(.A(G953), .B1(new_n412), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n872), .B2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n912), .B1(G898), .B2(new_n224), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  OAI21_X1  g777(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n312), .A2(new_n313), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n869), .A2(new_n756), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n781), .A2(new_n632), .A3(new_n685), .A4(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT125), .B1(new_n809), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT125), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n971), .B(new_n968), .C1(new_n798), .C2(new_n808), .ZN(new_n972));
  AOI22_X1  g786(.A1(new_n817), .A2(new_n820), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n672), .A2(new_n695), .A3(new_n883), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT123), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n689), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n974), .B1(new_n978), .B2(KEYINPUT62), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT62), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n977), .A2(KEYINPUT124), .A3(new_n980), .A4(new_n689), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n973), .A2(new_n979), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n966), .B1(new_n983), .B2(new_n224), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n966), .B1(new_n662), .B2(new_n224), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n975), .B(KEYINPUT123), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n766), .A2(new_n680), .A3(new_n683), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT126), .B1(new_n798), .B2(new_n987), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n798), .A2(new_n987), .A3(KEYINPUT126), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n787), .B1(new_n798), .B2(new_n808), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n991), .A2(new_n784), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n821), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n985), .B1(new_n993), .B2(new_n224), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n224), .B1(G227), .B2(G900), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT127), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  OR3_X1    g811(.A1(new_n984), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n997), .B1(new_n984), .B2(new_n994), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(G72));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  NAND3_X1  g816(.A1(new_n821), .A2(new_n990), .A3(new_n992), .ZN(new_n1003));
  INV_X1    g817(.A(new_n872), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1005), .A2(new_n526), .A3(new_n547), .A4(new_n562), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n592), .A2(new_n563), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n901), .A2(new_n1002), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1006), .A2(new_n909), .A3(new_n1008), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n983), .A2(new_n1004), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n674), .B1(new_n1010), .B2(new_n1002), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1009), .A2(new_n1011), .ZN(G57));
endmodule


