//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NOR3_X1   g009(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  OAI22_X1  g012(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(KEYINPUT15), .A3(new_n215), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n215), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(KEYINPUT15), .B2(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT94), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n211), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n211), .A2(new_n219), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n210), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n216), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n208), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(KEYINPUT17), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(new_n207), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n227), .B(KEYINPUT95), .Z(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT18), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n207), .B(new_n223), .Z(new_n231));
  XNOR2_X1  g030(.A(new_n228), .B(KEYINPUT13), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n226), .A2(KEYINPUT18), .A3(new_n229), .ZN(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G141gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G169gat), .B(G197gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n233), .A2(new_n234), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n241), .B1(new_n233), .B2(new_n234), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT96), .ZN(new_n246));
  INV_X1    g045(.A(new_n244), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n247), .A2(KEYINPUT96), .A3(new_n242), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT92), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT31), .B(G50gat), .ZN(new_n252));
  INV_X1    g051(.A(G106gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G228gat), .A2(G233gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT84), .Z(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G141gat), .B(G148gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT2), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(G155gat), .B2(G162gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G141gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G148gat), .ZN(new_n267));
  INV_X1    g066(.A(G148gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G141gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G155gat), .B(G162gat), .ZN(new_n271));
  INV_X1    g070(.A(G155gat), .ZN(new_n272));
  INV_X1    g071(.A(G162gat), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT2), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n270), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n265), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G197gat), .B(G204gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT22), .ZN(new_n278));
  INV_X1    g077(.A(G211gat), .ZN(new_n279));
  INV_X1    g078(.A(G218gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G211gat), .B(G218gat), .Z(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT85), .ZN(new_n285));
  INV_X1    g084(.A(new_n282), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT79), .ZN(new_n287));
  INV_X1    g086(.A(new_n283), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT79), .B1(new_n282), .B2(new_n283), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT29), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n276), .B1(new_n292), .B2(KEYINPUT3), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n282), .A2(KEYINPUT78), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n282), .A2(KEYINPUT78), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n283), .A3(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT3), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n265), .A2(new_n275), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n258), .B1(new_n293), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT29), .B1(new_n291), .B2(new_n296), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n276), .B1(new_n304), .B2(KEYINPUT3), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n301), .A2(KEYINPUT86), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(KEYINPUT86), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n297), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n256), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n305), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(G22gat), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n265), .A2(new_n275), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n289), .A2(new_n290), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT85), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n284), .B(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n300), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n312), .B1(new_n316), .B2(new_n298), .ZN(new_n317));
  INV_X1    g116(.A(new_n302), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n257), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G22gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n308), .A3(new_n309), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G78gat), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n311), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n311), .B2(new_n322), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n255), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n322), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G78gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n322), .A3(new_n323), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n329), .A3(new_n254), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G1gat), .B(G29gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT0), .ZN(new_n333));
  XNOR2_X1  g132(.A(G57gat), .B(G85gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n337));
  INV_X1    g136(.A(G120gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G113gat), .ZN(new_n339));
  INV_X1    g138(.A(G113gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G120gat), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n337), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n341), .A3(new_n337), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G127gat), .B(G134gat), .Z(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(KEYINPUT1), .ZN(new_n348));
  OR3_X1    g147(.A1(new_n340), .A2(KEYINPUT74), .A3(G120gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n339), .A2(KEYINPUT74), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n341), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n346), .A2(new_n347), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n312), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n345), .A2(new_n344), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n347), .B1(new_n355), .B2(new_n342), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n348), .A2(new_n351), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n358), .A2(new_n299), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n312), .A2(new_n356), .A3(new_n357), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT4), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n354), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n365), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n358), .A2(new_n276), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n361), .ZN(new_n369));
  INV_X1    g168(.A(new_n365), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n364), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n366), .A2(KEYINPUT83), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n361), .A2(KEYINPUT4), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n353), .B1(new_n352), .B2(new_n312), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n299), .A3(new_n359), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(KEYINPUT83), .B(new_n371), .C1(new_n376), .C2(new_n370), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n336), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT90), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n359), .A2(new_n299), .ZN(new_n383));
  OAI211_X1 g182(.A(KEYINPUT4), .B(new_n361), .C1(new_n383), .C2(new_n352), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n370), .B1(new_n384), .B2(new_n354), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n382), .B1(new_n385), .B2(new_n364), .ZN(new_n386));
  INV_X1    g185(.A(new_n361), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n312), .B1(new_n356), .B2(new_n357), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n370), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT5), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n335), .B(new_n377), .C1(new_n386), .C2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n377), .B1(new_n386), .B2(new_n391), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(KEYINPUT90), .A3(new_n336), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(KEYINPUT6), .A3(new_n336), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT68), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n400));
  INV_X1    g199(.A(G169gat), .ZN(new_n401));
  INV_X1    g200(.A(G176gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT23), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT23), .ZN(new_n407));
  NAND2_X1  g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(G183gat), .A2(G190gat), .ZN(new_n410));
  AND2_X1   g209(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(new_n411), .B2(G190gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(G183gat), .A2(G190gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT24), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n413), .A2(KEYINPUT65), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT65), .B1(new_n413), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n409), .B1(new_n417), .B2(KEYINPUT66), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT66), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n412), .B(new_n419), .C1(new_n415), .C2(new_n416), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n400), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n413), .A2(new_n414), .ZN(new_n423));
  NAND3_X1  g222(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT67), .B(G190gat), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n423), .B(new_n424), .C1(new_n425), .C2(G183gat), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n422), .A2(new_n426), .A3(KEYINPUT25), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n399), .B1(new_n421), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n429));
  AND2_X1   g228(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT27), .B(G183gat), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n429), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G183gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT27), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G183gat), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n436), .A2(new_n438), .A3(KEYINPUT70), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT70), .B1(new_n436), .B2(new_n438), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT28), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n425), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n434), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n406), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n403), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n445), .A2(KEYINPUT71), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT71), .B1(new_n445), .B2(new_n447), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT72), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n434), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n438), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT70), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n433), .A2(KEYINPUT70), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n443), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n449), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT71), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT72), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n451), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n400), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n424), .B1(G183gat), .B2(G190gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT65), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n423), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n413), .A2(KEYINPUT65), .A3(new_n414), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n422), .B1(new_n470), .B2(new_n419), .ZN(new_n471));
  INV_X1    g270(.A(new_n420), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n427), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(KEYINPUT68), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(G226gat), .A2(G233gat), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n428), .A2(new_n464), .A3(new_n475), .A4(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(KEYINPUT29), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n417), .A2(KEYINPUT66), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(new_n420), .A3(new_n422), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n427), .B1(new_n481), .B2(new_n465), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n444), .A2(new_n450), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n297), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT80), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n482), .A2(new_n476), .A3(new_n483), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n428), .A2(new_n464), .A3(new_n475), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(new_n479), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n297), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT80), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n485), .A2(new_n493), .A3(new_n486), .ZN(new_n494));
  XOR2_X1   g293(.A(G8gat), .B(G36gat), .Z(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT81), .ZN(new_n496));
  XNOR2_X1  g295(.A(G64gat), .B(G92gat), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n496), .B(new_n497), .Z(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n488), .A2(new_n492), .A3(new_n494), .A4(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n488), .A2(new_n501), .A3(new_n492), .A4(new_n494), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n491), .B2(new_n486), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n297), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n502), .A2(new_n507), .A3(new_n498), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n397), .A2(new_n398), .A3(new_n500), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n493), .B1(new_n485), .B2(new_n486), .ZN(new_n510));
  AOI211_X1 g309(.A(KEYINPUT80), .B(new_n297), .C1(new_n478), .C2(new_n484), .ZN(new_n511));
  AOI211_X1 g310(.A(new_n486), .B(new_n489), .C1(new_n490), .C2(new_n479), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n499), .B1(new_n513), .B2(new_n501), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n511), .A2(new_n512), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n488), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT37), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n503), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n331), .B1(new_n509), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT88), .B1(new_n363), .B2(new_n365), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n376), .A2(new_n521), .A3(new_n370), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT39), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n368), .A2(new_n365), .A3(new_n361), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT39), .B1(new_n526), .B2(KEYINPUT89), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n527), .B1(KEYINPUT89), .B2(new_n526), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(new_n520), .A3(new_n522), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n529), .A3(new_n335), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT40), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n525), .A2(new_n529), .A3(KEYINPUT40), .A4(new_n335), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n532), .A2(new_n381), .A3(new_n396), .A4(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT82), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n500), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n513), .A2(new_n499), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n500), .A2(new_n536), .A3(new_n535), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n534), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n251), .B1(new_n519), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n398), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n395), .A2(KEYINPUT90), .A3(new_n336), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT90), .B1(new_n395), .B2(new_n336), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n543), .B1(new_n546), .B2(new_n394), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n502), .A2(new_n498), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n501), .B1(new_n515), .B2(new_n488), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n504), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n547), .A2(new_n500), .A3(new_n550), .A4(new_n508), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n500), .A2(new_n536), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT30), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n516), .A2(new_n498), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n540), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n534), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n551), .A2(new_n557), .A3(KEYINPUT92), .A4(new_n331), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n326), .A2(new_n330), .ZN(new_n560));
  INV_X1    g359(.A(new_n379), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n392), .A2(new_n393), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n398), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n560), .B1(new_n555), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT77), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(KEYINPUT77), .A2(KEYINPUT36), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n490), .A2(new_n352), .ZN(new_n570));
  INV_X1    g369(.A(G227gat), .ZN(new_n571));
  INV_X1    g370(.A(G233gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n428), .A2(new_n464), .A3(new_n475), .A4(new_n358), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G15gat), .B(G43gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT75), .ZN(new_n577));
  XNOR2_X1  g376(.A(G71gat), .B(G99gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT33), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT76), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n575), .A2(KEYINPUT76), .A3(KEYINPUT32), .A4(new_n580), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n573), .B1(new_n570), .B2(new_n574), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT34), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n575), .A2(KEYINPUT32), .ZN(new_n588));
  INV_X1    g387(.A(new_n575), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n588), .B(new_n579), .C1(new_n589), .C2(KEYINPUT33), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n585), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n587), .B1(new_n585), .B2(new_n590), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n568), .B(new_n569), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n585), .A2(new_n590), .ZN(new_n594));
  INV_X1    g393(.A(new_n587), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n585), .A2(new_n587), .A3(new_n590), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n596), .A2(new_n566), .A3(new_n567), .A4(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n565), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT87), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n565), .A2(new_n593), .A3(new_n598), .A4(KEYINPUT87), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n559), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n591), .A2(new_n592), .ZN(new_n604));
  INV_X1    g403(.A(new_n540), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n605), .A2(new_n537), .A3(new_n538), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n604), .A2(new_n606), .A3(new_n563), .A4(new_n331), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n596), .A2(new_n597), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(new_n560), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT35), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n544), .A2(new_n545), .A3(new_n562), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n610), .B1(new_n611), .B2(new_n543), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(new_n555), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n607), .A2(KEYINPUT35), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n250), .B1(new_n603), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G64gat), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT97), .B1(new_n617), .B2(G57gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n619));
  INV_X1    g418(.A(G57gat), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(G64gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(G57gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT98), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n618), .A2(new_n621), .A3(new_n625), .A4(new_n622), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT9), .ZN(new_n629));
  NAND2_X1  g428(.A1(G71gat), .A2(G78gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n620), .A2(G64gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n622), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT9), .ZN(new_n635));
  INV_X1    g434(.A(new_n628), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n632), .A2(KEYINPUT99), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n624), .A2(new_n626), .B1(new_n630), .B2(new_n629), .ZN(new_n640));
  INV_X1    g439(.A(new_n637), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT100), .B(KEYINPUT21), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G231gat), .A2(G233gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G127gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G183gat), .B(G211gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n638), .A2(new_n642), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n208), .B1(new_n650), .B2(KEYINPUT21), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT102), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT101), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n272), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n652), .B(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n649), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT7), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(KEYINPUT103), .A2(KEYINPUT7), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n662), .A2(G85gat), .A3(G92gat), .A4(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(G85gat), .ZN(new_n665));
  INV_X1    g464(.A(G92gat), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n660), .B(new_n661), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(G99gat), .A2(G106gat), .ZN(new_n668));
  AOI22_X1  g467(.A1(KEYINPUT8), .A2(new_n668), .B1(new_n665), .B2(new_n666), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(G99gat), .B(G106gat), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n671), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(KEYINPUT104), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677));
  INV_X1    g476(.A(new_n675), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n674), .A2(new_n671), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n225), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n676), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n223), .ZN(new_n683));
  NAND3_X1  g482(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(G190gat), .B(G218gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(G134gat), .B(G162gat), .Z(new_n688));
  AOI21_X1  g487(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  OR3_X1    g489(.A1(new_n687), .A2(KEYINPUT105), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n690), .B(KEYINPUT105), .Z(new_n692));
  NAND2_X1  g491(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n659), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT10), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n680), .B2(new_n676), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n650), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n638), .A2(new_n642), .B1(new_n673), .B2(new_n675), .ZN(new_n701));
  AOI211_X1 g500(.A(new_n679), .B(new_n678), .C1(new_n632), .C2(new_n637), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n696), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n697), .A2(KEYINPUT106), .A3(new_n650), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(G230gat), .A2(G233gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OR3_X1    g506(.A1(new_n701), .A2(new_n702), .A3(new_n706), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(G120gat), .B(G148gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT107), .ZN(new_n711));
  XOR2_X1   g510(.A(G176gat), .B(G204gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n709), .A2(new_n713), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n695), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n616), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n564), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g520(.A1(new_n616), .A2(new_n555), .A3(new_n717), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n203), .A2(new_n206), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(KEYINPUT42), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT108), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n725), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n722), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1325gat));
  AOI21_X1  g528(.A(G15gat), .B1(new_n719), .B2(new_n604), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT109), .Z(new_n731));
  NAND2_X1  g530(.A1(new_n593), .A2(new_n598), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n719), .A2(G15gat), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT110), .ZN(G1326gat));
  NOR2_X1   g534(.A1(new_n718), .A2(new_n331), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT43), .B(G22gat), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1327gat));
  NOR3_X1   g537(.A1(new_n659), .A2(new_n694), .A3(new_n716), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n616), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n740), .A2(G29gat), .A3(new_n563), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT45), .Z(new_n742));
  NAND2_X1  g541(.A1(new_n603), .A2(new_n615), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n694), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n599), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n614), .B1(new_n559), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n744), .B1(new_n748), .B2(new_n694), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n659), .A2(new_n245), .A3(new_n716), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n746), .A2(new_n749), .A3(KEYINPUT111), .A4(new_n750), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n753), .A2(new_n564), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n742), .B1(new_n212), .B2(new_n755), .ZN(G1328gat));
  NOR3_X1   g555(.A1(new_n740), .A2(G36gat), .A3(new_n606), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT46), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n753), .A2(new_n555), .A3(new_n754), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n213), .B2(new_n759), .ZN(G1329gat));
  NOR3_X1   g559(.A1(new_n740), .A2(G43gat), .A3(new_n608), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n732), .ZN(new_n763));
  OAI21_X1  g562(.A(G43gat), .B1(new_n751), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n764), .A3(KEYINPUT47), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n753), .A2(new_n732), .A3(new_n754), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G43gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n762), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n761), .B1(new_n767), .B2(G43gat), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n772), .A2(KEYINPUT112), .A3(KEYINPUT47), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n765), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(KEYINPUT113), .B(new_n765), .C1(new_n771), .C2(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(G1330gat));
  NOR3_X1   g577(.A1(new_n740), .A2(G50gat), .A3(new_n331), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(G50gat), .B1(new_n751), .B2(new_n331), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n753), .A2(new_n560), .A3(new_n754), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n779), .B1(new_n784), .B2(G50gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n785), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g585(.A(new_n748), .ZN(new_n787));
  INV_X1    g586(.A(new_n245), .ZN(new_n788));
  INV_X1    g587(.A(new_n716), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n695), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n564), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n555), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n796));
  XOR2_X1   g595(.A(KEYINPUT49), .B(G64gat), .Z(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n795), .B2(new_n797), .ZN(G1333gat));
  OAI21_X1  g597(.A(G71gat), .B1(new_n791), .B2(new_n763), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n608), .A2(G71gat), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n791), .B2(new_n800), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g601(.A1(new_n792), .A2(new_n560), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g603(.A1(new_n746), .A2(new_n749), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n659), .A2(new_n788), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n716), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n805), .A2(KEYINPUT115), .A3(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(G85gat), .B1(new_n813), .B2(new_n563), .ZN(new_n814));
  INV_X1    g613(.A(new_n694), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n787), .A2(new_n815), .A3(new_n806), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n816), .A2(KEYINPUT51), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n789), .B1(new_n816), .B2(KEYINPUT51), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n665), .A3(new_n564), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n814), .A2(new_n821), .ZN(G1336gat));
  OAI21_X1  g621(.A(G92gat), .B1(new_n809), .B2(new_n606), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n555), .A2(new_n666), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n823), .B(new_n824), .C1(new_n819), .C2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n819), .A2(new_n825), .ZN(new_n827));
  INV_X1    g626(.A(new_n813), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n555), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n827), .B1(new_n829), .B2(G92gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n826), .B1(new_n830), .B2(new_n824), .ZN(G1337gat));
  AOI21_X1  g630(.A(G99gat), .B1(new_n820), .B2(new_n604), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n732), .A2(G99gat), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n828), .B2(new_n833), .ZN(G1338gat));
  NAND3_X1  g633(.A1(new_n811), .A2(new_n560), .A3(new_n812), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G106gat), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT116), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n838), .A3(G106gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n820), .A2(new_n253), .A3(new_n560), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n843), .ZN(new_n845));
  OAI21_X1  g644(.A(G106gat), .B1(new_n809), .B2(new_n331), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  OAI22_X1  g646(.A1(new_n841), .A2(new_n842), .B1(new_n844), .B2(new_n847), .ZN(G1339gat));
  NAND2_X1  g647(.A1(new_n717), .A2(new_n245), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT118), .B1(new_n705), .B2(new_n706), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n697), .A2(new_n650), .A3(KEYINPUT106), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT106), .B1(new_n697), .B2(new_n650), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  INV_X1    g653(.A(new_n706), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n703), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n850), .A2(new_n856), .A3(KEYINPUT54), .A4(new_n707), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n855), .B1(new_n853), .B2(new_n703), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n713), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n857), .A2(new_n860), .A3(KEYINPUT55), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(new_n715), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n857), .A2(new_n860), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT55), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT119), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n866), .B(KEYINPUT55), .C1(new_n857), .C2(new_n860), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n862), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n862), .B(KEYINPUT120), .C1(new_n865), .C2(new_n867), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n788), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n226), .A2(new_n229), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n231), .A2(new_n232), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n239), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n242), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n716), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n815), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n815), .A2(new_n876), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n870), .A2(new_n879), .A3(new_n871), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT121), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n659), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n878), .A2(KEYINPUT121), .A3(new_n880), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n849), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n609), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n555), .A2(new_n563), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(new_n340), .A3(new_n250), .ZN(new_n889));
  INV_X1    g688(.A(new_n888), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n788), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n340), .B2(new_n891), .ZN(G1340gat));
  NOR2_X1   g691(.A1(new_n888), .A2(new_n789), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(new_n338), .ZN(G1341gat));
  NAND2_X1  g693(.A1(new_n890), .A2(new_n659), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g695(.A1(new_n815), .A2(new_n606), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(G134gat), .A3(new_n563), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n886), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT56), .Z(new_n900));
  OAI21_X1  g699(.A(G134gat), .B1(new_n888), .B2(new_n694), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1343gat));
  NAND2_X1  g701(.A1(new_n763), .A2(new_n887), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n885), .B2(new_n560), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n560), .A2(KEYINPUT57), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n877), .B(KEYINPUT122), .Z(new_n907));
  NAND2_X1  g706(.A1(new_n863), .A2(new_n864), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n249), .A2(new_n862), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n815), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n882), .B1(new_n910), .B2(new_n880), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n906), .B1(new_n911), .B2(new_n849), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n904), .B1(new_n905), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(G141gat), .B1(new_n913), .B2(new_n250), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n250), .A2(G141gat), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n885), .A2(new_n560), .A3(new_n904), .A4(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n788), .B(new_n904), .C1(new_n905), .C2(new_n912), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G141gat), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n917), .B(KEYINPUT123), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n919), .B1(new_n923), .B2(KEYINPUT58), .ZN(new_n924));
  AOI211_X1 g723(.A(KEYINPUT124), .B(new_n915), .C1(new_n921), .C2(new_n922), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n918), .B1(new_n924), .B2(new_n925), .ZN(G1344gat));
  NAND2_X1  g725(.A1(new_n885), .A2(new_n560), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n903), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n268), .A3(new_n716), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n878), .A2(new_n880), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n882), .A3(new_n881), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n906), .B1(new_n934), .B2(new_n849), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n879), .B(new_n862), .C1(new_n865), .C2(new_n867), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n882), .B1(new_n910), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n250), .A2(new_n717), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT57), .B1(new_n940), .B2(new_n560), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n904), .A2(new_n716), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n268), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT125), .B1(new_n942), .B2(new_n943), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n930), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n913), .A2(new_n789), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n949), .A2(KEYINPUT59), .A3(new_n268), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n929), .B1(new_n948), .B2(new_n950), .ZN(G1345gat));
  OAI21_X1  g750(.A(G155gat), .B1(new_n913), .B2(new_n882), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n928), .A2(new_n272), .A3(new_n659), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1346gat));
  OAI21_X1  g753(.A(G162gat), .B1(new_n913), .B2(new_n694), .ZN(new_n955));
  OR4_X1    g754(.A1(G162gat), .A2(new_n732), .A3(new_n563), .A4(new_n897), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n927), .B2(new_n956), .ZN(G1347gat));
  NOR2_X1   g756(.A1(new_n606), .A2(new_n564), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n886), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(G169gat), .B1(new_n959), .B2(new_n788), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n886), .A2(new_n958), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n961), .A2(new_n401), .A3(new_n250), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n960), .A2(new_n962), .ZN(G1348gat));
  NOR2_X1   g762(.A1(new_n961), .A2(new_n789), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(new_n402), .ZN(G1349gat));
  OAI21_X1  g764(.A(new_n435), .B1(new_n961), .B2(new_n882), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n959), .A2(new_n659), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n441), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT60), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n968), .B(new_n969), .ZN(G1350gat));
  NAND2_X1  g769(.A1(new_n959), .A2(new_n815), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n971), .A2(new_n425), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(G190gat), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n975), .B1(new_n973), .B2(new_n974), .ZN(G1351gat));
  AND4_X1   g775(.A1(new_n560), .A2(new_n885), .A3(new_n763), .A4(new_n958), .ZN(new_n977));
  AOI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n788), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n763), .A2(new_n958), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n942), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n249), .A2(G197gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(G1352gat));
  INV_X1    g781(.A(G204gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n977), .A2(new_n983), .A3(new_n716), .ZN(new_n984));
  XOR2_X1   g783(.A(new_n984), .B(KEYINPUT62), .Z(new_n985));
  NAND2_X1  g784(.A1(new_n980), .A2(new_n716), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n985), .B1(new_n987), .B2(new_n983), .ZN(G1353gat));
  NAND3_X1  g787(.A1(new_n977), .A2(new_n279), .A3(new_n659), .ZN(new_n989));
  INV_X1    g788(.A(new_n979), .ZN(new_n990));
  OAI211_X1 g789(.A(new_n659), .B(new_n990), .C1(new_n935), .C2(new_n941), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(G211gat), .B1(new_n991), .B2(new_n992), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n995), .A2(KEYINPUT63), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT63), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n993), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n989), .B1(new_n996), .B2(new_n998), .ZN(G1354gat));
  NAND3_X1  g798(.A1(new_n977), .A2(new_n280), .A3(new_n815), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n1001));
  INV_X1    g800(.A(new_n1001), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n1003));
  NOR3_X1   g802(.A1(new_n1002), .A2(new_n694), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1000), .B1(new_n1004), .B2(new_n280), .ZN(G1355gat));
endmodule


