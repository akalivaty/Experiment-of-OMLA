//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n562, new_n563, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT67), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n461), .A2(new_n463), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n464), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT66), .ZN(new_n478));
  OAI21_X1  g053(.A(G2105), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n469), .A2(new_n465), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n470), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(new_n464), .A2(G126), .ZN(new_n489));
  OR2_X1    g064(.A1(KEYINPUT68), .A2(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT68), .A2(G114), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(G2104), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n465), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI22_X1  g070(.A1(new_n493), .A2(new_n494), .B1(new_n495), .B2(new_n466), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n469), .A2(new_n494), .A3(new_n495), .ZN(new_n497));
  AND2_X1   g072(.A1(G102), .A2(G2104), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n465), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n507), .B2(KEYINPUT6), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT69), .B(G651), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n508), .A2(G50), .B1(G75), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n509), .A2(new_n513), .A3(G62), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  INV_X1    g090(.A(new_n503), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n516), .B(new_n513), .C1(new_n509), .C2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n521), .A2(KEYINPUT70), .A3(new_n516), .A4(new_n513), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n512), .B(new_n514), .C1(new_n515), .C2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND3_X1  g100(.A1(new_n520), .A2(new_n522), .A3(G89), .ZN(new_n526));
  OAI211_X1 g101(.A(G543), .B(new_n516), .C1(new_n509), .C2(new_n517), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n526), .A2(new_n529), .A3(new_n531), .A4(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT5), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G543), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n537), .A3(G64), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT71), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n538), .A2(new_n542), .A3(new_n539), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n541), .A2(new_n509), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n520), .A2(new_n522), .A3(G90), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n528), .A2(G52), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n541), .A2(KEYINPUT72), .A3(new_n509), .A4(new_n543), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND3_X1  g126(.A1(new_n520), .A2(new_n522), .A3(G81), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n507), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n528), .A2(G43), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT73), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G188));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n520), .A2(new_n522), .A3(G91), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n567), .B(new_n568), .C1(new_n527), .C2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n502), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n566), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n567), .B1(new_n527), .B2(new_n569), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n508), .A2(KEYINPUT74), .A3(G53), .A4(G543), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT9), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n565), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n566), .A2(new_n570), .A3(new_n572), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n574), .A2(KEYINPUT9), .A3(new_n575), .ZN(new_n579));
  NOR3_X1   g154(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT75), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(G299));
  OAI21_X1  g156(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n528), .A2(G49), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n582), .B(new_n583), .C1(new_n523), .C2(new_n584), .ZN(G288));
  NAND3_X1  g160(.A1(new_n520), .A2(new_n522), .A3(G86), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n528), .A2(G48), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(new_n507), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n528), .A2(G47), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n591), .B1(new_n507), .B2(new_n592), .C1(new_n523), .C2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT76), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  XOR2_X1   g172(.A(KEYINPUT77), .B(KEYINPUT10), .Z(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n523), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n535), .A2(new_n537), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n528), .A2(G54), .B1(G651), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n520), .A2(new_n522), .A3(G92), .A4(new_n598), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n601), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n597), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n597), .B1(new_n609), .B2(G868), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n609), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g196(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n482), .A2(G123), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n470), .A2(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(new_n465), .B2(G111), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n626), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2430), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT78), .B(KEYINPUT14), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT79), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT80), .Z(new_n649));
  INV_X1    g224(.A(G14), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n645), .B2(new_n647), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XNOR2_X1  g228(.A(G2072), .B(G2078), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT81), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  INV_X1    g235(.A(new_n656), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(new_n657), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(KEYINPUT17), .A3(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n664));
  OAI221_X1 g239(.A(new_n663), .B1(new_n661), .B2(new_n657), .C1(new_n664), .C2(new_n655), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n632), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n625), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n673), .A2(new_n675), .A3(new_n677), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n680), .B(new_n681), .C1(new_n679), .C2(new_n678), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(G1986), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT22), .B(G1981), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(G229));
  NOR2_X1   g265(.A1(G16), .A2(G22), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G166), .B2(G16), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT86), .B(G1971), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G6), .ZN(new_n696));
  AND3_X1   g271(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(G16), .A2(G23), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G288), .B2(new_n695), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT33), .ZN(new_n703));
  INV_X1    g278(.A(G1976), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n694), .B(new_n700), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(KEYINPUT87), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n707), .A2(new_n711), .A3(KEYINPUT34), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n708), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n595), .A2(G16), .ZN(new_n714));
  OR2_X1    g289(.A1(G16), .A2(G24), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT85), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1986), .ZN(new_n718));
  OR2_X1    g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n719), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT82), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n482), .A2(G119), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n470), .A2(G131), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n721), .A2(KEYINPUT83), .A3(new_n722), .A4(new_n723), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G25), .B(new_n728), .S(G29), .Z(new_n729));
  XOR2_X1   g304(.A(KEYINPUT35), .B(G1991), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT84), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n729), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n713), .A2(new_n718), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT88), .B(KEYINPUT36), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI22_X1  g311(.A1(G129), .A2(new_n482), .B1(new_n470), .B2(G141), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT26), .Z(new_n740));
  NAND3_X1  g315(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G32), .B(new_n741), .S(G29), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT27), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1996), .ZN(new_n744));
  INV_X1    g319(.A(new_n735), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n713), .A2(new_n745), .A3(new_n718), .A4(new_n733), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n695), .A2(G4), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n609), .B2(new_n695), .ZN(new_n748));
  INV_X1    g323(.A(G1348), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n695), .A2(G19), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n557), .B2(new_n695), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT89), .B(G1341), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G29), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(G26), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n482), .A2(G128), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n470), .A2(G140), .ZN(new_n758));
  NOR2_X1   g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n756), .B1(new_n761), .B2(G29), .ZN(new_n762));
  MUX2_X1   g337(.A(new_n756), .B(new_n762), .S(KEYINPUT28), .Z(new_n763));
  XOR2_X1   g338(.A(KEYINPUT90), .B(G2067), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n750), .A2(new_n754), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT91), .ZN(new_n767));
  AND2_X1   g342(.A1(KEYINPUT24), .A2(G34), .ZN(new_n768));
  NOR2_X1   g343(.A1(KEYINPUT24), .A2(G34), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n755), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n480), .B2(new_n755), .ZN(new_n771));
  INV_X1    g346(.A(G2084), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT92), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n695), .A2(G5), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G171), .B2(new_n695), .ZN(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n755), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n755), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT95), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n780), .B(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n774), .B(new_n778), .C1(G2090), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n755), .A2(G27), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G164), .B2(new_n755), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(G2078), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n787), .A2(G2078), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n788), .B(new_n789), .C1(new_n772), .C2(new_n771), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT31), .B(G11), .Z(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT30), .B(G28), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n755), .B2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G1966), .ZN(new_n794));
  NAND2_X1  g369(.A1(G168), .A2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G16), .B2(G21), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n790), .B(new_n793), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n794), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT93), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n785), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(G299), .A2(G16), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n695), .A2(KEYINPUT23), .A3(G20), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT23), .ZN(new_n803));
  INV_X1    g378(.A(G20), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G16), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(G1956), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n784), .A2(G2090), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n807), .A2(KEYINPUT96), .A3(new_n808), .ZN(new_n812));
  AND4_X1   g387(.A1(new_n767), .A2(new_n800), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n736), .A2(new_n744), .A3(new_n746), .A4(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(G29), .A2(G33), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT25), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n470), .A2(G139), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n465), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n815), .B1(new_n820), .B2(new_n755), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(G2072), .Z(new_n822));
  NOR2_X1   g397(.A1(new_n631), .A2(new_n755), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n814), .A2(new_n822), .A3(new_n823), .ZN(G311));
  AND3_X1   g399(.A1(new_n736), .A2(new_n746), .A3(new_n813), .ZN(new_n825));
  INV_X1    g400(.A(new_n822), .ZN(new_n826));
  INV_X1    g401(.A(new_n823), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n825), .A2(new_n826), .A3(new_n827), .A4(new_n744), .ZN(G150));
  XOR2_X1   g403(.A(KEYINPUT97), .B(G55), .Z(new_n829));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  INV_X1    g405(.A(G67), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n603), .B2(new_n831), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n528), .A2(new_n829), .B1(new_n509), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n520), .A2(new_n522), .A3(G93), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND4_X1  g412(.A1(new_n835), .A2(new_n554), .A3(new_n552), .A4(new_n555), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n556), .A2(new_n834), .A3(new_n833), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n609), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n837), .B1(new_n844), .B2(G860), .ZN(G145));
  XNOR2_X1  g420(.A(new_n480), .B(new_n631), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n500), .B(new_n761), .Z(new_n848));
  XOR2_X1   g423(.A(new_n741), .B(new_n820), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n623), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n852));
  INV_X1    g427(.A(G142), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n466), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n482), .A2(G130), .ZN(new_n855));
  OR2_X1    g430(.A1(G106), .A2(G2105), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n470), .A2(KEYINPUT98), .A3(G142), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n854), .A2(new_n855), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n728), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n726), .A2(new_n727), .A3(new_n859), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n851), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n864), .A3(new_n623), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT100), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n867), .A2(new_n869), .A3(KEYINPUT100), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n850), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n850), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n873), .A2(new_n875), .A3(G162), .ZN(new_n876));
  INV_X1    g451(.A(new_n850), .ZN(new_n877));
  INV_X1    g452(.A(new_n872), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(new_n870), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n487), .B1(new_n879), .B2(new_n874), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n847), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  OAI21_X1  g457(.A(G162), .B1(new_n873), .B2(new_n875), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n879), .A2(new_n487), .A3(new_n874), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n846), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g462(.A1(new_n835), .A2(new_n612), .ZN(new_n888));
  XNOR2_X1  g463(.A(G303), .B(G288), .ZN(new_n889));
  NAND2_X1  g464(.A1(G290), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G288), .ZN(new_n891));
  XNOR2_X1  g466(.A(G303), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n595), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(G305), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n896), .A2(KEYINPUT102), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(KEYINPUT102), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n890), .A2(new_n893), .A3(new_n697), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n895), .A2(new_n897), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n895), .A2(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n900), .B1(new_n902), .B2(new_n898), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT101), .B1(new_n577), .B2(new_n580), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n573), .A2(new_n565), .A3(new_n576), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT75), .B1(new_n578), .B2(new_n579), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n609), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(G299), .A2(new_n907), .A3(new_n608), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n840), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(new_n618), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n909), .A2(KEYINPUT41), .A3(new_n910), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT41), .B1(new_n909), .B2(new_n910), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n914), .B1(new_n917), .B2(new_n913), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n903), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n888), .B1(new_n919), .B2(new_n612), .ZN(G331));
  NAND2_X1  g495(.A1(G331), .A2(KEYINPUT103), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n922), .B(new_n888), .C1(new_n919), .C2(new_n612), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(G295));
  AND2_X1   g499(.A1(new_n546), .A2(new_n549), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n547), .A2(new_n548), .ZN(new_n926));
  AOI21_X1  g501(.A(G286), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(G168), .A2(G301), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n840), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n925), .A2(G286), .A3(new_n926), .ZN(new_n931));
  NAND2_X1  g506(.A1(G168), .A2(G301), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n839), .A4(new_n838), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n912), .A2(KEYINPUT104), .A3(new_n932), .A4(new_n931), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT106), .B1(new_n936), .B2(new_n911), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT41), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n911), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n909), .A2(KEYINPUT41), .A3(new_n910), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n929), .A2(new_n933), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n934), .A2(new_n935), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n910), .A4(new_n909), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G37), .B1(new_n946), .B2(new_n902), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n911), .A2(new_n941), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(new_n917), .B2(new_n936), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n948), .B1(new_n950), .B2(new_n901), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n936), .A2(new_n939), .A3(new_n940), .ZN(new_n952));
  INV_X1    g527(.A(new_n949), .ZN(new_n953));
  AND4_X1   g528(.A1(new_n948), .A2(new_n952), .A3(new_n901), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n947), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n952), .A2(new_n953), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n902), .ZN(new_n960));
  OAI211_X1 g535(.A(KEYINPUT43), .B(new_n960), .C1(new_n951), .C2(new_n954), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT107), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n957), .A2(new_n964), .A3(new_n958), .A4(new_n961), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n958), .B1(new_n955), .B2(KEYINPUT43), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n956), .B(new_n960), .C1(new_n951), .C2(new_n954), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n952), .A2(new_n901), .A3(new_n953), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT105), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n956), .A4(new_n960), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n966), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n963), .A2(new_n965), .A3(new_n973), .ZN(G397));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n500), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT109), .B(G40), .Z(new_n979));
  AND4_X1   g554(.A1(new_n479), .A2(new_n473), .A3(new_n474), .A4(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n761), .B(G2067), .Z(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT110), .ZN(new_n984));
  INV_X1    g559(.A(G1996), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n741), .B(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n984), .B(new_n986), .C1(new_n731), .C2(new_n728), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n731), .B2(new_n728), .ZN(new_n988));
  INV_X1    g563(.A(G1986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n988), .B1(new_n989), .B2(new_n595), .ZN(new_n990));
  NOR2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n982), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n573), .A2(KEYINPUT116), .A3(new_n993), .A4(new_n576), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(KEYINPUT116), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n993), .A2(KEYINPUT116), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n995), .B(new_n996), .C1(new_n578), .C2(new_n579), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT45), .B1(new_n500), .B2(new_n975), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n977), .B(G1384), .C1(new_n496), .C2(new_n499), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n981), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT56), .B(G2072), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n496), .B2(new_n499), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n980), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n980), .B(KEYINPUT113), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n999), .B(new_n1004), .C1(new_n1013), .C2(G1956), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n980), .A2(new_n1005), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(G2067), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(new_n1007), .A3(new_n980), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1019), .B2(new_n749), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(new_n608), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1004), .B1(new_n1013), .B2(G1956), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1022), .A2(new_n998), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1023), .B2(KEYINPUT117), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n998), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1015), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1025), .A2(new_n1014), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT61), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g607(.A(KEYINPUT119), .B(KEYINPUT61), .C1(new_n1025), .C2(new_n1014), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1020), .A2(new_n609), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1020), .A2(new_n609), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(KEYINPUT60), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1036), .A2(KEYINPUT60), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1005), .A2(KEYINPUT45), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n978), .A2(new_n985), .A3(new_n980), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1043), .A2(KEYINPUT118), .A3(new_n985), .A4(new_n980), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT58), .B(G1341), .Z(new_n1045));
  NAND2_X1  g620(.A1(new_n1016), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1047), .A2(new_n1048), .A3(new_n557), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1047), .B2(new_n557), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1037), .B(new_n1038), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1014), .A2(KEYINPUT61), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT120), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1014), .A2(new_n1054), .A3(KEYINPUT61), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1028), .B1(new_n1034), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G303), .A2(G8), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G2090), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1013), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1971), .B1(new_n1043), .B2(new_n980), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1061), .B1(new_n1066), .B2(G8), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1008), .A2(new_n1009), .A3(G2090), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1061), .B(G8), .C1(new_n1064), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n589), .A2(KEYINPUT111), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G1981), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n697), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT49), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT112), .ZN(new_n1074));
  NAND3_X1  g649(.A1(G305), .A2(G1981), .A3(new_n1070), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1073), .A2(KEYINPUT112), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1077), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1072), .A2(new_n1079), .A3(new_n1075), .A4(new_n1074), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G8), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n980), .B2(new_n1005), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n704), .B2(G288), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT52), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n704), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1083), .B(new_n1087), .C1(new_n704), .C2(G288), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1069), .A2(new_n1084), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT125), .B1(new_n1067), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1061), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1064), .B1(new_n1013), .B2(new_n1062), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(new_n1082), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1084), .A2(new_n1088), .A3(new_n1086), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1069), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1090), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G2078), .ZN(new_n1098));
  AND4_X1   g673(.A1(G40), .A2(new_n978), .A3(new_n1098), .A4(new_n1039), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n475), .B(KEYINPUT123), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1099), .A2(KEYINPUT53), .A3(new_n479), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n978), .A2(new_n1098), .A3(new_n980), .A4(new_n1039), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1102), .A2(new_n1103), .B1(new_n1019), .B2(new_n777), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(G301), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1102), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1043), .A2(KEYINPUT53), .A3(new_n1098), .A4(new_n980), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1019), .A2(new_n777), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G171), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1105), .A2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(KEYINPUT124), .A3(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT114), .B(G2084), .Z(new_n1114));
  NAND4_X1  g689(.A1(new_n1018), .A2(new_n1007), .A3(new_n980), .A4(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(G168), .C1(new_n1002), .C2(G1966), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(G8), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1116), .A2(new_n1117), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n978), .A2(new_n980), .A3(new_n1039), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1123), .A2(new_n1114), .B1(new_n1124), .B2(new_n794), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(new_n1082), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(G286), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1097), .A2(new_n1113), .A3(new_n1128), .A4(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT54), .B1(new_n1109), .B2(G171), .ZN(new_n1133));
  AOI21_X1  g708(.A(G301), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1058), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1125), .A2(new_n1082), .A3(G286), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1093), .A2(new_n1069), .A3(new_n1095), .A4(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT63), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT115), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT115), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1138), .A2(new_n1142), .A3(new_n1139), .ZN(new_n1143));
  OAI21_X1  g718(.A(G8), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1139), .B1(new_n1144), .B2(new_n1091), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1145), .A2(new_n1095), .A3(new_n1069), .A4(new_n1137), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1141), .A2(new_n1143), .A3(new_n1146), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1120), .A2(new_n1121), .B1(G286), .B2(new_n1126), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1110), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1128), .A2(KEYINPUT62), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n1097), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1069), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1095), .A2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1081), .A2(G1976), .A3(G288), .ZN(new_n1155));
  NOR2_X1   g730(.A1(G305), .A2(G1981), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1083), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1147), .A2(new_n1152), .A3(new_n1154), .A4(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n992), .B1(new_n1136), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n984), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n982), .B1(new_n1160), .B2(new_n741), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT46), .ZN(new_n1162));
  INV_X1    g737(.A(new_n982), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1163), .B2(G1996), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n982), .A2(KEYINPUT46), .A3(new_n985), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1161), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT47), .Z(new_n1167));
  NOR2_X1   g742(.A1(new_n728), .A2(new_n731), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n984), .A2(new_n1168), .A3(new_n986), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n761), .A2(G2067), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1163), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n988), .A2(new_n1163), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1172), .B(KEYINPUT126), .Z(new_n1173));
  NAND2_X1  g748(.A1(new_n991), .A2(new_n982), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT48), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1167), .B(new_n1171), .C1(new_n1173), .C2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1159), .A2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g752(.A1(new_n886), .A2(G319), .A3(new_n957), .A4(new_n961), .ZN(new_n1179));
  NOR3_X1   g753(.A1(G401), .A2(G227), .A3(G229), .ZN(new_n1180));
  INV_X1    g754(.A(new_n1180), .ZN(new_n1181));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1181), .ZN(G308));
  AND2_X1   g756(.A1(new_n957), .A2(new_n961), .ZN(new_n1183));
  NAND4_X1  g757(.A1(new_n1183), .A2(G319), .A3(new_n886), .A4(new_n1180), .ZN(G225));
endmodule


