//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n608, new_n611,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g034(.A(G125), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n467), .C1(new_n468), .C2(new_n461), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n469), .A2(KEYINPUT66), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT66), .B1(new_n469), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n467), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT68), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n467), .B1(new_n462), .B2(new_n463), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(G124), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n468), .B2(new_n461), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n489), .B(new_n492), .C1(new_n461), .C2(new_n468), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n467), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n484), .B2(G126), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  OR2_X1    g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  XOR2_X1   g081(.A(KEYINPUT69), .B(G88), .Z(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n501), .B2(new_n502), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n512), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G89), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n505), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n520), .A2(new_n521), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(new_n511), .A2(G52), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n505), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n515), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G171));
  NAND2_X1  g111(.A1(new_n511), .A2(G43), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n505), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n515), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT71), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  NAND2_X1  g123(.A1(new_n504), .A2(G65), .ZN(new_n549));
  INV_X1    g124(.A(G78), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT72), .B1(new_n550), .B2(new_n510), .ZN(new_n551));
  OR3_X1    g126(.A1(new_n550), .A2(new_n510), .A3(KEYINPUT72), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n553), .A2(G651), .B1(new_n506), .B2(G91), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n512), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n511), .A2(new_n557), .A3(G53), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n554), .A2(new_n559), .A3(KEYINPUT73), .ZN(new_n560));
  AOI21_X1  g135(.A(KEYINPUT73), .B1(new_n554), .B2(new_n559), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  OAI221_X1 g138(.A(new_n508), .B1(new_n509), .B2(new_n512), .C1(new_n515), .C2(new_n514), .ZN(G303));
  OAI21_X1  g139(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT74), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n506), .A2(G87), .B1(G49), .B2(new_n511), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(new_n511), .A2(G48), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n505), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n504), .A2(G61), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n573), .B1(new_n576), .B2(G651), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  NOR3_X1   g153(.A1(new_n578), .A2(KEYINPUT75), .A3(new_n515), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n572), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n580), .A2(KEYINPUT76), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n580), .A2(KEYINPUT76), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OR3_X1    g159(.A1(new_n584), .A2(KEYINPUT77), .A3(new_n515), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT77), .B1(new_n584), .B2(new_n515), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n506), .A2(G85), .B1(G47), .B2(new_n511), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n506), .A2(KEYINPUT10), .A3(G92), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n505), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n504), .A2(G66), .ZN(new_n595));
  INV_X1    g170(.A(G79), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT78), .B1(new_n596), .B2(new_n510), .ZN(new_n597));
  OR3_X1    g172(.A1(new_n596), .A2(new_n510), .A3(KEYINPUT78), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n511), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n589), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n589), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(KEYINPUT79), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(KEYINPUT79), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n606), .B(new_n607), .C1(G868), .C2(new_n608), .ZN(G297));
  OAI211_X1 g184(.A(new_n606), .B(new_n607), .C1(G868), .C2(new_n608), .ZN(G280));
  INV_X1    g185(.A(G860), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n601), .B1(G559), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT80), .ZN(G148));
  OR2_X1    g188(.A1(new_n601), .A2(G559), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g192(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n477), .A2(G135), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n467), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n625));
  AND3_X1   g200(.A1(new_n484), .A2(new_n625), .A3(G123), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n484), .B2(G123), .ZN(new_n627));
  OAI221_X1 g202(.A(new_n622), .B1(new_n623), .B2(new_n624), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  AOI22_X1  g203(.A1(G2100), .A2(new_n621), .B1(new_n628), .B2(G2096), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n621), .A2(G2100), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n629), .B(new_n630), .C1(G2096), .C2(new_n628), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT82), .Z(G156));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n638), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n645), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(G401));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  NOR2_X1   g224(.A1(G2072), .A2(G2078), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n442), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n652), .B2(KEYINPUT84), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(KEYINPUT84), .B2(new_n652), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n651), .B(KEYINPUT17), .ZN(new_n657));
  INV_X1    g232(.A(new_n649), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n654), .B(new_n656), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n652), .A2(new_n649), .A3(new_n655), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT18), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n657), .A2(new_n658), .A3(new_n655), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n671), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  AOI211_X1 g250(.A(new_n673), .B(new_n675), .C1(new_n668), .C2(new_n672), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT85), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G229));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G22), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G166), .B2(new_n685), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT88), .ZN(new_n688));
  INV_X1    g263(.A(G1971), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  MUX2_X1   g266(.A(G23), .B(G288), .S(G16), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT33), .B(G1976), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT87), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n690), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  MUX2_X1   g271(.A(G6), .B(G305), .S(G16), .Z(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT32), .B(G1981), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT34), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G25), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n477), .A2(G131), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n484), .A2(G119), .ZN(new_n708));
  OR2_X1    g283(.A1(G95), .A2(G2105), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n709), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(new_n705), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G290), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(new_n685), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n685), .B2(G24), .ZN(new_n718));
  INV_X1    g293(.A(G1986), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n715), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n719), .B2(new_n718), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n703), .A2(new_n704), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT36), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n685), .A2(G4), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n602), .B2(new_n685), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G1348), .Z(new_n726));
  NOR2_X1   g301(.A1(new_n542), .A2(new_n685), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n685), .B2(G19), .ZN(new_n728));
  INV_X1    g303(.A(G1341), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NOR2_X1   g306(.A1(G29), .A2(G33), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT25), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(new_n467), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n734), .B(new_n736), .C1(G139), .C2(new_n477), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n732), .B1(new_n737), .B2(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G2072), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n726), .A2(new_n730), .A3(new_n731), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n484), .A2(G128), .ZN(new_n741));
  INV_X1    g316(.A(G140), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n467), .A2(G116), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n741), .B1(new_n742), .B2(new_n476), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n705), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2067), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n685), .A2(G5), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G171), .B2(new_n685), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1961), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT31), .B(G11), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT90), .ZN(new_n755));
  INV_X1    g330(.A(G28), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT30), .ZN(new_n757));
  AOI21_X1  g332(.A(G29), .B1(new_n756), .B2(KEYINPUT30), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n759), .B1(new_n705), .B2(new_n628), .C1(new_n738), .C2(G2072), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n740), .A2(new_n750), .A3(new_n753), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G29), .A2(G32), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT26), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n475), .A2(G2105), .ZN(new_n765));
  INV_X1    g340(.A(G129), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n768));
  INV_X1    g343(.A(G141), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n476), .B2(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n762), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT27), .B(G1996), .Z(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G168), .A2(new_n685), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n685), .B2(G21), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n776), .B1(new_n779), .B2(G1966), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n705), .A2(G27), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n705), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT91), .ZN(new_n783));
  INV_X1    g358(.A(G2078), .ZN(new_n784));
  INV_X1    g359(.A(G2084), .ZN(new_n785));
  INV_X1    g360(.A(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(G29), .B1(new_n786), .B2(KEYINPUT24), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(KEYINPUT24), .B2(new_n786), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n473), .B2(new_n705), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n783), .A2(new_n784), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n761), .A2(new_n780), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n705), .A2(G35), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n705), .ZN(new_n793));
  INV_X1    g368(.A(G2090), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n685), .A2(G20), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT23), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n608), .B2(new_n685), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1956), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n789), .A2(new_n785), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n774), .B2(new_n775), .ZN(new_n803));
  OAI221_X1 g378(.A(new_n803), .B1(new_n784), .B2(new_n783), .C1(new_n779), .C2(G1966), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n791), .A2(new_n797), .A3(new_n801), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n723), .A2(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  AOI22_X1  g382(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n808), .A2(KEYINPUT93), .A3(new_n515), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT94), .B(G93), .Z(new_n811));
  AOI22_X1  g386(.A1(new_n506), .A2(new_n811), .B1(G55), .B2(new_n511), .ZN(new_n812));
  OAI21_X1  g387(.A(KEYINPUT93), .B1(new_n808), .B2(new_n515), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(new_n611), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT37), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n602), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n542), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n810), .A2(new_n814), .B1(new_n541), .B2(new_n539), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n819), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT95), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n611), .B1(new_n824), .B2(KEYINPUT39), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n817), .B1(new_n826), .B2(new_n827), .ZN(G145));
  XNOR2_X1  g403(.A(new_n486), .B(new_n628), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n473), .B(KEYINPUT96), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n484), .A2(G130), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n467), .A2(G118), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G142), .B2(new_n477), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n619), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n711), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT98), .Z(new_n839));
  MUX2_X1   g414(.A(new_n771), .B(new_n773), .S(new_n737), .Z(new_n840));
  INV_X1    g415(.A(G126), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n765), .A2(new_n841), .B1(new_n495), .B2(new_n496), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n843));
  INV_X1    g418(.A(new_n493), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n492), .B1(new_n475), .B2(new_n489), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n491), .A2(KEYINPUT97), .A3(new_n493), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n745), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n840), .B(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT99), .B1(new_n839), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n839), .A2(new_n850), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n839), .A2(KEYINPUT99), .A3(new_n850), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n831), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n850), .A2(new_n838), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT100), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n831), .B1(new_n839), .B2(new_n850), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n855), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g437(.A(new_n822), .B(new_n614), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n554), .A2(new_n559), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT73), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n554), .A2(new_n559), .A3(KEYINPUT73), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n602), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n601), .B1(new_n560), .B2(new_n561), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(G299), .A2(KEYINPUT101), .A3(new_n602), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(KEYINPUT41), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n869), .A2(new_n870), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n864), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n872), .A2(new_n873), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n864), .B2(new_n880), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(KEYINPUT42), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n883));
  NAND2_X1  g458(.A1(G288), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n566), .A2(KEYINPUT102), .A3(new_n567), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(G305), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G290), .B(G303), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n884), .B(new_n885), .C1(new_n581), .C2(new_n582), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n887), .B2(new_n889), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n881), .A2(KEYINPUT42), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n882), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n882), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(G868), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(G868), .B2(new_n815), .ZN(G295));
  OAI21_X1  g473(.A(new_n897), .B1(G868), .B2(new_n815), .ZN(G331));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n872), .A2(new_n876), .A3(new_n873), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n901), .A2(KEYINPUT105), .B1(KEYINPUT41), .B2(new_n875), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n872), .A2(new_n903), .A3(new_n876), .A4(new_n873), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n820), .A2(G301), .A3(new_n821), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(G301), .B1(new_n820), .B2(new_n821), .ZN(new_n909));
  OAI21_X1  g484(.A(G286), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n822), .A2(G171), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(G168), .A3(new_n907), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n905), .A2(new_n906), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n890), .B2(new_n891), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n887), .A2(new_n889), .ZN(new_n918));
  INV_X1    g493(.A(new_n888), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(KEYINPUT104), .A3(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n913), .B1(new_n902), .B2(new_n904), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n913), .A2(new_n880), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT106), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n915), .B(new_n923), .C1(new_n924), .C2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n910), .A2(new_n912), .A3(new_n874), .A4(new_n877), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n892), .A3(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n929), .A2(new_n860), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n900), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n917), .A2(new_n922), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n928), .B2(new_n925), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n929), .A2(new_n860), .ZN(new_n934));
  XNOR2_X1  g509(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n927), .A2(new_n930), .A3(new_n935), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n936), .B1(new_n933), .B2(new_n934), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n938), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n939), .B1(new_n938), .B2(new_n943), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(G397));
  INV_X1    g521(.A(KEYINPUT127), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n848), .B2(G1384), .ZN(new_n949));
  OAI211_X1 g524(.A(G40), .B(new_n466), .C1(new_n471), .C2(new_n472), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT108), .ZN(new_n952));
  INV_X1    g527(.A(G2067), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n745), .B(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1996), .ZN(new_n955));
  INV_X1    g530(.A(new_n771), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n952), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n773), .A2(new_n951), .A3(new_n955), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n711), .B(new_n714), .Z(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n952), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n951), .ZN(new_n963));
  XNOR2_X1  g538(.A(G290), .B(new_n719), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT55), .ZN(new_n969));
  INV_X1    g544(.A(G8), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n969), .B1(G166), .B2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(G303), .A2(KEYINPUT109), .A3(KEYINPUT55), .A4(G8), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n491), .A2(KEYINPUT97), .A3(new_n493), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT97), .B1(new_n491), .B2(new_n493), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n498), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(KEYINPUT45), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(G1384), .B1(new_n494), .B2(new_n498), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n979), .A2(KEYINPUT45), .ZN(new_n980));
  INV_X1    g555(.A(new_n950), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n689), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n950), .B1(new_n984), .B2(new_n979), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n846), .A2(new_n847), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n986), .B2(new_n498), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n985), .B(new_n794), .C1(new_n987), .C2(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n970), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n984), .B1(new_n976), .B2(new_n977), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n979), .A2(new_n984), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n981), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n995), .A2(new_n794), .B1(new_n982), .B2(new_n689), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT113), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n973), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n950), .B1(new_n987), .B2(KEYINPUT45), .ZN(new_n999));
  AOI21_X1  g574(.A(G1971), .B1(new_n999), .B2(new_n980), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n984), .B1(new_n848), .B2(G1384), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n1002));
  AOI211_X1 g577(.A(G2090), .B(new_n950), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(G8), .B(new_n973), .C1(new_n1000), .C2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n566), .A2(G1976), .A3(new_n567), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1005), .A2(KEYINPUT111), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(KEYINPUT111), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g583(.A(KEYINPUT110), .B(new_n970), .C1(new_n987), .C2(new_n981), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n981), .A2(new_n976), .A3(new_n977), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(G8), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1008), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT52), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT112), .B(G1976), .Z(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(G288), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1008), .B(new_n1016), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n848), .A2(G1384), .A3(new_n950), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT110), .B1(new_n1018), .B2(new_n970), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1011), .A2(new_n1010), .A3(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n572), .B(new_n1022), .C1(new_n577), .C2(new_n579), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n578), .A2(new_n515), .ZN(new_n1024));
  OAI21_X1  g599(.A(G1981), .B1(new_n571), .B2(new_n1024), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1023), .A2(KEYINPUT49), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT49), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1021), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1004), .A2(new_n1014), .A3(new_n1017), .A4(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n998), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n950), .A2(G2084), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n950), .B1(KEYINPUT45), .B2(new_n979), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1966), .B1(new_n949), .B2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(G8), .B(G168), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT63), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1966), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT45), .B1(new_n976), .B2(new_n977), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n979), .A2(KEYINPUT45), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n981), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1040), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT50), .B1(new_n976), .B2(new_n977), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1002), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1032), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1048), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1049));
  OAI21_X1  g624(.A(G8), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1029), .A2(new_n1017), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1021), .B2(new_n1008), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1052), .A2(new_n1056), .A3(new_n1057), .A4(new_n1004), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT63), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1037), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n950), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1061), .A2(new_n794), .B1(new_n982), .B2(new_n689), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1051), .B1(new_n1062), .B2(new_n970), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT114), .B1(new_n1030), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1058), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1039), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1004), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1029), .ZN(new_n1069));
  OR2_X1    g644(.A1(G288), .A2(G1976), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1023), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1068), .A2(new_n1056), .B1(new_n1071), .B2(new_n1021), .ZN(new_n1072));
  OAI21_X1  g647(.A(G8), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n970), .B1(new_n527), .B2(new_n528), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1073), .A2(KEYINPUT122), .A3(KEYINPUT51), .A4(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT51), .B1(new_n1074), .B2(KEYINPUT122), .ZN(new_n1077));
  OAI211_X1 g652(.A(G8), .B(new_n1077), .C1(new_n1048), .C2(G286), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n1048), .B2(new_n1074), .ZN(new_n1080));
  AOI211_X1 g655(.A(KEYINPUT121), .B(new_n1075), .C1(new_n1044), .C2(new_n1047), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1076), .B(new_n1078), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT62), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1074), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT121), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1048), .A2(new_n1079), .A3(new_n1074), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1030), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n991), .A2(new_n997), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1051), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n981), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1094));
  INV_X1    g669(.A(G1961), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n978), .A2(new_n980), .A3(new_n784), .A4(new_n981), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(G2078), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n949), .A2(new_n1035), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1096), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G171), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1091), .A2(new_n1093), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1072), .B1(new_n1090), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1067), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1096), .A2(new_n1099), .A3(G301), .A4(new_n1101), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1108), .A2(KEYINPUT54), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1061), .B2(G1961), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1094), .A2(KEYINPUT123), .A3(new_n1095), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n999), .A2(new_n949), .A3(new_n1100), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1111), .A2(new_n1112), .A3(new_n1099), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G171), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1091), .A2(new_n1116), .A3(new_n1093), .A4(new_n1082), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1103), .B1(new_n1114), .B2(G171), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT124), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n865), .A2(KEYINPUT57), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n554), .B2(new_n559), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1956), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n992), .B2(new_n994), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1126), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1128), .A2(new_n1130), .A3(new_n1126), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1134), .A2(KEYINPUT61), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n542), .A2(KEYINPUT119), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n978), .A2(new_n980), .A3(new_n955), .A4(new_n981), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(new_n729), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1011), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1137), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1138), .A2(new_n1137), .A3(new_n1141), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1136), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1133), .A2(new_n1135), .B1(new_n1145), .B2(KEYINPUT59), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT115), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1011), .B2(G2067), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1018), .A2(KEYINPUT115), .A3(new_n953), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1148), .B(new_n1149), .C1(new_n1061), .C2(G1348), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n601), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT120), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1150), .A2(KEYINPUT120), .A3(new_n1151), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1153), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1126), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT61), .B1(new_n1160), .B2(new_n1134), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1144), .ZN(new_n1163));
  OAI211_X1 g738(.A(KEYINPUT119), .B(new_n542), .C1(new_n1163), .C2(new_n1142), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1161), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1156), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1166), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1146), .A2(new_n1157), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1150), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1133), .B1(new_n601), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1134), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1077), .A2(new_n1173), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1174), .A2(new_n1076), .B1(new_n1109), .B2(new_n1115), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1175), .A2(new_n1176), .A3(new_n1120), .A4(new_n1031), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1122), .A2(new_n1172), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n965), .B1(new_n1107), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n954), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n952), .B1(new_n771), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT46), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n951), .A2(new_n955), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1183), .A2(new_n1182), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT125), .ZN(new_n1187));
  OR3_X1    g762(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1185), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1189));
  AOI21_X1  g764(.A(KEYINPUT47), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n719), .A3(new_n716), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT48), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n962), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n712), .A2(new_n714), .ZN(new_n1194));
  OAI22_X1  g769(.A1(new_n960), .A2(new_n1194), .B1(G2067), .B2(new_n745), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n952), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1190), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1188), .A2(KEYINPUT47), .A3(new_n1189), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n947), .B1(new_n1179), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1199), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n1202), .A2(new_n1190), .A3(new_n1197), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1031), .A2(new_n1083), .A3(new_n1104), .A4(new_n1089), .ZN(new_n1204));
  OAI211_X1 g779(.A(new_n1204), .B(new_n1072), .C1(new_n1039), .C2(new_n1066), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1175), .A2(new_n1120), .A3(new_n1031), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1206), .A2(KEYINPUT124), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1205), .B1(new_n1207), .B2(new_n1177), .ZN(new_n1208));
  OAI211_X1 g783(.A(KEYINPUT127), .B(new_n1203), .C1(new_n1208), .C2(new_n965), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1201), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g785(.A1(new_n665), .A2(G319), .ZN(new_n1212));
  NOR3_X1   g786(.A1(G229), .A2(G401), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n940), .A2(new_n941), .ZN(new_n1214));
  AND3_X1   g788(.A1(new_n1213), .A2(new_n861), .A3(new_n1214), .ZN(G308));
  NAND3_X1  g789(.A1(new_n1213), .A2(new_n861), .A3(new_n1214), .ZN(G225));
endmodule


