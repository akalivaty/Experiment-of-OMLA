

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761;

  NOR2_X1 U363 ( .A1(n706), .A2(n705), .ZN(n702) );
  XNOR2_X2 U364 ( .A(KEYINPUT64), .B(G953), .ZN(n637) );
  XNOR2_X2 U365 ( .A(n388), .B(G101), .ZN(n499) );
  XNOR2_X2 U366 ( .A(KEYINPUT3), .B(G119), .ZN(n388) );
  INV_X1 U367 ( .A(n710), .ZN(n587) );
  AND2_X1 U368 ( .A1(n391), .A2(KEYINPUT56), .ZN(n390) );
  XNOR2_X1 U369 ( .A(n598), .B(KEYINPUT80), .ZN(n679) );
  XNOR2_X1 U370 ( .A(n382), .B(n381), .ZN(n725) );
  XNOR2_X1 U371 ( .A(n527), .B(n526), .ZN(n684) );
  AND2_X1 U372 ( .A1(n411), .A2(n408), .ZN(n407) );
  XNOR2_X1 U373 ( .A(n433), .B(n432), .ZN(n586) );
  XNOR2_X1 U374 ( .A(n509), .B(n508), .ZN(n744) );
  XNOR2_X2 U375 ( .A(n733), .B(n447), .ZN(n642) );
  XNOR2_X2 U376 ( .A(n437), .B(n436), .ZN(n733) );
  NOR2_X1 U377 ( .A1(n528), .A2(n705), .ZN(n588) );
  NOR2_X1 U378 ( .A1(G902), .A2(n665), .ZN(n433) );
  INV_X1 U379 ( .A(G107), .ZN(n434) );
  INV_X1 U380 ( .A(n662), .ZN(n398) );
  INV_X1 U381 ( .A(n600), .ZN(n353) );
  XNOR2_X1 U382 ( .A(n558), .B(KEYINPUT84), .ZN(n576) );
  NOR2_X1 U383 ( .A1(G953), .A2(G237), .ZN(n467) );
  INV_X1 U384 ( .A(G143), .ZN(n460) );
  XNOR2_X1 U385 ( .A(G131), .B(G122), .ZN(n468) );
  XOR2_X1 U386 ( .A(KEYINPUT68), .B(G140), .Z(n508) );
  XNOR2_X1 U387 ( .A(n478), .B(n342), .ZN(n745) );
  XNOR2_X1 U388 ( .A(KEYINPUT4), .B(G131), .ZN(n428) );
  INV_X1 U389 ( .A(G237), .ZN(n448) );
  INV_X1 U390 ( .A(n589), .ZN(n370) );
  NAND2_X1 U391 ( .A1(n406), .A2(n404), .ZN(n403) );
  NAND2_X1 U392 ( .A1(n362), .A2(n613), .ZN(n751) );
  XNOR2_X1 U393 ( .A(n364), .B(n363), .ZN(n362) );
  INV_X1 U394 ( .A(KEYINPUT48), .ZN(n363) );
  XNOR2_X1 U395 ( .A(G113), .B(G104), .ZN(n462) );
  XNOR2_X1 U396 ( .A(G104), .B(G107), .ZN(n424) );
  XNOR2_X1 U397 ( .A(n745), .B(n429), .ZN(n503) );
  INV_X1 U398 ( .A(G146), .ZN(n429) );
  NAND2_X1 U399 ( .A1(n401), .A2(n351), .ZN(n399) );
  OR2_X1 U400 ( .A1(n643), .A2(G210), .ZN(n400) );
  INV_X1 U401 ( .A(KEYINPUT33), .ZN(n381) );
  NAND2_X1 U402 ( .A1(n701), .A2(n379), .ZN(n382) );
  NOR2_X1 U403 ( .A1(n546), .A2(n380), .ZN(n379) );
  XNOR2_X1 U404 ( .A(n585), .B(KEYINPUT41), .ZN(n724) );
  NOR2_X1 U405 ( .A1(n579), .A2(n584), .ZN(n580) );
  XNOR2_X1 U406 ( .A(n591), .B(n590), .ZN(n592) );
  NOR2_X1 U407 ( .A1(n653), .A2(G902), .ZN(n521) );
  INV_X1 U408 ( .A(n637), .ZN(n752) );
  XNOR2_X1 U409 ( .A(n481), .B(n480), .ZN(n373) );
  NOR2_X1 U410 ( .A1(n643), .A2(KEYINPUT56), .ZN(n395) );
  NAND2_X1 U411 ( .A1(n398), .A2(n397), .ZN(n391) );
  NOR2_X1 U412 ( .A1(n679), .A2(n695), .ZN(n599) );
  INV_X1 U413 ( .A(G224), .ZN(n438) );
  INV_X1 U414 ( .A(n584), .ZN(n691) );
  NOR2_X1 U415 ( .A1(n405), .A2(KEYINPUT85), .ZN(n404) );
  NOR2_X1 U416 ( .A1(n417), .A2(n410), .ZN(n409) );
  INV_X1 U417 ( .A(KEYINPUT85), .ZN(n410) );
  NAND2_X1 U418 ( .A1(n357), .A2(n356), .ZN(n378) );
  AND2_X1 U419 ( .A1(n575), .A2(n559), .ZN(n356) );
  INV_X1 U420 ( .A(KEYINPUT44), .ZN(n377) );
  XNOR2_X1 U421 ( .A(n368), .B(G143), .ZN(n440) );
  INV_X1 U422 ( .A(G128), .ZN(n368) );
  INV_X1 U423 ( .A(KEYINPUT65), .ZN(n626) );
  NAND2_X1 U424 ( .A1(G234), .A2(G237), .ZN(n453) );
  XNOR2_X1 U425 ( .A(n578), .B(n361), .ZN(n584) );
  INV_X1 U426 ( .A(KEYINPUT38), .ZN(n361) );
  NAND2_X1 U427 ( .A1(n616), .A2(n449), .ZN(n416) );
  NAND2_X1 U428 ( .A1(n615), .A2(n415), .ZN(n414) );
  INV_X1 U429 ( .A(n449), .ZN(n415) );
  NAND2_X1 U430 ( .A1(n588), .A2(n343), .ZN(n591) );
  XOR2_X1 U431 ( .A(G113), .B(G116), .Z(n495) );
  XNOR2_X1 U432 ( .A(G137), .B(G110), .ZN(n511) );
  XNOR2_X1 U433 ( .A(G128), .B(G119), .ZN(n510) );
  XNOR2_X1 U434 ( .A(n483), .B(n482), .ZN(n516) );
  NAND2_X1 U435 ( .A1(n752), .A2(G234), .ZN(n483) );
  INV_X1 U436 ( .A(KEYINPUT9), .ZN(n479) );
  XNOR2_X1 U437 ( .A(n440), .B(n367), .ZN(n478) );
  INV_X1 U438 ( .A(G134), .ZN(n367) );
  XNOR2_X1 U439 ( .A(n470), .B(n421), .ZN(n471) );
  INV_X1 U440 ( .A(n751), .ZN(n385) );
  NOR2_X1 U441 ( .A1(n725), .A2(n564), .ZN(n548) );
  NAND2_X1 U442 ( .A1(n371), .A2(n369), .ZN(n579) );
  XNOR2_X1 U443 ( .A(n537), .B(n538), .ZN(n371) );
  NOR2_X1 U444 ( .A1(n561), .A2(n370), .ZN(n369) );
  XNOR2_X1 U445 ( .A(n484), .B(n499), .ZN(n437) );
  XNOR2_X1 U446 ( .A(KEYINPUT16), .B(G110), .ZN(n435) );
  INV_X1 U447 ( .A(G953), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n503), .B(n383), .ZN(n665) );
  XNOR2_X1 U449 ( .A(n427), .B(n384), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n430), .B(G101), .ZN(n384) );
  XNOR2_X1 U451 ( .A(n359), .B(n349), .ZN(n756) );
  NOR2_X1 U452 ( .A1(n724), .A2(n360), .ZN(n359) );
  NOR2_X1 U453 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U454 ( .A1(n525), .A2(n524), .ZN(n555) );
  INV_X1 U455 ( .A(KEYINPUT102), .ZN(n526) );
  NOR2_X1 U456 ( .A1(n398), .A2(n656), .ZN(n660) );
  AND2_X1 U457 ( .A1(n396), .A2(n394), .ZN(n393) );
  XOR2_X1 U458 ( .A(n344), .B(n428), .Z(n342) );
  INV_X1 U459 ( .A(n643), .ZN(n397) );
  AND2_X1 U460 ( .A1(n587), .A2(n589), .ZN(n343) );
  XOR2_X1 U461 ( .A(KEYINPUT69), .B(G137), .Z(n344) );
  OR2_X1 U462 ( .A1(n689), .A2(n628), .ZN(n345) );
  AND2_X1 U463 ( .A1(n606), .A2(n543), .ZN(n346) );
  AND2_X1 U464 ( .A1(n413), .A2(n416), .ZN(n347) );
  AND2_X1 U465 ( .A1(n416), .A2(n690), .ZN(n348) );
  XOR2_X1 U466 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n349) );
  XNOR2_X1 U467 ( .A(KEYINPUT46), .B(KEYINPUT83), .ZN(n350) );
  AND2_X1 U468 ( .A1(n400), .A2(n654), .ZN(n351) );
  XNOR2_X2 U469 ( .A(n602), .B(n452), .ZN(n595) );
  XNOR2_X1 U470 ( .A(n378), .B(n377), .ZN(n376) );
  XNOR2_X2 U471 ( .A(n493), .B(n420), .ZN(n419) );
  XNOR2_X2 U472 ( .A(n505), .B(n630), .ZN(n710) );
  AND2_X1 U473 ( .A1(n601), .A2(n352), .ZN(n609) );
  NOR2_X1 U474 ( .A1(n757), .A2(n353), .ZN(n352) );
  NOR2_X2 U475 ( .A1(n592), .A2(n593), .ZN(n597) );
  XNOR2_X2 U476 ( .A(n354), .B(KEYINPUT45), .ZN(n619) );
  NAND2_X1 U477 ( .A1(n376), .A2(n577), .ZN(n354) );
  XNOR2_X2 U478 ( .A(n387), .B(n434), .ZN(n484) );
  XNOR2_X2 U479 ( .A(n355), .B(KEYINPUT0), .ZN(n547) );
  NOR2_X2 U480 ( .A1(n595), .A2(n459), .ZN(n355) );
  INV_X1 U481 ( .A(n576), .ZN(n357) );
  NAND2_X1 U482 ( .A1(n358), .A2(n625), .ZN(n627) );
  NAND2_X1 U483 ( .A1(n618), .A2(n619), .ZN(n358) );
  NAND2_X1 U484 ( .A1(n597), .A2(n596), .ZN(n598) );
  INV_X1 U485 ( .A(n597), .ZN(n360) );
  NAND2_X1 U486 ( .A1(n347), .A2(n417), .ZN(n578) );
  NAND2_X1 U487 ( .A1(n366), .A2(n365), .ZN(n364) );
  XNOR2_X1 U488 ( .A(n594), .B(n350), .ZN(n365) );
  XNOR2_X1 U489 ( .A(n609), .B(KEYINPUT70), .ZN(n366) );
  XNOR2_X1 U490 ( .A(n486), .B(n372), .ZN(n658) );
  XNOR2_X1 U491 ( .A(n478), .B(n373), .ZN(n372) );
  NAND2_X1 U492 ( .A1(n374), .A2(n684), .ZN(n604) );
  NOR2_X1 U493 ( .A1(n546), .A2(n375), .ZN(n374) );
  NAND2_X1 U494 ( .A1(n588), .A2(n589), .ZN(n375) );
  NAND2_X1 U495 ( .A1(n701), .A2(n702), .ZN(n563) );
  INV_X1 U496 ( .A(n702), .ZN(n380) );
  XNOR2_X1 U497 ( .A(n426), .B(n423), .ZN(n427) );
  XNOR2_X1 U498 ( .A(n627), .B(n626), .ZN(n629) );
  NAND2_X1 U499 ( .A1(n629), .A2(n345), .ZN(n657) );
  XNOR2_X2 U500 ( .A(n521), .B(n520), .ZN(n706) );
  NAND2_X1 U501 ( .A1(n619), .A2(n385), .ZN(n689) );
  AND2_X1 U502 ( .A1(n619), .A2(n386), .ZN(n741) );
  XNOR2_X2 U503 ( .A(G122), .B(G116), .ZN(n387) );
  NAND2_X1 U504 ( .A1(n662), .A2(n402), .ZN(n401) );
  NAND2_X1 U505 ( .A1(n393), .A2(n389), .ZN(G51) );
  NAND2_X1 U506 ( .A1(n392), .A2(n390), .ZN(n389) );
  INV_X1 U507 ( .A(n399), .ZN(n392) );
  NAND2_X1 U508 ( .A1(n398), .A2(n395), .ZN(n394) );
  NAND2_X1 U509 ( .A1(n399), .A2(n644), .ZN(n396) );
  AND2_X1 U510 ( .A1(n643), .A2(G210), .ZN(n402) );
  NAND2_X2 U511 ( .A1(n407), .A2(n403), .ZN(n602) );
  INV_X1 U512 ( .A(n417), .ZN(n405) );
  INV_X1 U513 ( .A(n412), .ZN(n406) );
  INV_X1 U514 ( .A(n409), .ZN(n408) );
  NAND2_X1 U515 ( .A1(n412), .A2(KEYINPUT85), .ZN(n411) );
  NAND2_X1 U516 ( .A1(n413), .A2(n348), .ZN(n412) );
  OR2_X2 U517 ( .A1(n642), .A2(n414), .ZN(n413) );
  NAND2_X1 U518 ( .A1(n642), .A2(n449), .ZN(n417) );
  NAND2_X1 U519 ( .A1(n419), .A2(n346), .ZN(n545) );
  NAND2_X1 U520 ( .A1(n419), .A2(n418), .ZN(n525) );
  INV_X1 U521 ( .A(n701), .ZN(n418) );
  INV_X1 U522 ( .A(KEYINPUT22), .ZN(n420) );
  XNOR2_X2 U523 ( .A(n553), .B(n552), .ZN(n761) );
  XOR2_X1 U524 ( .A(n469), .B(n468), .Z(n421) );
  AND2_X1 U525 ( .A1(n519), .A2(G217), .ZN(n422) );
  XOR2_X1 U526 ( .A(n425), .B(n424), .Z(n423) );
  XNOR2_X1 U527 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n464) );
  XNOR2_X1 U528 ( .A(n479), .B(KEYINPUT100), .ZN(n480) );
  INV_X1 U529 ( .A(KEYINPUT8), .ZN(n482) );
  XNOR2_X1 U530 ( .A(KEYINPUT106), .B(KEYINPUT28), .ZN(n590) );
  XNOR2_X1 U531 ( .A(n431), .B(G469), .ZN(n432) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n646) );
  XNOR2_X1 U533 ( .A(n473), .B(n645), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(n568) );
  XOR2_X1 U535 ( .A(n508), .B(G110), .Z(n426) );
  XOR2_X1 U536 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n425) );
  NAND2_X1 U537 ( .A1(G227), .A2(n752), .ZN(n430) );
  XNOR2_X1 U538 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n431) );
  XNOR2_X2 U539 ( .A(n586), .B(KEYINPUT1), .ZN(n701) );
  XNOR2_X1 U540 ( .A(n462), .B(n435), .ZN(n436) );
  NOR2_X1 U541 ( .A1(n637), .A2(n438), .ZN(n439) );
  XNOR2_X1 U542 ( .A(n440), .B(n439), .ZN(n446) );
  XNOR2_X2 U543 ( .A(G146), .B(G125), .ZN(n463) );
  XNOR2_X1 U544 ( .A(KEYINPUT18), .B(KEYINPUT77), .ZN(n441) );
  XNOR2_X1 U545 ( .A(n463), .B(n441), .ZN(n444) );
  XNOR2_X1 U546 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n442) );
  XNOR2_X1 U547 ( .A(n442), .B(KEYINPUT88), .ZN(n443) );
  XNOR2_X1 U548 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U549 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U550 ( .A(KEYINPUT15), .B(G902), .ZN(n615) );
  INV_X1 U551 ( .A(n615), .ZN(n616) );
  INV_X1 U552 ( .A(G902), .ZN(n504) );
  NAND2_X1 U553 ( .A1(n504), .A2(n448), .ZN(n450) );
  NAND2_X1 U554 ( .A1(n450), .A2(G210), .ZN(n449) );
  NAND2_X1 U555 ( .A1(n450), .A2(G214), .ZN(n690) );
  XNOR2_X1 U556 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n451) );
  XNOR2_X1 U557 ( .A(n451), .B(KEYINPUT66), .ZN(n452) );
  XNOR2_X1 U558 ( .A(n453), .B(KEYINPUT14), .ZN(n457) );
  NAND2_X1 U559 ( .A1(G952), .A2(n457), .ZN(n454) );
  XOR2_X1 U560 ( .A(KEYINPUT89), .B(n454), .Z(n723) );
  NOR2_X1 U561 ( .A1(G953), .A2(n723), .ZN(n456) );
  INV_X1 U562 ( .A(KEYINPUT90), .ZN(n455) );
  XNOR2_X1 U563 ( .A(n456), .B(n455), .ZN(n532) );
  NAND2_X1 U564 ( .A1(G902), .A2(n457), .ZN(n529) );
  XNOR2_X1 U565 ( .A(G898), .B(KEYINPUT91), .ZN(n738) );
  NAND2_X1 U566 ( .A1(G953), .A2(n738), .ZN(n734) );
  OR2_X1 U567 ( .A1(n529), .A2(n734), .ZN(n458) );
  AND2_X1 U568 ( .A1(n532), .A2(n458), .ZN(n459) );
  XNOR2_X1 U569 ( .A(n460), .B(G140), .ZN(n461) );
  XNOR2_X1 U570 ( .A(n462), .B(n461), .ZN(n466) );
  XNOR2_X1 U571 ( .A(n463), .B(KEYINPUT10), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(n464), .ZN(n465) );
  XOR2_X1 U573 ( .A(n466), .B(n465), .Z(n472) );
  XOR2_X1 U574 ( .A(KEYINPUT73), .B(n467), .Z(n496) );
  NAND2_X1 U575 ( .A1(G214), .A2(n496), .ZN(n470) );
  XOR2_X1 U576 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n469) );
  NOR2_X1 U577 ( .A1(G902), .A2(n646), .ZN(n475) );
  XNOR2_X1 U578 ( .A(KEYINPUT13), .B(KEYINPUT97), .ZN(n473) );
  INV_X1 U579 ( .A(G475), .ZN(n645) );
  XOR2_X1 U580 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n477) );
  XNOR2_X1 U581 ( .A(KEYINPUT101), .B(KEYINPUT98), .ZN(n476) );
  XNOR2_X1 U582 ( .A(n477), .B(n476), .ZN(n481) );
  NAND2_X1 U583 ( .A1(G217), .A2(n516), .ZN(n485) );
  XNOR2_X1 U584 ( .A(n485), .B(n484), .ZN(n486) );
  NAND2_X1 U585 ( .A1(n658), .A2(n504), .ZN(n487) );
  INV_X1 U586 ( .A(G478), .ZN(n656) );
  XNOR2_X1 U587 ( .A(n487), .B(n656), .ZN(n567) );
  INV_X1 U588 ( .A(n567), .ZN(n539) );
  NOR2_X1 U589 ( .A1(n568), .A2(n539), .ZN(n583) );
  NAND2_X1 U590 ( .A1(G234), .A2(n615), .ZN(n488) );
  XNOR2_X1 U591 ( .A(KEYINPUT20), .B(n488), .ZN(n519) );
  AND2_X1 U592 ( .A1(n519), .A2(G221), .ZN(n490) );
  INV_X1 U593 ( .A(KEYINPUT21), .ZN(n489) );
  XNOR2_X1 U594 ( .A(n490), .B(n489), .ZN(n705) );
  INV_X1 U595 ( .A(n705), .ZN(n491) );
  AND2_X1 U596 ( .A1(n583), .A2(n491), .ZN(n492) );
  NAND2_X1 U597 ( .A1(n547), .A2(n492), .ZN(n493) );
  INV_X1 U598 ( .A(n525), .ZN(n523) );
  XNOR2_X1 U599 ( .A(KEYINPUT5), .B(KEYINPUT93), .ZN(n494) );
  XNOR2_X1 U600 ( .A(n495), .B(n494), .ZN(n498) );
  NAND2_X1 U601 ( .A1(n496), .A2(G210), .ZN(n497) );
  XNOR2_X1 U602 ( .A(n498), .B(n497), .ZN(n501) );
  INV_X1 U603 ( .A(n499), .ZN(n500) );
  XNOR2_X1 U604 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U605 ( .A(n503), .B(n502), .ZN(n633) );
  NAND2_X1 U606 ( .A1(n633), .A2(n504), .ZN(n505) );
  INV_X1 U607 ( .A(G472), .ZN(n630) );
  INV_X1 U608 ( .A(KEYINPUT6), .ZN(n506) );
  XNOR2_X1 U609 ( .A(n710), .B(n506), .ZN(n546) );
  INV_X1 U610 ( .A(n507), .ZN(n509) );
  XNOR2_X1 U611 ( .A(n510), .B(KEYINPUT23), .ZN(n514) );
  XOR2_X1 U612 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n512) );
  XNOR2_X1 U613 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U614 ( .A(n513), .B(n514), .Z(n515) );
  XNOR2_X1 U615 ( .A(n744), .B(n515), .ZN(n518) );
  NAND2_X1 U616 ( .A1(G221), .A2(n516), .ZN(n517) );
  XNOR2_X1 U617 ( .A(n518), .B(n517), .ZN(n653) );
  XNOR2_X1 U618 ( .A(KEYINPUT25), .B(n422), .ZN(n520) );
  INV_X1 U619 ( .A(n706), .ZN(n528) );
  AND2_X1 U620 ( .A1(n546), .A2(n528), .ZN(n522) );
  NAND2_X1 U621 ( .A1(n523), .A2(n522), .ZN(n572) );
  XNOR2_X1 U622 ( .A(n572), .B(G101), .ZN(G3) );
  NAND2_X1 U623 ( .A1(n710), .A2(n706), .ZN(n524) );
  XOR2_X1 U624 ( .A(G110), .B(n555), .Z(G12) );
  XOR2_X1 U625 ( .A(KEYINPUT103), .B(KEYINPUT43), .Z(n535) );
  NAND2_X1 U626 ( .A1(n567), .A2(n568), .ZN(n527) );
  NOR2_X1 U627 ( .A1(G900), .A2(n529), .ZN(n530) );
  NAND2_X1 U628 ( .A1(n530), .A2(n637), .ZN(n531) );
  NAND2_X1 U629 ( .A1(n532), .A2(n531), .ZN(n589) );
  NOR2_X1 U630 ( .A1(n604), .A2(n701), .ZN(n533) );
  NAND2_X1 U631 ( .A1(n533), .A2(n690), .ZN(n534) );
  XNOR2_X1 U632 ( .A(n535), .B(n534), .ZN(n536) );
  AND2_X1 U633 ( .A1(n536), .A2(n578), .ZN(n612) );
  XOR2_X1 U634 ( .A(n612), .B(G140), .Z(G42) );
  NAND2_X1 U635 ( .A1(n586), .A2(n702), .ZN(n561) );
  XOR2_X1 U636 ( .A(KEYINPUT30), .B(KEYINPUT104), .Z(n538) );
  NAND2_X1 U637 ( .A1(n690), .A2(n587), .ZN(n537) );
  NAND2_X1 U638 ( .A1(n568), .A2(n539), .ZN(n549) );
  NOR2_X1 U639 ( .A1(n579), .A2(n549), .ZN(n541) );
  INV_X1 U640 ( .A(n578), .ZN(n540) );
  NAND2_X1 U641 ( .A1(n541), .A2(n540), .ZN(n600) );
  XNOR2_X1 U642 ( .A(n600), .B(G143), .ZN(G45) );
  INV_X1 U643 ( .A(KEYINPUT87), .ZN(n542) );
  XNOR2_X1 U644 ( .A(n701), .B(n542), .ZN(n606) );
  AND2_X1 U645 ( .A1(n706), .A2(n546), .ZN(n543) );
  XNOR2_X1 U646 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n544) );
  XNOR2_X1 U647 ( .A(n545), .B(n544), .ZN(n554) );
  XOR2_X1 U648 ( .A(n554), .B(G119), .Z(G21) );
  INV_X1 U649 ( .A(n547), .ZN(n564) );
  XNOR2_X1 U650 ( .A(n548), .B(KEYINPUT34), .ZN(n551) );
  XOR2_X1 U651 ( .A(n549), .B(KEYINPUT78), .Z(n550) );
  NAND2_X1 U652 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U653 ( .A(KEYINPUT35), .B(KEYINPUT82), .ZN(n552) );
  INV_X1 U654 ( .A(KEYINPUT67), .ZN(n559) );
  INV_X1 U655 ( .A(n554), .ZN(n557) );
  INV_X1 U656 ( .A(n555), .ZN(n556) );
  NAND2_X1 U657 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U658 ( .A1(n559), .A2(n576), .ZN(n560) );
  NAND2_X1 U659 ( .A1(n761), .A2(n560), .ZN(n574) );
  NOR2_X1 U660 ( .A1(n561), .A2(n587), .ZN(n562) );
  AND2_X1 U661 ( .A1(n562), .A2(n547), .ZN(n672) );
  OR2_X1 U662 ( .A1(n710), .A2(n563), .ZN(n700) );
  OR2_X1 U663 ( .A1(n564), .A2(n700), .ZN(n566) );
  XNOR2_X1 U664 ( .A(KEYINPUT94), .B(KEYINPUT31), .ZN(n565) );
  XNOR2_X1 U665 ( .A(n566), .B(n565), .ZN(n687) );
  OR2_X1 U666 ( .A1(n672), .A2(n687), .ZN(n570) );
  OR2_X1 U667 ( .A1(n568), .A2(n567), .ZN(n676) );
  INV_X1 U668 ( .A(n676), .ZN(n686) );
  NOR2_X1 U669 ( .A1(n684), .A2(n686), .ZN(n695) );
  INV_X1 U670 ( .A(n695), .ZN(n569) );
  NAND2_X1 U671 ( .A1(n570), .A2(n569), .ZN(n571) );
  AND2_X1 U672 ( .A1(n572), .A2(n571), .ZN(n573) );
  AND2_X1 U673 ( .A1(n574), .A2(n573), .ZN(n577) );
  INV_X1 U674 ( .A(n761), .ZN(n575) );
  INV_X1 U675 ( .A(n684), .ZN(n680) );
  XNOR2_X1 U676 ( .A(n580), .B(KEYINPUT39), .ZN(n610) );
  NOR2_X1 U677 ( .A1(n680), .A2(n610), .ZN(n582) );
  XNOR2_X1 U678 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n581) );
  XNOR2_X1 U679 ( .A(n582), .B(n581), .ZN(n759) );
  INV_X1 U680 ( .A(n583), .ZN(n693) );
  NAND2_X1 U681 ( .A1(n691), .A2(n690), .ZN(n694) );
  NOR2_X1 U682 ( .A1(n693), .A2(n694), .ZN(n585) );
  XNOR2_X1 U683 ( .A(n586), .B(KEYINPUT105), .ZN(n593) );
  NAND2_X1 U684 ( .A1(n759), .A2(n756), .ZN(n594) );
  INV_X1 U685 ( .A(n595), .ZN(n596) );
  XNOR2_X1 U686 ( .A(n599), .B(KEYINPUT47), .ZN(n601) );
  INV_X1 U687 ( .A(n602), .ZN(n603) );
  XNOR2_X1 U688 ( .A(n605), .B(KEYINPUT36), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U690 ( .A(n608), .B(KEYINPUT109), .ZN(n757) );
  NOR2_X1 U691 ( .A1(n676), .A2(n610), .ZN(n611) );
  XNOR2_X1 U692 ( .A(n611), .B(KEYINPUT110), .ZN(n760) );
  NOR2_X1 U693 ( .A1(n760), .A2(n612), .ZN(n613) );
  AND2_X1 U694 ( .A1(KEYINPUT2), .A2(KEYINPUT81), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n621) );
  INV_X1 U696 ( .A(n621), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n624) );
  NOR2_X1 U698 ( .A1(n751), .A2(n624), .ZN(n618) );
  INV_X1 U699 ( .A(KEYINPUT81), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n620), .A2(KEYINPUT2), .ZN(n622) );
  AND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n623) );
  OR2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  INV_X1 U703 ( .A(KEYINPUT2), .ZN(n628) );
  NOR2_X1 U704 ( .A1(n657), .A2(n630), .ZN(n635) );
  XNOR2_X1 U705 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n631), .B(KEYINPUT62), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U708 ( .A(n635), .B(n634), .ZN(n638) );
  INV_X1 U709 ( .A(G952), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n637), .A2(n636), .ZN(n654) );
  NAND2_X1 U711 ( .A1(n638), .A2(n654), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n639), .B(KEYINPUT63), .ZN(G57) );
  INV_X2 U713 ( .A(n657), .ZN(n662) );
  XNOR2_X1 U714 ( .A(KEYINPUT86), .B(KEYINPUT54), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n640), .B(KEYINPUT55), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n642), .B(n641), .ZN(n643) );
  INV_X1 U717 ( .A(KEYINPUT56), .ZN(n644) );
  NOR2_X1 U718 ( .A1(n657), .A2(n645), .ZN(n648) );
  XOR2_X1 U719 ( .A(n646), .B(KEYINPUT59), .Z(n647) );
  XNOR2_X1 U720 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n649), .A2(n654), .ZN(n651) );
  INV_X1 U722 ( .A(KEYINPUT60), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n651), .B(n650), .ZN(G60) );
  NAND2_X1 U724 ( .A1(n662), .A2(G217), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n653), .B(n652), .ZN(n655) );
  INV_X1 U726 ( .A(n654), .ZN(n668) );
  NOR2_X1 U727 ( .A1(n655), .A2(n668), .ZN(G66) );
  XOR2_X1 U728 ( .A(n658), .B(KEYINPUT123), .Z(n659) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U730 ( .A1(n661), .A2(n668), .ZN(G63) );
  NAND2_X1 U731 ( .A1(n662), .A2(G469), .ZN(n667) );
  XOR2_X1 U732 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT58), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n667), .B(n666), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(G54) );
  XOR2_X1 U737 ( .A(G104), .B(KEYINPUT113), .Z(n671) );
  NAND2_X1 U738 ( .A1(n672), .A2(n684), .ZN(n670) );
  XNOR2_X1 U739 ( .A(n671), .B(n670), .ZN(G6) );
  XOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n674) );
  NAND2_X1 U741 ( .A1(n672), .A2(n686), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U743 ( .A(G107), .B(n675), .ZN(G9) );
  NOR2_X1 U744 ( .A1(n679), .A2(n676), .ZN(n678) );
  XNOR2_X1 U745 ( .A(G128), .B(KEYINPUT29), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n678), .B(n677), .ZN(G30) );
  XNOR2_X1 U747 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U749 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U750 ( .A(G146), .B(n683), .ZN(G48) );
  NAND2_X1 U751 ( .A1(n687), .A2(n684), .ZN(n685) );
  XNOR2_X1 U752 ( .A(n685), .B(G113), .ZN(G15) );
  NAND2_X1 U753 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n688), .B(G116), .ZN(G18) );
  XOR2_X1 U755 ( .A(KEYINPUT2), .B(n689), .Z(n730) );
  NOR2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U760 ( .A(n698), .B(KEYINPUT120), .ZN(n699) );
  NOR2_X1 U761 ( .A1(n725), .A2(n699), .ZN(n720) );
  INV_X1 U762 ( .A(n700), .ZN(n715) );
  XNOR2_X1 U763 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n704) );
  NOR2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U765 ( .A(n704), .B(n703), .ZN(n713) );
  NAND2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n709) );
  XNOR2_X1 U767 ( .A(KEYINPUT49), .B(KEYINPUT117), .ZN(n707) );
  XNOR2_X1 U768 ( .A(n707), .B(KEYINPUT116), .ZN(n708) );
  XNOR2_X1 U769 ( .A(n709), .B(n708), .ZN(n711) );
  NAND2_X1 U770 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U772 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U773 ( .A(n716), .B(KEYINPUT119), .ZN(n717) );
  XNOR2_X1 U774 ( .A(KEYINPUT51), .B(n717), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n724), .A2(n718), .ZN(n719) );
  NOR2_X1 U776 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U777 ( .A(n721), .B(KEYINPUT52), .ZN(n722) );
  NOR2_X1 U778 ( .A1(n723), .A2(n722), .ZN(n728) );
  NOR2_X1 U779 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U780 ( .A(KEYINPUT121), .B(n726), .Z(n727) );
  NOR2_X1 U781 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n731), .A2(G953), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n732), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U785 ( .A(KEYINPUT125), .B(n733), .Z(n735) );
  NAND2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n743) );
  XOR2_X1 U787 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n737) );
  NAND2_X1 U788 ( .A1(G224), .A2(G953), .ZN(n736) );
  XNOR2_X1 U789 ( .A(n737), .B(n736), .ZN(n739) );
  NOR2_X1 U790 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U791 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n743), .B(n742), .ZN(G69) );
  XOR2_X1 U793 ( .A(n745), .B(n744), .Z(n750) );
  XOR2_X1 U794 ( .A(G227), .B(n750), .Z(n746) );
  NAND2_X1 U795 ( .A1(n746), .A2(G900), .ZN(n747) );
  XNOR2_X1 U796 ( .A(KEYINPUT126), .B(n747), .ZN(n748) );
  NAND2_X1 U797 ( .A1(n748), .A2(G953), .ZN(n749) );
  XOR2_X1 U798 ( .A(KEYINPUT127), .B(n749), .Z(n755) );
  XOR2_X1 U799 ( .A(n751), .B(n750), .Z(n753) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n755), .A2(n754), .ZN(G72) );
  XNOR2_X1 U802 ( .A(G137), .B(n756), .ZN(G39) );
  XNOR2_X1 U803 ( .A(G125), .B(n757), .ZN(n758) );
  XNOR2_X1 U804 ( .A(n758), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U805 ( .A(G131), .B(n759), .ZN(G33) );
  XOR2_X1 U806 ( .A(G134), .B(n760), .Z(G36) );
  XOR2_X1 U807 ( .A(n761), .B(G122), .Z(G24) );
endmodule

