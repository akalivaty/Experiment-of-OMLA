//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n212), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G68), .B2(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G107), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n208), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n206), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n211), .B(new_n231), .C1(new_n233), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT64), .B(G250), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G257), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n206), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT22), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n206), .A2(G107), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT23), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT84), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT84), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n256), .A2(new_n262), .A3(new_n258), .A4(new_n259), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(KEYINPUT24), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n232), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT24), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n260), .A2(KEYINPUT84), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n264), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n205), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(G13), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n266), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n205), .A2(G33), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT25), .ZN(new_n276));
  INV_X1    g0076(.A(new_n270), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G13), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n276), .B1(new_n278), .B2(G107), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n272), .A2(KEYINPUT25), .A3(new_n218), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n275), .A2(G107), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n205), .B(G45), .C1(new_n282), .C2(KEYINPUT5), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT79), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT5), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n282), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n284), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(G264), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n213), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n215), .A2(G1698), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n295), .B(new_n296), .C1(new_n253), .C2(new_n254), .ZN(new_n297));
  INV_X1    g0097(.A(G294), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT85), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT85), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G294), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n301), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n292), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n283), .B1(new_n287), .B2(new_n288), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G274), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n293), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(G200), .B2(new_n308), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n269), .A2(new_n281), .A3(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n265), .A2(new_n232), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n253), .A2(new_n254), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT7), .B1(new_n314), .B2(new_n206), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT7), .ZN(new_n316));
  NOR4_X1   g0116(.A1(new_n253), .A2(new_n254), .A3(new_n316), .A4(G20), .ZN(new_n317));
  OAI21_X1  g0117(.A(G68), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(G58), .A2(G68), .ZN(new_n319));
  NOR2_X1   g0119(.A1(G58), .A2(G68), .ZN(new_n320));
  OAI21_X1  g0120(.A(G20), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(G20), .A2(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G159), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n313), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT73), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n321), .B2(new_n323), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n321), .A2(new_n330), .A3(new_n323), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n253), .A2(new_n254), .A3(G20), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT72), .B1(new_n335), .B2(KEYINPUT7), .ZN(new_n336));
  OR2_X1    g0136(.A1(KEYINPUT3), .A2(G33), .ZN(new_n337));
  NAND2_X1  g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n206), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(new_n316), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n317), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G68), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n334), .B(KEYINPUT16), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n329), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT8), .B(G58), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT75), .A3(new_n270), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT75), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n346), .B2(new_n277), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n273), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n272), .A2(new_n346), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n345), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n223), .A2(G1698), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n356), .B1(G223), .B2(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n357));
  INV_X1    g0157(.A(G33), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n358), .B2(new_n212), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n304), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G274), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n292), .A2(G232), .A3(new_n361), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT76), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n363), .B2(new_n364), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n360), .B(G179), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n368), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(new_n366), .B1(new_n304), .B2(new_n359), .ZN(new_n371));
  INV_X1    g0171(.A(G169), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n355), .A2(KEYINPUT18), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT77), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT18), .ZN(new_n376));
  INV_X1    g0176(.A(new_n373), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n353), .B1(new_n329), .B2(new_n344), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT77), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n355), .A2(new_n380), .A3(KEYINPUT18), .A4(new_n373), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n375), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n371), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n371), .A2(G190), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n378), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n378), .A2(KEYINPUT17), .A3(new_n384), .A4(new_n385), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n382), .A2(new_n390), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n391), .A2(KEYINPUT78), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT13), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n228), .A2(G1698), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n394), .B1(G226), .B2(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n304), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n292), .A2(new_n361), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT69), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n292), .A2(KEYINPUT69), .A3(new_n361), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(G238), .A3(new_n402), .ZN(new_n403));
  AND4_X1   g0203(.A1(new_n393), .A2(new_n398), .A3(new_n363), .A4(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n397), .A2(new_n304), .B1(G274), .B2(new_n362), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n393), .B1(new_n405), .B2(new_n403), .ZN(new_n406));
  OAI21_X1  g0206(.A(G169), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT14), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n404), .A2(new_n406), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G179), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n398), .A2(new_n363), .A3(new_n403), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT13), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n405), .A2(new_n393), .A3(new_n403), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT14), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(G169), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n408), .A2(new_n410), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n206), .A2(G33), .A3(G77), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n322), .A2(G50), .B1(G20), .B2(new_n343), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n313), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT71), .B(KEYINPUT11), .Z(new_n421));
  XNOR2_X1  g0221(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n313), .A2(new_n270), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT12), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n272), .B2(new_n343), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n278), .A2(KEYINPUT12), .A3(G68), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n422), .B1(new_n343), .B2(new_n423), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n417), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n409), .B2(G190), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT70), .B1(new_n409), .B2(new_n383), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT70), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n414), .A2(new_n431), .A3(G200), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n391), .A2(KEYINPUT78), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n392), .A2(new_n428), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT67), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n346), .A2(G20), .A3(new_n358), .ZN(new_n437));
  INV_X1    g0237(.A(G150), .ZN(new_n438));
  INV_X1    g0238(.A(new_n322), .ZN(new_n439));
  NOR3_X1   g0239(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n438), .A2(new_n439), .B1(new_n440), .B2(new_n206), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n266), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n423), .A2(G50), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT65), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n278), .A2(new_n222), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n443), .B2(new_n445), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n442), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT9), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n337), .A2(new_n338), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n294), .A2(G222), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G223), .A2(G1698), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n304), .B1(new_n451), .B2(G77), .ZN(new_n455));
  OAI221_X1 g0255(.A(new_n363), .B1(new_n223), .B2(new_n399), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(new_n309), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(new_n448), .B2(new_n449), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(G200), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n450), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n436), .B1(new_n460), .B2(KEYINPUT66), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT10), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n460), .A2(new_n436), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n436), .B(KEYINPUT10), .C1(new_n460), .C2(KEYINPUT66), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G238), .A2(G1698), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n451), .B(new_n467), .C1(new_n228), .C2(G1698), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n304), .C1(G107), .C2(new_n451), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n469), .B(new_n363), .C1(new_n225), .C2(new_n399), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n470), .A2(G179), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n278), .A2(G77), .ZN(new_n472));
  XOR2_X1   g0272(.A(KEYINPUT15), .B(G87), .Z(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(new_n206), .A3(G33), .ZN(new_n474));
  OAI221_X1 g0274(.A(new_n474), .B1(new_n206), .B2(new_n224), .C1(new_n439), .C2(new_n346), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n475), .B2(new_n266), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n423), .A2(new_n224), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n470), .A2(new_n372), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n471), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n456), .A2(new_n372), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n448), .B(new_n482), .C1(G179), .C2(new_n456), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n476), .B(new_n478), .C1(new_n309), .C2(new_n470), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n470), .A2(G200), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n466), .A2(new_n481), .A3(new_n483), .A4(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT68), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n489), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n435), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(G244), .B1(new_n253), .B2(new_n254), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n494), .A2(G1698), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(G244), .C1(new_n254), .C2(new_n253), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(G250), .B1(new_n253), .B2(new_n254), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n294), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n304), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n306), .A2(new_n304), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT80), .B1(new_n503), .B2(G257), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT80), .ZN(new_n505));
  NOR4_X1   g0305(.A1(new_n306), .A2(new_n505), .A3(new_n215), .A4(new_n304), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n307), .B(new_n502), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G200), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT81), .ZN(new_n509));
  INV_X1    g0309(.A(new_n507), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G190), .ZN(new_n511));
  OAI21_X1  g0311(.A(G107), .B1(new_n315), .B2(new_n317), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n218), .A2(KEYINPUT6), .A3(G97), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n214), .A2(new_n218), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(new_n202), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G20), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n512), .B(new_n517), .C1(new_n224), .C2(new_n439), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n266), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n278), .A2(G97), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n275), .A2(G97), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT81), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n507), .A2(new_n524), .A3(G200), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n509), .A2(new_n511), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n225), .A2(G1698), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n451), .B(new_n527), .C1(G238), .C2(G1698), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G116), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n292), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n213), .A2(KEYINPUT82), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n205), .B(G45), .C1(new_n531), .C2(G274), .ZN(new_n532));
  INV_X1    g0332(.A(G45), .ZN(new_n533));
  OAI211_X1 g0333(.A(KEYINPUT82), .B(G250), .C1(new_n533), .C2(G1), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n304), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G190), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n451), .A2(new_n206), .A3(G68), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n396), .A2(new_n206), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n539), .B(KEYINPUT19), .C1(new_n203), .C2(G87), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n396), .A2(G20), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n538), .B(new_n540), .C1(KEYINPUT19), .C2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n473), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n542), .A2(new_n266), .B1(new_n272), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(G200), .B1(new_n530), .B2(new_n535), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n275), .A2(G87), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n537), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n275), .A2(new_n473), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G179), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n536), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n372), .B1(new_n530), .B2(new_n535), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n507), .A2(new_n372), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n493), .A2(new_n494), .B1(G33), .B2(G283), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n494), .B1(new_n451), .B2(G250), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n498), .C1(new_n294), .C2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(new_n304), .B1(G274), .B2(new_n306), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n503), .A2(KEYINPUT80), .A3(G257), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n290), .A2(G257), .A3(new_n292), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n505), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n564), .A3(new_n550), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n555), .A2(new_n556), .A3(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n526), .A2(new_n554), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n308), .A2(new_n550), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G169), .B2(new_n308), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n269), .B2(new_n281), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n278), .A2(G116), .A3(new_n313), .A4(new_n274), .ZN(new_n571));
  INV_X1    g0371(.A(G116), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n272), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n265), .A2(new_n232), .B1(G20), .B2(new_n572), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n496), .B(new_n206), .C1(G33), .C2(new_n214), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT20), .B1(new_n574), .B2(new_n575), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n571), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n294), .A2(G257), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n451), .B(new_n579), .C1(new_n219), .C2(new_n294), .ZN(new_n580));
  INV_X1    g0380(.A(G303), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n314), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n304), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n290), .A2(G270), .A3(new_n292), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(new_n307), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n585), .A2(KEYINPUT21), .A3(G169), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n550), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n578), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(G169), .A3(new_n578), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT83), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(KEYINPUT83), .A3(new_n590), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n588), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n585), .A2(new_n309), .ZN(new_n596));
  AOI211_X1 g0396(.A(new_n578), .B(new_n596), .C1(G200), .C2(new_n585), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n570), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n312), .A2(new_n492), .A3(new_n567), .A4(new_n598), .ZN(G372));
  AND2_X1   g0399(.A1(new_n556), .A2(new_n565), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n554), .A2(new_n600), .A3(KEYINPUT26), .A4(new_n555), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT26), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n547), .A2(new_n553), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n566), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n526), .A2(new_n312), .A3(new_n554), .A4(new_n566), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n570), .A2(new_n595), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n553), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n492), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g0409(.A(new_n609), .B(KEYINPUT86), .Z(new_n610));
  INV_X1    g0410(.A(KEYINPUT87), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n374), .A2(new_n379), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n471), .A2(new_n479), .A3(new_n480), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n433), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n614), .A2(new_n428), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n388), .A2(new_n389), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n611), .B(new_n612), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n614), .B2(new_n428), .ZN(new_n618));
  INV_X1    g0418(.A(new_n612), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT87), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n617), .A2(new_n466), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n483), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT88), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT88), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(new_n624), .A3(new_n483), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n610), .A2(new_n626), .ZN(G369));
  NOR2_X1   g0427(.A1(new_n271), .A2(G20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n205), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G213), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(G343), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n570), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n570), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n269), .A2(new_n281), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n312), .B1(new_n639), .B2(new_n635), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n595), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n578), .A3(new_n634), .ZN(new_n643));
  INV_X1    g0443(.A(new_n578), .ZN(new_n644));
  OAI22_X1  g0444(.A1(new_n595), .A2(new_n597), .B1(new_n644), .B2(new_n635), .ZN(new_n645));
  XNOR2_X1  g0445(.A(KEYINPUT89), .B(G330), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g0448(.A(new_n648), .B(KEYINPUT90), .Z(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n642), .A2(new_n634), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n637), .B1(new_n641), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(G399));
  INV_X1    g0453(.A(new_n209), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G41), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G1), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n234), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT28), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n608), .A2(new_n635), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT29), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n567), .A2(new_n598), .A3(new_n312), .A4(new_n635), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT30), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n293), .A2(new_n305), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n585), .A2(new_n666), .A3(new_n550), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n560), .A2(new_n564), .A3(new_n536), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n665), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n510), .A2(KEYINPUT30), .A3(new_n667), .A4(new_n536), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT91), .ZN(new_n672));
  INV_X1    g0472(.A(new_n308), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n507), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n550), .A3(new_n585), .ZN(new_n675));
  INV_X1    g0475(.A(new_n536), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n308), .B1(new_n560), .B2(new_n564), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n672), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n670), .B(new_n671), .C1(new_n675), .C2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT31), .B1(new_n679), .B2(new_n634), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(KEYINPUT31), .A3(new_n634), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n664), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n646), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n663), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n660), .B1(new_n686), .B2(G1), .ZN(G364));
  NAND2_X1  g0487(.A1(new_n643), .A2(new_n645), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n646), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n628), .A2(G45), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n656), .A2(G1), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n690), .A2(new_n647), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n232), .B1(G20), .B2(new_n372), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n206), .A2(G179), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(new_n309), .A3(G200), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT99), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n451), .B1(new_n703), .B2(G283), .ZN(new_n704));
  INV_X1    g0504(.A(G326), .ZN(new_n705));
  NAND2_X1  g0505(.A1(G20), .A2(G179), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT93), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(G190), .A3(G200), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n309), .A3(G200), .ZN(new_n709));
  XOR2_X1   g0509(.A(KEYINPUT33), .B(G317), .Z(new_n710));
  OAI221_X1 g0510(.A(new_n704), .B1(new_n705), .B2(new_n708), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n309), .A2(G200), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n707), .A2(KEYINPUT94), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT94), .B1(new_n707), .B2(new_n712), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n711), .B1(G322), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G190), .A2(G200), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n707), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n697), .A2(new_n717), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n718), .A2(G311), .B1(G329), .B2(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n697), .A2(G190), .A3(G200), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n299), .A2(new_n301), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n712), .A2(new_n550), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI221_X1 g0527(.A(new_n722), .B1(new_n581), .B2(new_n723), .C1(new_n724), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n718), .A2(KEYINPUT95), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n707), .A2(new_n717), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n733), .A2(G77), .B1(G58), .B2(new_n715), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT96), .Z(new_n735));
  INV_X1    g0535(.A(new_n723), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G87), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n727), .A2(new_n214), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n451), .B1(new_n708), .B2(new_n222), .C1(new_n702), .C2(new_n218), .ZN(new_n739));
  INV_X1    g0539(.A(new_n709), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n738), .B(new_n739), .C1(G68), .C2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT98), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n720), .A2(G159), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n735), .A2(new_n737), .A3(new_n741), .A4(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n696), .B1(new_n728), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n689), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n747), .A2(new_n692), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n248), .A2(G45), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n654), .A2(new_n451), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(G45), .C2(new_n234), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n209), .A2(G355), .A3(new_n451), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n756), .B(new_n757), .C1(G116), .C2(new_n209), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT92), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n750), .A2(new_n695), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n694), .B1(new_n753), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(G396));
  INV_X1    g0563(.A(new_n708), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n733), .A2(G116), .B1(G303), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n766), .B2(new_n709), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT100), .Z(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(G311), .B2(new_n720), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n702), .A2(new_n212), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n738), .B1(new_n715), .B2(G294), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n451), .B1(new_n736), .B2(G107), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n769), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n702), .A2(new_n343), .B1(new_n227), .B2(new_n727), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n715), .A2(G143), .B1(G150), .B2(new_n740), .ZN(new_n776));
  INV_X1    g0576(.A(G137), .ZN(new_n777));
  INV_X1    g0577(.A(new_n733), .ZN(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n776), .B1(new_n777), .B2(new_n708), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT34), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n314), .B(new_n775), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n720), .A2(G132), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n780), .A2(new_n781), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n736), .A2(G50), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n774), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n695), .A2(new_n748), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n787), .A2(new_n695), .B1(new_n224), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n479), .A2(new_n634), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n484), .B2(new_n486), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n481), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n613), .A2(new_n635), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT101), .ZN(new_n794));
  AND3_X1   g0594(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(new_n792), .B2(new_n793), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n748), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n789), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n693), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT102), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n792), .A2(new_n793), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(KEYINPUT101), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n608), .A2(new_n805), .A3(new_n635), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n805), .B1(new_n608), .B2(new_n635), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n809), .A2(new_n646), .A3(new_n683), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n684), .B1(new_n807), .B2(new_n808), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n800), .B(new_n801), .C1(new_n812), .C2(new_n693), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n693), .B1(new_n810), .B2(new_n811), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n692), .B1(new_n789), .B2(new_n798), .ZN(new_n815));
  OAI21_X1  g0615(.A(KEYINPUT102), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n813), .A2(new_n816), .ZN(G384));
  INV_X1    g0617(.A(KEYINPUT38), .ZN(new_n818));
  AND3_X1   g0618(.A1(new_n321), .A2(new_n330), .A3(new_n323), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n331), .ZN(new_n820));
  INV_X1    g0620(.A(new_n317), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n335), .A2(KEYINPUT72), .A3(KEYINPUT7), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n340), .B1(new_n339), .B2(new_n316), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n820), .B1(new_n824), .B2(G68), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n344), .B(new_n266), .C1(new_n825), .C2(new_n327), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n354), .ZN(new_n827));
  INV_X1    g0627(.A(new_n632), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n382), .B2(new_n390), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n329), .A2(new_n344), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n831), .A2(new_n353), .B1(new_n373), .B2(new_n828), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT37), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n832), .A2(new_n833), .A3(new_n386), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n827), .A2(new_n373), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n835), .A2(new_n829), .A3(new_n386), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n834), .B1(KEYINPUT37), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n818), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n313), .B1(new_n825), .B2(KEYINPUT16), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n334), .B1(new_n342), .B2(new_n343), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n328), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n353), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n386), .B1(new_n842), .B2(new_n632), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n377), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT37), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n832), .A2(new_n833), .A3(new_n386), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n381), .A2(new_n379), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n616), .B1(new_n848), .B2(new_n375), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(KEYINPUT38), .C1(new_n849), .C2(new_n829), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n838), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n427), .A2(new_n634), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n428), .A2(new_n433), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT103), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT103), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n428), .A2(new_n433), .A3(new_n855), .A4(new_n852), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n417), .A2(new_n427), .A3(new_n634), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n679), .A2(KEYINPUT31), .A3(new_n634), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n859), .A2(new_n680), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n797), .B1(new_n860), .B2(new_n664), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n851), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT40), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n683), .A2(new_n805), .A3(new_n858), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n355), .A2(new_n828), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n390), .B2(new_n612), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n833), .B1(new_n832), .B2(new_n386), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n834), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n818), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n863), .B1(new_n850), .B2(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n862), .A2(new_n863), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT104), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n492), .A2(new_n683), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n646), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n623), .A2(new_n625), .B1(new_n492), .B2(new_n662), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n850), .A2(new_n869), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n428), .A2(new_n634), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n838), .A2(new_n850), .A3(KEYINPUT39), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n854), .A2(new_n856), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n793), .A2(new_n806), .B1(new_n883), .B2(new_n857), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n851), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n619), .A2(new_n632), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n882), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n876), .B(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n889), .A2(KEYINPUT105), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(KEYINPUT105), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n875), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n892), .B1(new_n205), .B2(new_n628), .C1(new_n890), .C2(new_n875), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n572), .B1(new_n516), .B2(KEYINPUT35), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n894), .B(new_n233), .C1(KEYINPUT35), .C2(new_n516), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT36), .ZN(new_n896));
  OAI21_X1  g0696(.A(G77), .B1(new_n227), .B2(new_n343), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n897), .A2(new_n234), .B1(G50), .B2(new_n343), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(G1), .A3(new_n271), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n893), .A2(new_n896), .A3(new_n899), .ZN(G367));
  NAND2_X1  g0700(.A1(new_n703), .A2(G77), .ZN(new_n901));
  INV_X1    g0701(.A(G143), .ZN(new_n902));
  OAI221_X1 g0702(.A(new_n901), .B1(new_n902), .B2(new_n708), .C1(new_n778), .C2(new_n222), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n726), .A2(G68), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n904), .B1(new_n227), .B2(new_n723), .C1(new_n777), .C2(new_n719), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n903), .A2(new_n314), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n715), .ZN(new_n907));
  OAI221_X1 g0707(.A(new_n906), .B1(new_n438), .B2(new_n907), .C1(new_n779), .C2(new_n709), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n715), .A2(G303), .B1(G311), .B2(new_n764), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT109), .ZN(new_n910));
  OAI221_X1 g0710(.A(new_n314), .B1(new_n218), .B2(new_n727), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n702), .A2(new_n214), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT110), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n736), .A2(KEYINPUT46), .A3(G116), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT46), .B1(new_n736), .B2(G116), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n909), .A2(new_n910), .B1(G317), .B2(new_n720), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n918), .B(new_n919), .C1(new_n766), .C2(new_n778), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n709), .A2(new_n724), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n908), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT47), .Z(new_n923));
  NOR2_X1   g0723(.A1(new_n923), .A2(new_n696), .ZN(new_n924));
  INV_X1    g0724(.A(new_n755), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n760), .B1(new_n209), .B2(new_n543), .C1(new_n244), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n544), .A2(new_n546), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n634), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n554), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n553), .A2(new_n928), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n693), .B(new_n926), .C1(new_n931), .C2(new_n751), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n924), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n691), .A2(G1), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n600), .A2(new_n555), .A3(new_n634), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n936), .A2(KEYINPUT107), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n526), .B(new_n566), .C1(new_n523), .C2(new_n635), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(KEYINPUT107), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n652), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT44), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n652), .A2(new_n940), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT45), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n943), .A2(new_n945), .A3(new_n650), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n650), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n641), .B(new_n651), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(new_n647), .Z(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(new_n685), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT108), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n948), .A2(KEYINPUT108), .A3(new_n951), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n685), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n655), .B(KEYINPUT41), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n935), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n649), .A2(new_n940), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT106), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n641), .A2(new_n651), .A3(new_n940), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT42), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n940), .A2(new_n570), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n634), .B1(new_n967), .B2(new_n566), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n966), .A2(new_n969), .B1(KEYINPUT43), .B2(new_n931), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n963), .A2(new_n964), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n971), .B1(new_n963), .B2(new_n964), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n933), .B1(new_n958), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(G387));
  INV_X1    g0777(.A(new_n657), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n209), .A3(new_n451), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(G107), .B2(new_n209), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT111), .Z(new_n981));
  NOR3_X1   g0781(.A1(new_n346), .A2(KEYINPUT50), .A3(G50), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n978), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(G68), .A2(G77), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT50), .B1(new_n346), .B2(G50), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n983), .A2(new_n533), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n755), .B(new_n986), .C1(new_n240), .C2(new_n533), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n692), .B1(new_n988), .B2(new_n760), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT112), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n736), .A2(G77), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n438), .B2(new_n719), .C1(new_n907), .C2(new_n222), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n314), .B(new_n992), .C1(G159), .C2(new_n764), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n727), .A2(new_n543), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n994), .B(new_n912), .C1(new_n347), .C2(new_n740), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n993), .B(new_n995), .C1(new_n343), .C2(new_n730), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT113), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n715), .A2(G317), .B1(G311), .B2(new_n740), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n764), .A2(G322), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n778), .C2(new_n581), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT48), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n766), .B2(new_n727), .C1(new_n724), .C2(new_n723), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT49), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n314), .B1(new_n719), .B2(new_n705), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n703), .B2(G116), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n997), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n990), .B1(new_n641), .B2(new_n751), .C1(new_n1006), .C2(new_n696), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n950), .A2(new_n685), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n655), .B(KEYINPUT114), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n950), .B2(new_n685), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1007), .B1(new_n935), .B2(new_n950), .C1(new_n1008), .C2(new_n1011), .ZN(G393));
  OAI221_X1 g0812(.A(new_n760), .B1(new_n214), .B2(new_n209), .C1(new_n925), .C2(new_n251), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n940), .B2(new_n751), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n715), .A2(G311), .B1(G317), .B2(new_n764), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT52), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G107), .B2(new_n703), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n740), .A2(G303), .B1(G116), .B2(new_n726), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT115), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n720), .A2(G322), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n314), .B1(new_n298), .B2(new_n730), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G283), .B2(new_n736), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n727), .A2(new_n224), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n715), .A2(G159), .B1(G150), .B2(new_n764), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(KEYINPUT51), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n347), .B2(new_n733), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n451), .B1(new_n343), .B2(new_n723), .C1(new_n709), .C2(new_n222), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n770), .B(new_n1029), .C1(new_n1026), .C2(KEYINPUT51), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1028), .B(new_n1030), .C1(new_n902), .C2(new_n719), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1024), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n692), .B(new_n1014), .C1(new_n695), .C2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n948), .B2(new_n934), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n954), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n1035), .A2(new_n952), .B1(new_n951), .B2(new_n948), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1034), .B1(new_n1036), .B2(new_n1009), .ZN(G390));
  OAI211_X1 g0837(.A(new_n879), .B(new_n881), .C1(new_n884), .C2(new_n880), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n861), .A2(G330), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n858), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n806), .A2(new_n793), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n858), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n880), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1042), .A2(new_n850), .A3(new_n1043), .A4(new_n869), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n1038), .A2(new_n1040), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n861), .A2(new_n646), .A3(new_n858), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n858), .B1(new_n806), .B2(new_n793), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n806), .A2(new_n793), .A3(new_n858), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n1039), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n861), .A2(new_n646), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1051), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n1049), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n490), .A2(new_n491), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n435), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1057), .A2(G330), .A3(new_n1058), .A4(new_n683), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n876), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1010), .B1(new_n1048), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n1048), .B2(new_n1060), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n788), .A2(new_n346), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n879), .A2(new_n881), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n748), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n736), .A2(G150), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT53), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n314), .B1(new_n715), .B2(G132), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n222), .B2(new_n702), .ZN(new_n1071));
  XOR2_X1   g0871(.A(KEYINPUT54), .B(G143), .Z(new_n1072));
  AOI211_X1 g0872(.A(new_n1069), .B(new_n1071), .C1(new_n733), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n720), .A2(G125), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n726), .A2(G159), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G128), .A2(new_n764), .B1(new_n740), .B2(G137), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n702), .A2(new_n343), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1025), .B(new_n1078), .C1(new_n733), .C2(G97), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n740), .A2(G107), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n715), .A2(G116), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n737), .B1(new_n708), .B2(new_n766), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n451), .B(new_n1082), .C1(G294), .C2(new_n720), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n696), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  OR3_X1    g0885(.A1(new_n1067), .A2(new_n692), .A3(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1048), .A2(new_n935), .B1(new_n1064), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1062), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(G378));
  NAND2_X1  g0889(.A1(new_n448), .A2(new_n828), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n466), .A2(new_n483), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1092), .B1(new_n466), .B2(new_n483), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n466), .A2(new_n483), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n1091), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1090), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n1099), .A3(new_n1093), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n748), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n222), .B1(new_n253), .B2(G41), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n715), .A2(G128), .B1(G150), .B2(new_n726), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n736), .A2(new_n1072), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT116), .Z(new_n1106));
  AOI22_X1  g0906(.A1(new_n740), .A2(G132), .B1(new_n718), .B2(G137), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G125), .B2(new_n764), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT59), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n703), .A2(G159), .ZN(new_n1112));
  AOI21_X1  g0912(.A(G33), .B1(new_n720), .B2(G124), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1111), .A2(new_n282), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1103), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n715), .A2(G107), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n740), .A2(G97), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1117), .A2(new_n314), .A3(new_n991), .A4(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n764), .A2(G116), .B1(G68), .B2(new_n726), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n766), .B2(new_n719), .C1(new_n543), .C2(new_n730), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n702), .A2(new_n227), .ZN(new_n1122));
  NOR4_X1   g0922(.A1(new_n1119), .A2(new_n1121), .A3(G41), .A4(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT58), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n695), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n788), .A2(new_n222), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1102), .A2(new_n693), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n887), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1101), .B1(new_n871), .B2(G330), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n838), .A2(new_n850), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n683), .A2(new_n805), .A3(new_n858), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n863), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n864), .A2(new_n870), .ZN(new_n1134));
  AND4_X1   g0934(.A1(G330), .A2(new_n1133), .A3(new_n1134), .A4(new_n1101), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1129), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT118), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(KEYINPUT118), .B(new_n1129), .C1(new_n1130), .C2(new_n1135), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1133), .A2(new_n1134), .A3(G330), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1101), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n871), .A2(G330), .A3(new_n1101), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n887), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT117), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1142), .A2(new_n1143), .A3(KEYINPUT117), .A4(new_n887), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1138), .A2(new_n1139), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1128), .B1(new_n1148), .B2(new_n934), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n492), .A2(new_n662), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n626), .A2(new_n1150), .A3(new_n1059), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1056), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1048), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT57), .B1(new_n1148), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1136), .A2(new_n1144), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(KEYINPUT57), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1010), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1149), .B1(new_n1155), .B2(new_n1158), .ZN(G375));
  AOI21_X1  g0959(.A(new_n1122), .B1(new_n740), .B2(new_n1072), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n764), .A2(G132), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT121), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G150), .B2(new_n718), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n726), .A2(G50), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n720), .A2(G128), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n907), .A2(new_n777), .B1(new_n779), .B2(new_n723), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n451), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n733), .A2(G107), .B1(G294), .B2(new_n764), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n572), .B2(new_n709), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT119), .Z(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(new_n994), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n715), .A2(G283), .B1(G303), .B2(new_n720), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n214), .C2(new_n723), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n901), .A2(new_n314), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT120), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1171), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n695), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n693), .C1(new_n749), .C2(new_n858), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n343), .B2(new_n788), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n934), .B2(new_n1056), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n956), .B1(new_n1152), .B2(new_n1056), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1060), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(G381));
  OR2_X1    g0987(.A1(G387), .A2(G381), .ZN(new_n1188));
  OR2_X1    g0988(.A1(G393), .A2(G396), .ZN(new_n1189));
  OR2_X1    g0989(.A1(G390), .A2(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(G375), .A2(G378), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1188), .A2(G384), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(G407));
  INV_X1    g0993(.A(KEYINPUT122), .ZN(new_n1194));
  OAI21_X1  g0994(.A(G213), .B1(new_n1191), .B2(G343), .ZN(new_n1195));
  OR3_X1    g0995(.A1(new_n1192), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1194), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(G409));
  NAND2_X1  g0998(.A1(G375), .A2(G378), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n633), .A2(G213), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1156), .A2(new_n934), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1148), .A2(new_n956), .A3(new_n1154), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1088), .A2(new_n1127), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n813), .A2(new_n816), .A3(KEYINPUT123), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT123), .B1(new_n813), .B2(new_n816), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1151), .A2(new_n1153), .A3(KEYINPUT60), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(new_n1010), .A3(new_n1060), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT60), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1184), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1184), .B(new_n1206), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n633), .A2(G213), .A3(G2897), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1214), .B(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1204), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT61), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT125), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT125), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1220), .B(KEYINPUT61), .C1(new_n1204), .C2(new_n1216), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT62), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1199), .A2(new_n1200), .A3(new_n1203), .A4(new_n1214), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT126), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1222), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1219), .A2(new_n1221), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT127), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(G393), .B(new_n762), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT124), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n976), .A2(new_n1230), .A3(G390), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n976), .A2(G390), .A3(new_n1229), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n933), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n686), .B1(new_n1035), .B2(new_n952), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n934), .B1(new_n1234), .B2(new_n956), .ZN(new_n1235));
  OAI211_X1 g1035(.A(G390), .B(new_n1233), .C1(new_n1235), .C2(new_n974), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1230), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n976), .A2(G390), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1231), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT127), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n1226), .B2(new_n1225), .C1(new_n1219), .C2(new_n1221), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1228), .A2(new_n1241), .A3(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1241), .A2(KEYINPUT61), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1217), .A2(KEYINPUT63), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1223), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT63), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1245), .B(new_n1247), .C1(new_n1248), .C2(new_n1223), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(new_n1249), .ZN(G405));
  NAND2_X1  g1050(.A1(new_n1191), .A2(new_n1199), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1241), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1239), .B1(new_n1237), .B2(new_n1232), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1191), .B(new_n1199), .C1(new_n1253), .C2(new_n1231), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1214), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1252), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1255), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(G402));
endmodule


