//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  NOR2_X1   g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT14), .Z(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT95), .B(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G29gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n207), .A2(KEYINPUT97), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT96), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n207), .A2(KEYINPUT97), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n215), .B(new_n205), .C1(new_n211), .C2(KEYINPUT96), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n209), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT17), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT98), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT98), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(new_n221), .A3(new_n218), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(G1gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G1gat), .B2(new_n224), .ZN(new_n227));
  INV_X1    g026(.A(G8gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n217), .A2(new_n218), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n223), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT99), .ZN(new_n233));
  INV_X1    g032(.A(new_n229), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n217), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n231), .A2(KEYINPUT18), .A3(new_n233), .A4(new_n235), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n234), .B(new_n217), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n233), .B(KEYINPUT13), .Z(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(G169gat), .B(G197gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT94), .B(KEYINPUT11), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT12), .Z(new_n249));
  NAND2_X1  g048(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n249), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n238), .A2(new_n239), .A3(new_n242), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G78gat), .B(G106gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT31), .B(G50gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  INV_X1    g056(.A(G141gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT79), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT79), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G141gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n261), .A3(G148gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT80), .ZN(new_n263));
  INV_X1    g062(.A(G148gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(G141gat), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269));
  INV_X1    g068(.A(G155gat), .ZN(new_n270));
  INV_X1    g069(.A(G162gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n269), .B1(new_n272), .B2(KEYINPUT2), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT2), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(G141gat), .B2(G148gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(new_n269), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT78), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n258), .A2(new_n264), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(new_n275), .A3(new_n277), .ZN(new_n284));
  INV_X1    g083(.A(new_n269), .ZN(new_n285));
  NOR2_X1   g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT78), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n274), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT22), .ZN(new_n290));
  XOR2_X1   g089(.A(KEYINPUT74), .B(G211gat), .Z(new_n291));
  INV_X1    g090(.A(G218gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294));
  XOR2_X1   g093(.A(G197gat), .B(G204gat), .Z(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n294), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT74), .B(G211gat), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT22), .B1(new_n299), .B2(G218gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n300), .B2(new_n295), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT29), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n289), .B1(new_n302), .B2(KEYINPUT3), .ZN(new_n303));
  NAND2_X1  g102(.A1(G228gat), .A2(G233gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n297), .A2(new_n301), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT3), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n274), .B(new_n310), .C1(new_n282), .C2(new_n288), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT81), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n281), .B1(new_n279), .B2(new_n280), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n284), .A2(new_n287), .A3(KEYINPUT78), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n314), .A2(new_n315), .B1(new_n268), .B2(new_n273), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(KEYINPUT81), .A3(new_n310), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT83), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n309), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI211_X1 g119(.A(KEYINPUT83), .B(KEYINPUT29), .C1(new_n313), .C2(new_n317), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n307), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G22gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n294), .B1(new_n293), .B2(new_n296), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n324), .B2(KEYINPUT82), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT82), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n297), .A2(new_n326), .A3(new_n301), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT3), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n318), .A2(new_n308), .B1(new_n328), .B2(new_n316), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n304), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n322), .A2(new_n323), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n323), .B1(new_n322), .B2(new_n330), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n257), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT84), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(KEYINPUT84), .B(new_n257), .C1(new_n331), .C2(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT86), .ZN(new_n338));
  AOI211_X1 g137(.A(KEYINPUT85), .B(new_n323), .C1(new_n322), .C2(new_n330), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n330), .ZN(new_n340));
  INV_X1    g139(.A(new_n257), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n311), .A2(new_n312), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT81), .B1(new_n316), .B2(new_n310), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n308), .B1(new_n347), .B2(KEYINPUT83), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n318), .A2(new_n319), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n306), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n325), .A2(new_n327), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n289), .B1(new_n351), .B2(KEYINPUT3), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n309), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n305), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(G22gat), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT85), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n338), .B1(new_n343), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT85), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n358), .B(G22gat), .C1(new_n350), .C2(new_n354), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(new_n341), .A3(new_n340), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n332), .A2(new_n358), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n360), .A2(KEYINPUT86), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n337), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT87), .ZN(new_n364));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(G183gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT27), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G183gat), .ZN(new_n369));
  INV_X1    g168(.A(G190gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT27), .B(G183gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(KEYINPUT28), .A3(new_n370), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT26), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n379), .A2(new_n382), .B1(G183gat), .B2(G190gat), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT66), .ZN(new_n385));
  NAND2_X1  g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n378), .B1(new_n386), .B2(KEYINPUT24), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n366), .A2(G190gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n370), .A2(G183gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n387), .B1(new_n390), .B2(KEYINPUT24), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n380), .B2(KEYINPUT65), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT65), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n394), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT64), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT66), .B1(new_n391), .B2(new_n396), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT25), .ZN(new_n399));
  OAI22_X1  g198(.A1(new_n385), .A2(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n391), .A2(new_n396), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT64), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(KEYINPUT66), .A3(KEYINPUT25), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n384), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n365), .B1(new_n405), .B2(KEYINPUT29), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT75), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n400), .A2(new_n404), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n376), .A2(KEYINPUT67), .A3(new_n383), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT67), .B1(new_n376), .B2(new_n383), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n365), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n415), .B(new_n365), .C1(new_n405), .C2(KEYINPUT29), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n407), .A2(new_n308), .A3(new_n414), .A4(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n413), .A2(KEYINPUT29), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n412), .A2(new_n418), .B1(new_n405), .B2(new_n413), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n309), .ZN(new_n420));
  XOR2_X1   g219(.A(G8gat), .B(G36gat), .Z(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT76), .ZN(new_n422));
  XNOR2_X1  g221(.A(G64gat), .B(G92gat), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n422), .B(new_n423), .Z(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n417), .A2(new_n420), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT30), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT30), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n417), .A2(new_n428), .A3(new_n420), .A4(new_n425), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431));
  NOR2_X1   g230(.A1(G127gat), .A2(G134gat), .ZN(new_n432));
  XOR2_X1   g231(.A(KEYINPUT68), .B(G127gat), .Z(new_n433));
  AOI21_X1  g232(.A(new_n432), .B1(new_n433), .B2(G134gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(G113gat), .B(G120gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT69), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT1), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n435), .A2(KEYINPUT69), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n434), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(G120gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G113gat), .ZN(new_n442));
  XOR2_X1   g241(.A(KEYINPUT70), .B(G113gat), .Z(new_n443));
  OAI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(new_n441), .ZN(new_n444));
  INV_X1    g243(.A(new_n432), .ZN(new_n445));
  NAND2_X1  g244(.A1(G127gat), .A2(G134gat), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT1), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n440), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n431), .B1(new_n449), .B2(new_n289), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT1), .B1(new_n435), .B2(KEYINPUT69), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(KEYINPUT69), .B2(new_n435), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n452), .A2(new_n434), .B1(new_n444), .B2(new_n447), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(KEYINPUT4), .A3(new_n316), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI221_X1 g255(.A(new_n449), .B1(new_n310), .B2(new_n316), .C1(new_n345), .C2(new_n346), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT5), .ZN(new_n458));
  NAND2_X1  g257(.A1(G225gat), .A2(G233gat), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n449), .B1(new_n310), .B2(new_n316), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n313), .B2(new_n317), .ZN(new_n462));
  INV_X1    g261(.A(new_n459), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n462), .A2(new_n463), .A3(new_n455), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n289), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n453), .A2(new_n316), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n463), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT5), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n460), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G1gat), .B(G29gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(KEYINPUT0), .ZN(new_n472));
  XNOR2_X1  g271(.A(G57gat), .B(G85gat), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n472), .B(new_n473), .Z(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n470), .A2(KEYINPUT6), .A3(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n460), .B(new_n474), .C1(new_n464), .C2(new_n469), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(KEYINPUT5), .A3(new_n468), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n474), .B1(new_n481), .B2(new_n460), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n476), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT77), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n417), .A2(new_n420), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n484), .B1(new_n485), .B2(new_n424), .ZN(new_n486));
  AOI211_X1 g285(.A(KEYINPUT77), .B(new_n425), .C1(new_n417), .C2(new_n420), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n430), .B(new_n483), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT86), .B1(new_n360), .B2(new_n361), .ZN(new_n489));
  INV_X1    g288(.A(new_n342), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n490), .A2(new_n356), .A3(new_n338), .A4(new_n359), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n337), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n364), .A2(new_n488), .A3(new_n494), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n408), .A2(new_n449), .A3(new_n411), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n449), .B1(new_n408), .B2(new_n411), .ZN(new_n497));
  INV_X1    g296(.A(G227gat), .ZN(new_n498));
  INV_X1    g297(.A(G233gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n496), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT32), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G15gat), .B(G43gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT72), .ZN(new_n506));
  XNOR2_X1  g305(.A(G71gat), .B(G99gat), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n506), .B(new_n507), .Z(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT33), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT73), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n509), .B1(new_n502), .B2(new_n503), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT71), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n412), .A2(new_n453), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n408), .A2(new_n449), .A3(new_n411), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n500), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT33), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n514), .A3(new_n518), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n512), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT71), .B1(new_n502), .B2(KEYINPUT33), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n508), .B1(new_n517), .B2(KEYINPUT32), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n512), .A4(new_n521), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n511), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n501), .B1(new_n496), .B2(new_n497), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT34), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n523), .A2(new_n521), .A3(new_n524), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT73), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n525), .ZN(new_n533));
  INV_X1    g332(.A(new_n529), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n534), .A3(new_n511), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(KEYINPUT36), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT36), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n534), .B1(new_n533), .B2(new_n511), .ZN(new_n538));
  INV_X1    g337(.A(new_n511), .ZN(new_n539));
  AOI211_X1 g338(.A(new_n529), .B(new_n539), .C1(new_n532), .C2(new_n525), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n537), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT88), .B1(new_n495), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n426), .A2(KEYINPUT30), .ZN(new_n544));
  INV_X1    g343(.A(new_n429), .ZN(new_n545));
  OAI22_X1  g344(.A1(new_n544), .A2(new_n545), .B1(new_n486), .B2(new_n487), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT39), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n547), .B(new_n463), .C1(new_n462), .C2(new_n455), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n459), .B1(new_n456), .B2(new_n457), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT89), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n467), .B2(new_n463), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT89), .A4(new_n459), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(KEYINPUT39), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n474), .B(new_n548), .C1(new_n549), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT40), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n463), .B1(new_n462), .B2(new_n455), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n557), .A2(KEYINPUT39), .A3(new_n551), .A4(new_n552), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n558), .A2(KEYINPUT40), .A3(new_n474), .A4(new_n548), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT90), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n470), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n481), .A2(KEYINPUT90), .A3(new_n460), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n474), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n492), .A2(new_n337), .B1(new_n546), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT37), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n417), .A2(new_n567), .A3(new_n420), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n424), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n417), .B2(new_n420), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT38), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT93), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT93), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n573), .B(KEYINPUT38), .C1(new_n569), .C2(new_n570), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n407), .A2(new_n309), .A3(new_n414), .A4(new_n416), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n567), .B1(new_n419), .B2(new_n308), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT38), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(new_n424), .A3(new_n568), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n578), .A2(KEYINPUT92), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(KEYINPUT92), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n572), .B(new_n574), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n563), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n475), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT91), .ZN(new_n584));
  INV_X1    g383(.A(new_n479), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT91), .B1(new_n564), .B2(new_n479), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n586), .A2(new_n587), .A3(new_n476), .A4(new_n426), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n566), .B1(new_n581), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n543), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n495), .A2(new_n542), .A3(KEYINPUT88), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n488), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n363), .A2(new_n530), .A3(new_n594), .A4(new_n535), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT35), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n479), .B1(new_n582), .B2(new_n475), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n597), .A2(new_n584), .B1(KEYINPUT6), .B2(new_n482), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT35), .B1(new_n598), .B2(new_n587), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n538), .A2(new_n540), .ZN(new_n600));
  INV_X1    g399(.A(new_n546), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .A4(new_n363), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n254), .B1(new_n593), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT101), .B(G85gat), .Z(new_n606));
  INV_X1    g405(.A(G92gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G85gat), .A2(G92gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT7), .ZN(new_n610));
  INV_X1    g409(.A(G99gat), .ZN(new_n611));
  INV_X1    g410(.A(G106gat), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT8), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G99gat), .B(G106gat), .Z(new_n615));
  OR3_X1    g414(.A1(new_n614), .A2(KEYINPUT102), .A3(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n615), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(KEYINPUT102), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n223), .A2(new_n230), .A3(new_n616), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n616), .ZN(new_n621));
  INV_X1    g420(.A(G232gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(new_n499), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n621), .A2(new_n217), .B1(KEYINPUT41), .B2(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(KEYINPUT103), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n605), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(KEYINPUT103), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632));
  INV_X1    g431(.A(new_n626), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n620), .A2(new_n624), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n605), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n628), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n631), .B1(new_n628), .B2(new_n636), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT9), .ZN(new_n640));
  INV_X1    g439(.A(G71gat), .ZN(new_n641));
  INV_X1    g440(.A(G78gat), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n643), .A2(KEYINPUT100), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(KEYINPUT100), .ZN(new_n645));
  XOR2_X1   g444(.A(G57gat), .B(G64gat), .Z(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(G71gat), .B(G78gat), .Z(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n648), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n644), .A2(new_n650), .A3(new_n645), .A4(new_n646), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT21), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G231gat), .A2(G233gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G127gat), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n229), .B1(new_n652), .B2(new_n653), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n270), .ZN(new_n661));
  XOR2_X1   g460(.A(G183gat), .B(G211gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n659), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n639), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(G230gat), .A2(G233gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT104), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  INV_X1    g471(.A(new_n652), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n619), .B2(new_n616), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n652), .B1(new_n617), .B2(new_n618), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n621), .A2(KEYINPUT10), .A3(new_n673), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n671), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n674), .A2(new_n670), .A3(new_n675), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n669), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT105), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n682), .A2(new_n670), .ZN(new_n683));
  OR3_X1    g482(.A1(new_n683), .A2(new_n669), .A3(new_n679), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n665), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n604), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT106), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n604), .A2(new_n691), .A3(new_n688), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n483), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  AND3_X1   g496(.A1(new_n693), .A2(new_n546), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n228), .B1(new_n693), .B2(new_n546), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT42), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(KEYINPUT42), .B2(new_n698), .ZN(G1325gat));
  INV_X1    g500(.A(G15gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n693), .A2(new_n702), .A3(new_n600), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n542), .B1(new_n690), .B2(new_n692), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n702), .ZN(G1326gat));
  NAND2_X1  g504(.A1(new_n364), .A2(new_n494), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n692), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n691), .B1(new_n604), .B2(new_n688), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT107), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n693), .A2(new_n712), .A3(new_n707), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT43), .B(G22gat), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n711), .B2(new_n713), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(G1327gat));
  INV_X1    g516(.A(G29gat), .ZN(new_n718));
  INV_X1    g517(.A(new_n664), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n685), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n639), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n604), .A2(new_n718), .A3(new_n694), .A4(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n723), .A2(KEYINPUT108), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(KEYINPUT108), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n724), .B2(new_n725), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n720), .A2(new_n253), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n593), .A2(new_n603), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n639), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT44), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n495), .A2(new_n542), .A3(new_n589), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n603), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n637), .B2(new_n638), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n628), .A2(new_n636), .ZN(new_n737));
  INV_X1    g536(.A(new_n631), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n628), .A2(new_n631), .A3(new_n636), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(KEYINPUT109), .A3(new_n740), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n729), .B1(new_n732), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n746), .A2(new_n694), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n727), .B(new_n728), .C1(new_n718), .C2(new_n747), .ZN(G1328gat));
  INV_X1    g547(.A(new_n206), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n746), .B2(new_n546), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n604), .A2(new_n749), .A3(new_n546), .A4(new_n722), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT46), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753));
  OR3_X1    g552(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n750), .B2(new_n752), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1329gat));
  INV_X1    g555(.A(G43gat), .ZN(new_n757));
  INV_X1    g556(.A(new_n542), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(new_n746), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n604), .ZN(new_n760));
  INV_X1    g559(.A(new_n600), .ZN(new_n761));
  NOR4_X1   g560(.A1(new_n760), .A2(G43gat), .A3(new_n761), .A4(new_n721), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n766), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n762), .B2(new_n759), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1330gat));
  NOR4_X1   g569(.A1(new_n760), .A2(G50gat), .A3(new_n706), .A4(new_n721), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n746), .A2(new_n707), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(G50gat), .ZN(new_n773));
  INV_X1    g572(.A(G50gat), .ZN(new_n774));
  INV_X1    g573(.A(new_n363), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n746), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT48), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n771), .A2(new_n777), .ZN(new_n778));
  OAI22_X1  g577(.A1(new_n773), .A2(KEYINPUT48), .B1(new_n776), .B2(new_n778), .ZN(G1331gat));
  NOR4_X1   g578(.A1(new_n664), .A2(new_n639), .A3(new_n686), .A4(new_n253), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n734), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n694), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g583(.A1(new_n781), .A2(new_n601), .ZN(new_n785));
  NOR2_X1   g584(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n786));
  AND2_X1   g585(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n785), .B2(new_n786), .ZN(G1333gat));
  NOR3_X1   g588(.A1(new_n781), .A2(G71gat), .A3(new_n761), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n782), .A2(new_n758), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(G71gat), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g592(.A1(new_n781), .A2(new_n706), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(new_n642), .ZN(G1335gat));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n495), .A2(new_n542), .A3(new_n589), .ZN(new_n797));
  AND4_X1   g596(.A1(new_n601), .A2(new_n363), .A3(new_n530), .A4(new_n535), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n798), .A2(new_n599), .B1(KEYINPUT35), .B2(new_n595), .ZN(new_n799));
  OAI211_X1 g598(.A(KEYINPUT112), .B(new_n639), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n719), .A2(new_n253), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT112), .B1(new_n734), .B2(new_n639), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n796), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n734), .A2(new_n639), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(KEYINPUT51), .A3(new_n801), .A4(new_n800), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n686), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n694), .A3(new_n606), .ZN(new_n810));
  INV_X1    g609(.A(new_n801), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n686), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT44), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n730), .B2(new_n639), .ZN(new_n814));
  INV_X1    g613(.A(new_n745), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n483), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n810), .B1(new_n817), .B2(new_n606), .ZN(G1336gat));
  NAND3_X1  g617(.A1(new_n685), .A2(new_n607), .A3(new_n546), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n804), .B2(new_n808), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT52), .B1(new_n820), .B2(KEYINPUT113), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n546), .B(new_n812), .C1(new_n814), .C2(new_n815), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n820), .B1(new_n823), .B2(G92gat), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n825), .B(KEYINPUT52), .C1(new_n820), .C2(KEYINPUT113), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n822), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n824), .B1(new_n822), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(G1337gat));
  OAI21_X1  g628(.A(G99gat), .B1(new_n816), .B2(new_n542), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n809), .A2(new_n611), .A3(new_n600), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1338gat));
  INV_X1    g631(.A(new_n816), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n612), .B1(new_n833), .B2(new_n707), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n809), .A2(new_n612), .A3(new_n775), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT53), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(KEYINPUT115), .A3(new_n775), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n816), .B2(new_n363), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n837), .A2(G106gat), .A3(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n835), .A2(KEYINPUT53), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(G1339gat));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n668), .B1(new_n678), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n682), .B2(new_n670), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n676), .A2(new_n677), .A3(new_n671), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n845), .B2(new_n847), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n684), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n845), .A2(new_n847), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT117), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT55), .B1(new_n856), .B2(new_n844), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT118), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n850), .A2(new_n851), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(KEYINPUT55), .A3(new_n844), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .A4(new_n684), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n858), .A2(new_n253), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n233), .B1(new_n231), .B2(new_n235), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n240), .A2(new_n241), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n248), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n252), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n685), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n742), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  AND4_X1   g668(.A1(new_n742), .A2(new_n858), .A3(new_n867), .A4(new_n862), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n664), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n688), .A2(new_n872), .A3(new_n254), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT116), .B1(new_n687), .B2(new_n253), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI211_X1 g674(.A(new_n761), .B(new_n707), .C1(new_n871), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n546), .A2(new_n483), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G113gat), .B1(new_n878), .B2(new_n254), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n483), .B1(new_n871), .B2(new_n875), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n880), .A2(new_n798), .ZN(new_n881));
  INV_X1    g680(.A(new_n443), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n253), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n879), .A2(new_n883), .ZN(G1340gat));
  NOR3_X1   g683(.A1(new_n878), .A2(new_n441), .A3(new_n686), .ZN(new_n885));
  AOI21_X1  g684(.A(G120gat), .B1(new_n881), .B2(new_n685), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(G1341gat));
  OAI21_X1  g686(.A(new_n433), .B1(new_n878), .B2(new_n664), .ZN(new_n888));
  INV_X1    g687(.A(new_n433), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n881), .A2(new_n889), .A3(new_n719), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1342gat));
  INV_X1    g690(.A(G134gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n881), .A2(new_n892), .A3(new_n639), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(KEYINPUT56), .ZN(new_n894));
  INV_X1    g693(.A(new_n639), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n878), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(KEYINPUT56), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(G1343gat));
  NAND2_X1  g697(.A1(new_n542), .A2(new_n877), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n873), .A2(new_n874), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT55), .B1(new_n850), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n856), .A2(KEYINPUT119), .A3(new_n844), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n860), .A2(new_n253), .A3(new_n684), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n868), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n895), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n742), .A2(new_n858), .A3(new_n867), .A4(new_n862), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n719), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n707), .B1(new_n900), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n899), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n871), .A2(new_n875), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n775), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n253), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n259), .A2(new_n261), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT58), .B1(new_n917), .B2(KEYINPUT120), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n542), .A2(new_n775), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n546), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n880), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n921), .A2(G141gat), .A3(new_n254), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n922), .B1(new_n915), .B2(new_n916), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n918), .B(new_n923), .ZN(G1344gat));
  NAND2_X1  g723(.A1(new_n912), .A2(new_n775), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT57), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n639), .A2(new_n867), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n852), .A2(new_n857), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n719), .B1(new_n907), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n687), .A2(new_n253), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n927), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n906), .A2(new_n895), .B1(new_n929), .B2(new_n928), .ZN(new_n934));
  OAI221_X1 g733(.A(KEYINPUT122), .B1(new_n253), .B2(new_n687), .C1(new_n934), .C2(new_n719), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n706), .A2(KEYINPUT57), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n685), .B1(new_n899), .B2(KEYINPUT121), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n938), .B1(new_n899), .B2(KEYINPUT121), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n926), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n940), .A2(KEYINPUT123), .ZN(new_n941));
  OAI21_X1  g740(.A(G148gat), .B1(new_n940), .B2(KEYINPUT123), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT59), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n265), .A2(new_n266), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(KEYINPUT59), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n911), .A2(new_n914), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(new_n686), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n921), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n945), .A3(new_n685), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1345gat));
  AOI21_X1  g751(.A(G155gat), .B1(new_n950), .B2(new_n719), .ZN(new_n953));
  INV_X1    g752(.A(new_n947), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n664), .A2(new_n270), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT124), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n953), .B1(new_n954), .B2(new_n956), .ZN(G1346gat));
  AOI21_X1  g756(.A(G162gat), .B1(new_n950), .B2(new_n639), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n743), .A2(new_n271), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n954), .B2(new_n959), .ZN(G1347gat));
  AOI21_X1  g759(.A(new_n694), .B1(new_n871), .B2(new_n875), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n761), .A2(new_n775), .A3(new_n601), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(G169gat), .B1(new_n964), .B2(new_n253), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n601), .A2(new_n694), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n876), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n253), .A2(G169gat), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(G1348gat));
  INV_X1    g768(.A(G176gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n964), .A2(new_n970), .A3(new_n685), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n967), .A2(new_n685), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n972), .B2(new_n970), .ZN(G1349gat));
  AOI21_X1  g772(.A(new_n366), .B1(new_n967), .B2(new_n719), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n964), .A2(new_n374), .A3(new_n719), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g775(.A(new_n976), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g776(.A(new_n370), .B1(new_n967), .B2(new_n639), .ZN(new_n978));
  XOR2_X1   g777(.A(new_n978), .B(KEYINPUT61), .Z(new_n979));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n370), .A3(new_n742), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1351gat));
  NOR2_X1   g780(.A1(new_n919), .A2(new_n601), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n961), .A2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(G197gat), .B1(new_n984), .B2(new_n253), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n926), .A2(new_n937), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n542), .A2(new_n966), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n253), .A2(G197gat), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(G1352gat));
  NOR3_X1   g790(.A1(new_n983), .A2(G204gat), .A3(new_n686), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT62), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT125), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n994), .B1(new_n988), .B2(new_n686), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(G204gat), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n988), .A2(new_n994), .A3(new_n686), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(G1353gat));
  NAND3_X1  g797(.A1(new_n984), .A2(new_n291), .A3(new_n719), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n926), .A2(new_n719), .A3(new_n937), .A4(new_n987), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n1000), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1001));
  AOI21_X1  g800(.A(KEYINPUT63), .B1(new_n1000), .B2(G211gat), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g804(.A(KEYINPUT126), .B(new_n999), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(G1354gat));
  AOI21_X1  g806(.A(G218gat), .B1(new_n984), .B2(new_n742), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n639), .A2(G218gat), .ZN(new_n1009));
  XOR2_X1   g808(.A(new_n1009), .B(KEYINPUT127), .Z(new_n1010));
  AOI21_X1  g809(.A(new_n1008), .B1(new_n989), .B2(new_n1010), .ZN(G1355gat));
endmodule


