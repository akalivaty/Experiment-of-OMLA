//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309, new_n1310;
  OAI21_X1  g0000(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n204), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G107), .A2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(G97), .A2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR4_X1   g0024(.A1(new_n217), .A2(new_n218), .A3(new_n221), .A4(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(KEYINPUT65), .A2(G68), .ZN(new_n226));
  NAND2_X1  g0026(.A1(KEYINPUT65), .A2(G68), .ZN(new_n227));
  AND2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G238), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n212), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  OR3_X1    g0031(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(new_n201), .ZN(new_n233));
  INV_X1    g0033(.A(G50), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G1), .A2(G13), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n236), .A2(new_n211), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(new_n212), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n239), .A2(G13), .ZN(new_n240));
  OAI211_X1 g0040(.A(new_n240), .B(G250), .C1(G257), .C2(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT0), .ZN(new_n242));
  NAND3_X1  g0042(.A1(new_n231), .A2(new_n238), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G232), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT2), .B(G226), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G250), .B(G257), .Z(new_n249));
  XNOR2_X1  g0049(.A(G264), .B(G270), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G358));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  INV_X1    g0053(.A(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(KEYINPUT67), .B(G107), .Z(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(G68), .B(G77), .ZN(new_n258));
  XNOR2_X1  g0058(.A(G50), .B(G58), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XOR2_X1   g0060(.A(new_n257), .B(new_n260), .Z(G351));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n236), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n211), .A2(G33), .ZN(new_n264));
  XOR2_X1   g0064(.A(new_n264), .B(KEYINPUT71), .Z(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n219), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n228), .A2(new_n211), .B1(new_n234), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n263), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT11), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n210), .A2(KEYINPUT69), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT69), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G1), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n263), .B1(new_n275), .B2(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G68), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G13), .A3(G20), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT12), .B1(new_n278), .B2(new_n228), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT74), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n278), .A2(KEYINPUT12), .A3(G68), .ZN(new_n281));
  OR2_X1    g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n271), .A2(new_n277), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n275), .A2(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n275), .A2(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n236), .B1(G33), .B2(G41), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G238), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT68), .B(G41), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n210), .B(G274), .C1(new_n292), .C2(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G97), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n223), .A2(G1698), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(G226), .B2(G1698), .ZN(new_n296));
  INV_X1    g0096(.A(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT3), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n294), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n287), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n291), .A2(new_n293), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT13), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT13), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n291), .A2(new_n306), .A3(new_n293), .A4(new_n303), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G190), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n284), .B(new_n309), .C1(new_n310), .C2(new_n308), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n308), .A2(KEYINPUT14), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT14), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n305), .A2(new_n307), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(G169), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n313), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n311), .B1(new_n319), .B2(new_n284), .ZN(new_n320));
  OAI21_X1  g0120(.A(G20), .B1(new_n204), .B2(G50), .ZN(new_n321));
  INV_X1    g0121(.A(G150), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT70), .B(G58), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT8), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(KEYINPUT8), .B2(G58), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n321), .B1(new_n322), .B2(new_n268), .C1(new_n325), .C2(new_n265), .ZN(new_n326));
  INV_X1    g0126(.A(new_n278), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n326), .A2(new_n263), .B1(new_n234), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n276), .A2(G50), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT3), .B(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G222), .A2(G1698), .ZN(new_n332));
  INV_X1    g0132(.A(G1698), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(G223), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(new_n287), .C1(G77), .C2(new_n331), .ZN(new_n336));
  INV_X1    g0136(.A(G226), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n336), .B(new_n293), .C1(new_n289), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n312), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n338), .A2(G179), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n330), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n328), .A2(KEYINPUT9), .A3(new_n329), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT9), .B1(new_n328), .B2(new_n329), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT10), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n338), .A2(G200), .ZN(new_n348));
  INV_X1    g0148(.A(G190), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n338), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n346), .A2(new_n347), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT9), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n330), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n353), .A2(new_n348), .A3(new_n343), .A4(new_n350), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT10), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n342), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n331), .A2(G232), .A3(new_n333), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT72), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n331), .A2(G1698), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n359), .A2(new_n290), .B1(new_n207), .B2(new_n331), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n287), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n361), .B(new_n293), .C1(new_n220), .C2(new_n289), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n362), .A2(G179), .ZN(new_n363));
  XOR2_X1   g0163(.A(KEYINPUT8), .B(G58), .Z(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n267), .B1(G20), .B2(G77), .ZN(new_n365));
  XOR2_X1   g0165(.A(KEYINPUT15), .B(G87), .Z(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n264), .B2(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(new_n263), .B1(new_n219), .B2(new_n327), .ZN(new_n369));
  INV_X1    g0169(.A(new_n276), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n369), .B1(new_n219), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n362), .A2(new_n312), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n363), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n362), .B2(G200), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n349), .B2(new_n362), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n356), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n320), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n356), .A2(KEYINPUT73), .A3(new_n373), .A4(new_n375), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n325), .A2(new_n327), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n370), .B2(new_n325), .ZN(new_n381));
  NOR2_X1   g0181(.A1(G223), .A2(G1698), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n333), .A2(G226), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n301), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G87), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT78), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n287), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n285), .A2(new_n286), .A3(G232), .A4(new_n288), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n387), .A2(new_n349), .A3(new_n293), .A4(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(KEYINPUT79), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n301), .B2(new_n211), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  AOI211_X1 g0192(.A(new_n392), .B(G20), .C1(new_n298), .C2(new_n300), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT75), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n392), .B1(new_n331), .B2(G20), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n299), .A2(G33), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT7), .B(new_n211), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(KEYINPUT75), .A3(G68), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n222), .A2(KEYINPUT70), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT70), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G58), .ZN(new_n406));
  AND4_X1   g0206(.A1(new_n226), .A2(new_n404), .A3(new_n406), .A4(new_n227), .ZN(new_n407));
  OAI21_X1  g0207(.A(G20), .B1(new_n407), .B2(new_n233), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT76), .ZN(new_n409));
  INV_X1    g0209(.A(G159), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n268), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n226), .A2(new_n404), .A3(new_n406), .A4(new_n227), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n211), .B1(new_n204), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT76), .B1(new_n415), .B2(new_n411), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n403), .A2(KEYINPUT16), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n263), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n415), .A2(new_n411), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n401), .A2(new_n228), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT16), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n419), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI211_X1 g0224(.A(new_n381), .B(new_n390), .C1(new_n418), .C2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT80), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n387), .A2(new_n293), .A3(new_n388), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n310), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT79), .A3(new_n389), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n425), .A2(new_n428), .A3(new_n429), .A4(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n409), .B1(new_n408), .B2(new_n412), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n415), .A2(KEYINPUT76), .A3(new_n411), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT75), .B1(new_n401), .B2(G68), .ZN(new_n436));
  INV_X1    g0236(.A(G68), .ZN(new_n437));
  AOI211_X1 g0237(.A(new_n395), .B(new_n437), .C1(new_n397), .C2(new_n400), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n434), .A2(new_n435), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n424), .B1(new_n439), .B2(new_n423), .ZN(new_n440));
  INV_X1    g0240(.A(new_n390), .ZN(new_n441));
  INV_X1    g0241(.A(new_n381), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n440), .A2(new_n432), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n426), .A3(new_n427), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n433), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n430), .A2(G169), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n387), .A2(G179), .A3(new_n293), .A4(new_n388), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT77), .B1(new_n440), .B2(new_n442), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT77), .ZN(new_n451));
  AOI211_X1 g0251(.A(new_n451), .B(new_n381), .C1(new_n418), .C2(new_n424), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n449), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(KEYINPUT18), .B(new_n449), .C1(new_n450), .C2(new_n452), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n445), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n378), .A2(new_n379), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n298), .A2(new_n300), .A3(G250), .A4(new_n333), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n298), .A2(new_n300), .A3(G257), .A4(G1698), .ZN(new_n461));
  XOR2_X1   g0261(.A(KEYINPUT88), .B(G294), .Z(new_n462));
  OAI211_X1 g0262(.A(new_n460), .B(new_n461), .C1(new_n462), .C2(new_n297), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n287), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT89), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n275), .A2(G45), .A3(G274), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n292), .B2(KEYINPUT5), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n288), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n463), .A2(KEYINPUT89), .A3(new_n287), .ZN(new_n472));
  INV_X1    g0272(.A(new_n469), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT68), .B(G41), .Z(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(G264), .B(new_n288), .C1(new_n476), .C2(new_n286), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n466), .A2(new_n471), .A3(new_n472), .A4(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n477), .A2(new_n471), .A3(new_n464), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n478), .A2(G190), .B1(new_n479), .B2(G200), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n275), .A2(G33), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n278), .A2(new_n419), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G107), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n278), .A2(G107), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n484), .B(KEYINPUT25), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n298), .A2(new_n300), .A3(new_n211), .A4(G87), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT87), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT22), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(KEYINPUT22), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n331), .A2(new_n211), .A3(G87), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n211), .A2(G107), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n493), .B(KEYINPUT23), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT24), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n491), .A2(KEYINPUT24), .A3(new_n492), .A4(new_n494), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(new_n263), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n480), .A2(new_n483), .A3(new_n485), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n286), .A2(G250), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n287), .B1(new_n501), .B2(new_n467), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n220), .A2(G1698), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n331), .B(new_n503), .C1(G238), .C2(G1698), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G116), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n288), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G190), .ZN(new_n508));
  OAI21_X1  g0308(.A(G200), .B1(new_n502), .B2(new_n506), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT81), .B(G97), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n215), .A3(new_n207), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT19), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n211), .B1(new_n294), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n331), .A2(new_n211), .A3(G68), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n512), .B1(new_n510), .B2(new_n264), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(new_n263), .B1(new_n327), .B2(new_n367), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n482), .A2(G87), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n508), .A2(new_n509), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n507), .A2(new_n317), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(new_n263), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n327), .A2(new_n367), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n482), .A2(new_n366), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n312), .B1(new_n502), .B2(new_n506), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n521), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n520), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n478), .A2(G169), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n479), .A2(G179), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n499), .A2(new_n483), .A3(new_n485), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n500), .A2(new_n528), .A3(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n278), .A2(new_n481), .A3(G116), .A4(new_n419), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n327), .A2(new_n254), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n211), .B(new_n537), .C1(new_n510), .C2(G33), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n262), .A2(new_n236), .B1(G20), .B2(new_n254), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n538), .A2(KEYINPUT20), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT20), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n535), .B(new_n536), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G270), .B(new_n288), .C1(new_n476), .C2(new_n286), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n331), .A2(G264), .A3(G1698), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n331), .A2(G257), .A3(new_n333), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n301), .A2(G303), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n287), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n543), .A2(new_n548), .A3(new_n471), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n542), .A2(G169), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT21), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n549), .A2(new_n317), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n542), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n542), .A2(new_n549), .A3(KEYINPUT21), .A4(G169), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n549), .A2(G200), .ZN(new_n557));
  INV_X1    g0357(.A(new_n542), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT86), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n549), .A2(new_n349), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n556), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n278), .A2(G97), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT6), .B1(new_n510), .B2(G107), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT6), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G97), .A2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n208), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT82), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n566), .A2(new_n572), .A3(new_n569), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n211), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n401), .A2(G107), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n219), .B2(new_n268), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n263), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT83), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n566), .A2(new_n572), .A3(new_n569), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n572), .B1(new_n566), .B2(new_n569), .ZN(new_n580));
  OAI21_X1  g0380(.A(G20), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n401), .A2(G107), .B1(G77), .B2(new_n267), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT83), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(new_n263), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n565), .B1(new_n578), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n286), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n287), .B1(new_n587), .B2(new_n470), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n470), .A2(new_n288), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n588), .A2(G257), .B1(new_n589), .B2(new_n468), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n298), .A2(new_n300), .A3(G244), .A4(new_n333), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT84), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT4), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n331), .A2(G244), .A3(new_n333), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(KEYINPUT84), .A2(KEYINPUT4), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n537), .B1(new_n359), .B2(new_n216), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n287), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n590), .A2(G190), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g0401(.A(new_n601), .B(KEYINPUT85), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n482), .A2(G97), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n590), .A2(new_n600), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n604), .A2(new_n310), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n586), .A2(new_n602), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n565), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n584), .B1(new_n583), .B2(new_n263), .ZN(new_n608));
  AOI211_X1 g0408(.A(KEYINPUT83), .B(new_n419), .C1(new_n581), .C2(new_n582), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n607), .B(new_n603), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n604), .A2(G169), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n604), .A2(new_n317), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n534), .A2(new_n564), .A3(new_n606), .A4(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n459), .A2(new_n615), .ZN(G372));
  AND2_X1   g0416(.A1(new_n552), .A2(new_n555), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n554), .A3(new_n533), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n526), .A2(KEYINPUT90), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n521), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT90), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n621), .B(new_n312), .C1(new_n502), .C2(new_n506), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n525), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n520), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n532), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n624), .B1(new_n625), .B2(new_n480), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n606), .A2(new_n614), .A3(new_n618), .A4(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n611), .B1(new_n586), .B2(new_n603), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  INV_X1    g0429(.A(new_n623), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n526), .A2(KEYINPUT90), .B1(new_n507), .B2(new_n317), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n518), .A2(new_n509), .A3(new_n519), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(new_n508), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n628), .A2(new_n629), .A3(new_n613), .A4(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n620), .A2(new_n623), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n610), .A2(new_n528), .A3(new_n612), .A4(new_n613), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT26), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n627), .A2(new_n634), .A3(new_n636), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n458), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n440), .A2(new_n442), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(KEYINPUT18), .A3(new_n449), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n381), .B1(new_n418), .B2(new_n424), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n454), .B1(new_n643), .B2(new_n448), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n319), .A2(new_n284), .ZN(new_n646));
  INV_X1    g0446(.A(new_n373), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n311), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n645), .B1(new_n648), .B2(new_n445), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n351), .A2(new_n355), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n342), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n640), .A2(new_n651), .ZN(G369));
  INV_X1    g0452(.A(G13), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(G20), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n275), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT27), .ZN(new_n656));
  OR3_X1    g0456(.A1(new_n655), .A2(KEYINPUT91), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G213), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n655), .B2(new_n656), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT91), .B1(new_n655), .B2(new_n656), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(new_n558), .ZN(new_n664));
  MUX2_X1   g0464(.A(new_n564), .B(new_n556), .S(new_n664), .Z(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G330), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n533), .A2(new_n663), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT93), .ZN(new_n669));
  INV_X1    g0469(.A(new_n663), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n532), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT92), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n533), .A3(new_n500), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n556), .A2(new_n663), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n533), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n674), .A2(new_n677), .B1(new_n678), .B2(new_n663), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n240), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n292), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G1), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n511), .A2(G116), .ZN(new_n685));
  INV_X1    g0485(.A(new_n235), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n684), .A2(new_n685), .B1(new_n686), .B2(new_n683), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n639), .A2(new_n663), .ZN(new_n689));
  XNOR2_X1  g0489(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT96), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n637), .A2(KEYINPUT26), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n610), .A2(new_n633), .A3(new_n612), .A4(new_n613), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n635), .B1(new_n695), .B2(KEYINPUT26), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n606), .A2(new_n614), .A3(new_n626), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT97), .B1(new_n678), .B2(new_n556), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT97), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n617), .A2(new_n699), .A3(new_n533), .A4(new_n554), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n694), .B(new_n696), .C1(new_n697), .C2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .A3(new_n663), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n689), .A2(KEYINPUT96), .A3(new_n690), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n693), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT94), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n477), .A2(new_n464), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n604), .A2(new_n707), .A3(new_n507), .ZN(new_n708));
  INV_X1    g0508(.A(new_n553), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT30), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n706), .B(new_n712), .C1(new_n708), .C2(new_n709), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n604), .A2(new_n479), .ZN(new_n714));
  INV_X1    g0514(.A(new_n507), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(new_n317), .A3(new_n549), .A4(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n711), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n670), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n718), .B(KEYINPUT31), .C1(new_n615), .C2(new_n670), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n720), .A3(new_n670), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n705), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n688), .B1(new_n724), .B2(G1), .ZN(G364));
  AOI21_X1  g0525(.A(new_n210), .B1(new_n654), .B2(G45), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n682), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n667), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G330), .B2(new_n665), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G13), .A2(G33), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OR3_X1    g0532(.A1(new_n665), .A2(G20), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n240), .A2(G355), .A3(new_n331), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n260), .A2(G45), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT98), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n681), .A2(new_n331), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n686), .B2(G45), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n734), .B1(G116), .B2(new_n240), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n732), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n236), .B1(G20), .B2(new_n312), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n211), .A2(G190), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n310), .A2(G179), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n317), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI22_X1  g0550(.A1(G283), .A2(new_n747), .B1(new_n750), .B2(G311), .ZN(new_n751));
  INV_X1    g0551(.A(G326), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n317), .A2(new_n310), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n211), .A2(new_n349), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n751), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n754), .A2(new_n745), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT99), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT99), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G303), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n301), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT101), .ZN(new_n763));
  INV_X1    g0563(.A(new_n462), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G190), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n744), .A2(new_n765), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n764), .A2(new_n767), .B1(new_n769), .B2(G329), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n753), .A2(new_n744), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT102), .B(KEYINPUT33), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(G317), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n763), .B(new_n770), .C1(new_n771), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n754), .A2(new_n748), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n756), .B(new_n774), .C1(G322), .C2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n760), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n778), .A2(G87), .B1(new_n323), .B2(new_n776), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n769), .A2(G159), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n301), .B1(new_n780), .B2(KEYINPUT32), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n747), .A2(G107), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n767), .A2(G97), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n437), .B2(new_n771), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT100), .Z(new_n786));
  NOR2_X1   g0586(.A1(new_n780), .A2(KEYINPUT32), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n755), .A2(new_n234), .B1(new_n749), .B2(new_n219), .ZN(new_n788));
  NOR4_X1   g0588(.A1(new_n783), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n741), .B1(new_n777), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n733), .A2(new_n728), .A3(new_n743), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n730), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT103), .ZN(G396));
  NAND2_X1  g0593(.A1(new_n670), .A2(new_n371), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n375), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n373), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n647), .A2(new_n663), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n689), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n796), .A2(new_n797), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n639), .A2(new_n663), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n723), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT105), .Z(new_n804));
  AOI21_X1  g0604(.A(new_n728), .B1(new_n723), .B2(new_n802), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n798), .A2(new_n731), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n301), .B1(new_n760), .B2(new_n207), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G87), .B2(new_n747), .ZN(new_n809));
  INV_X1    g0609(.A(new_n771), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G283), .ZN(new_n811));
  INV_X1    g0611(.A(new_n755), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G303), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n776), .A2(G294), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n814), .B(new_n784), .C1(new_n254), .C2(new_n749), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G311), .B2(new_n769), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n809), .A2(new_n811), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT104), .Z(new_n818));
  AOI22_X1  g0618(.A1(G143), .A2(new_n776), .B1(new_n750), .B2(G159), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n819), .B1(new_n820), .B2(new_n755), .C1(new_n322), .C2(new_n771), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT34), .Z(new_n822));
  INV_X1    g0622(.A(new_n767), .ZN(new_n823));
  INV_X1    g0623(.A(new_n323), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n769), .A2(G132), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n331), .B1(new_n437), .B2(new_n746), .C1(new_n760), .C2(new_n234), .ZN(new_n827));
  NOR4_X1   g0627(.A1(new_n822), .A2(new_n825), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n741), .B1(new_n818), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n741), .A2(new_n731), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n219), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n807), .A2(new_n728), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n806), .A2(new_n832), .ZN(G384));
  NAND2_X1  g0633(.A1(new_n571), .A2(new_n573), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n254), .B1(new_n834), .B2(KEYINPUT35), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n835), .B(new_n237), .C1(KEYINPUT35), .C2(new_n834), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT36), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n235), .A2(G77), .A3(new_n414), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(G50), .B2(new_n437), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n653), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n283), .A2(new_n670), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n311), .B(new_n841), .C1(new_n319), .C2(new_n284), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n313), .A2(new_n316), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n283), .B1(new_n843), .B2(new_n318), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n842), .B1(new_n844), .B2(new_n663), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n845), .A2(new_n719), .A3(new_n721), .A4(new_n800), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n662), .B1(new_n450), .B2(new_n452), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n448), .B1(new_n440), .B2(new_n442), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT106), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n443), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n425), .A2(KEYINPUT106), .A3(new_n432), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n848), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT37), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT107), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n450), .A2(new_n452), .B1(new_n449), .B2(new_n662), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT37), .B1(new_n425), .B2(new_n432), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n853), .A2(KEYINPUT107), .A3(KEYINPUT37), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n856), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n645), .A2(new_n433), .A3(new_n444), .ZN(new_n862));
  INV_X1    g0662(.A(new_n848), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n862), .A2(KEYINPUT108), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT108), .B1(new_n862), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT38), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n418), .A2(new_n263), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n439), .A2(new_n423), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n381), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n449), .A2(new_n662), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n443), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .B1(new_n857), .B2(new_n858), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n455), .A2(new_n456), .ZN(new_n875));
  INV_X1    g0675(.A(new_n445), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n868), .B(new_n874), .C1(new_n877), .C2(new_n662), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n847), .B(KEYINPUT40), .C1(new_n867), .C2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n641), .A2(new_n451), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n643), .A2(KEYINPUT77), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT18), .B1(new_n883), .B2(new_n449), .ZN(new_n884));
  INV_X1    g0684(.A(new_n456), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n876), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n871), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(new_n662), .A3(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n874), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n847), .B1(new_n878), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(KEYINPUT109), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT109), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n457), .A2(new_n661), .A3(new_n871), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n868), .B1(new_n895), .B2(new_n874), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n846), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(new_n898), .B2(KEYINPUT40), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n880), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n458), .A3(new_n722), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT109), .B1(new_n891), .B2(new_n892), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n898), .A2(new_n894), .A3(KEYINPUT40), .ZN(new_n903));
  OAI211_X1 g0703(.A(G330), .B(new_n879), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n458), .A2(G330), .A3(new_n722), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n901), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n646), .A2(new_n663), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n867), .A2(new_n878), .A3(KEYINPUT39), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT39), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n896), .B2(new_n897), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n910), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n645), .A2(new_n662), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n896), .A2(new_n897), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n646), .A2(new_n670), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n917), .A2(new_n842), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n801), .B2(new_n797), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n915), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n908), .B(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n458), .A2(new_n703), .A3(new_n693), .A4(new_n704), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n651), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n275), .A2(new_n654), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n837), .B1(new_n275), .B2(new_n840), .C1(new_n925), .C2(new_n926), .ZN(G367));
  INV_X1    g0727(.A(KEYINPUT114), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT44), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n610), .A2(new_n670), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n606), .A2(new_n614), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT110), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n931), .B(new_n932), .C1(new_n614), .C2(new_n663), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n628), .A2(KEYINPUT110), .A3(new_n613), .A4(new_n670), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n929), .B1(new_n679), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT93), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n668), .B(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT92), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n671), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n500), .A2(new_n533), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n677), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n678), .A2(new_n663), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n933), .A2(new_n934), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(KEYINPUT44), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n936), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT45), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n945), .B2(new_n946), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n679), .A2(new_n935), .A3(KEYINPUT45), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n948), .A2(new_n952), .A3(new_n675), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n675), .B1(new_n948), .B2(new_n952), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT113), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n666), .A2(new_n676), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(new_n674), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n724), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n705), .A2(new_n723), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT113), .B1(new_n961), .B2(new_n958), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n955), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n724), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n682), .B(KEYINPUT41), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n727), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n935), .A2(new_n667), .A3(new_n674), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT112), .Z(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT111), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n676), .B1(new_n669), .B2(new_n673), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n935), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT111), .B1(new_n946), .B2(new_n943), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT42), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT42), .B1(new_n972), .B2(new_n973), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n935), .A2(new_n678), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n670), .B1(new_n976), .B2(new_n614), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n663), .B1(new_n518), .B2(new_n519), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n624), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n635), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n978), .A2(KEYINPUT43), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n972), .A2(new_n973), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT42), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n976), .A2(new_n614), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n663), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT42), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n982), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT43), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n984), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n969), .B1(new_n983), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n984), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n978), .B2(new_n994), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n991), .A2(new_n993), .A3(new_n992), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n968), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n928), .B1(new_n966), .B2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n983), .A2(new_n996), .A3(new_n969), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n968), .B1(new_n999), .B2(new_n1000), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n965), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n963), .B2(new_n724), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1006), .B(KEYINPUT114), .C1(new_n727), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n331), .B1(new_n437), .B2(new_n823), .C1(new_n760), .C2(new_n824), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n768), .A2(new_n820), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n749), .A2(new_n234), .ZN(new_n1013));
  INV_X1    g0813(.A(G143), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n755), .A2(new_n1014), .B1(new_n746), .B2(new_n219), .ZN(new_n1015));
  NOR4_X1   g0815(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n322), .B2(new_n775), .C1(new_n410), .C2(new_n771), .ZN(new_n1017));
  XOR2_X1   g0817(.A(KEYINPUT115), .B(G311), .Z(new_n1018));
  OAI22_X1  g0818(.A1(new_n755), .A2(new_n1018), .B1(new_n775), .B2(new_n761), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n301), .B1(new_n746), .B2(new_n510), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n778), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT46), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n760), .B2(new_n254), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(new_n462), .C2(new_n771), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT116), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1019), .B(new_n1020), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G283), .A2(new_n750), .B1(new_n769), .B2(G317), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n1025), .C2(new_n1024), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n823), .A2(new_n207), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1017), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(KEYINPUT117), .B(KEYINPUT47), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n741), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n992), .A2(new_n740), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n737), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n742), .B1(new_n240), .B2(new_n367), .C1(new_n1036), .C2(new_n251), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n728), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1010), .A2(new_n1038), .ZN(G387));
  NAND2_X1  g0839(.A1(new_n960), .A2(new_n962), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n682), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT119), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(KEYINPUT119), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n724), .C2(new_n959), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n760), .A2(new_n219), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G159), .A2(new_n812), .B1(new_n776), .B2(G50), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n322), .B2(new_n768), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n823), .A2(new_n367), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1045), .A2(new_n1047), .A3(new_n301), .A4(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n325), .A2(new_n771), .B1(new_n437), .B2(new_n749), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT118), .Z(new_n1051));
  OAI211_X1 g0851(.A(new_n1049), .B(new_n1051), .C1(new_n206), .C2(new_n746), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G322), .A2(new_n812), .B1(new_n750), .B2(G303), .ZN(new_n1053));
  INV_X1    g0853(.A(G317), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n775), .C1(new_n771), .C2(new_n1018), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT48), .ZN(new_n1056));
  INV_X1    g0856(.A(G283), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1056), .B1(new_n1057), .B2(new_n823), .C1(new_n462), .C2(new_n760), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT49), .Z(new_n1059));
  OAI221_X1 g0859(.A(new_n301), .B1(new_n768), .B2(new_n752), .C1(new_n254), .C2(new_n746), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1052), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n741), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n364), .A2(new_n234), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT50), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n437), .A2(new_n219), .ZN(new_n1065));
  NOR4_X1   g0865(.A1(new_n1064), .A2(G45), .A3(new_n1065), .A4(new_n685), .ZN(new_n1066));
  INV_X1    g0866(.A(G45), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n737), .B1(new_n248), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n685), .A2(new_n240), .A3(new_n331), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n240), .A2(G107), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n742), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n669), .A2(new_n673), .A3(new_n740), .ZN(new_n1073));
  AND4_X1   g0873(.A1(new_n728), .A2(new_n1062), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n959), .B2(new_n727), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1044), .A2(new_n1075), .ZN(G393));
  NAND2_X1  g0876(.A1(new_n955), .A2(new_n727), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n946), .A2(new_n740), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n750), .A2(G294), .B1(new_n767), .B2(G116), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G317), .A2(new_n812), .B1(new_n776), .B2(G311), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT121), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n301), .B(new_n1079), .C1(new_n1081), .C2(KEYINPUT52), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(KEYINPUT52), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n769), .A2(G322), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n810), .A2(G303), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1083), .A2(new_n782), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1082), .B(new_n1086), .C1(G283), .C2(new_n778), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n810), .A2(G50), .B1(new_n750), .B2(new_n364), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n331), .B1(new_n768), .B2(new_n1014), .C1(new_n215), .C2(new_n746), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n778), .B2(new_n228), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT120), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n767), .A2(G77), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n755), .A2(new_n322), .B1(new_n775), .B2(new_n410), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  AND4_X1   g0894(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n741), .B1(new_n1087), .B2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n742), .B1(new_n240), .B2(new_n510), .C1(new_n257), .C2(new_n1036), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1078), .A2(new_n728), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n955), .B1(new_n960), .B2(new_n962), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n682), .B1(new_n1099), .B2(KEYINPUT122), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n955), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1040), .A2(new_n1101), .A3(KEYINPUT122), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n963), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1077), .B(new_n1098), .C1(new_n1100), .C2(new_n1103), .ZN(G390));
  AND3_X1   g0904(.A1(new_n853), .A2(KEYINPUT107), .A3(KEYINPUT37), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT107), .B1(new_n853), .B2(KEYINPUT37), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n859), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n862), .A2(new_n863), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT108), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n862), .A2(KEYINPUT108), .A3(new_n863), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n868), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n912), .A3(new_n897), .ZN(new_n1115));
  OAI21_X1  g0915(.A(KEYINPUT39), .B1(new_n878), .B2(new_n890), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n801), .A2(new_n797), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n845), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n909), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n702), .A2(new_n663), .A3(new_n796), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n797), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n910), .B1(new_n1122), .B2(new_n845), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n878), .B2(new_n867), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n798), .B1(new_n917), .B2(new_n842), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1126), .A2(G330), .A3(new_n719), .A4(new_n721), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT123), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1120), .A2(new_n1129), .A3(new_n1124), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n727), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1115), .A2(new_n1116), .A3(new_n731), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT54), .B(G143), .Z(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1137), .A2(new_n749), .B1(new_n820), .B2(new_n771), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G159), .B2(new_n767), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT124), .Z(new_n1140));
  AOI211_X1 g0940(.A(new_n301), .B(new_n1140), .C1(G125), .C2(new_n769), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n776), .A2(G132), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n747), .A2(G50), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n778), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT53), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n760), .B2(new_n322), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1144), .A2(new_n1146), .B1(G128), .B2(new_n812), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n755), .A2(new_n1057), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n778), .A2(G87), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n301), .B1(new_n771), .B2(new_n207), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G294), .B2(new_n769), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n775), .A2(new_n254), .B1(new_n749), .B2(new_n510), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G68), .B2(new_n747), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1150), .A2(new_n1092), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1148), .B1(new_n1149), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n741), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n325), .A2(new_n830), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1135), .A2(new_n728), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1134), .A2(new_n1159), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1121), .A2(new_n797), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n719), .A2(G330), .A3(new_n721), .A4(new_n800), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n918), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1161), .A2(new_n1163), .A3(new_n1127), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1163), .A2(new_n1127), .B1(new_n797), .B2(new_n801), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n923), .A2(new_n651), .A3(new_n906), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1133), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1131), .A2(new_n1168), .A3(new_n1132), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1170), .A2(new_n682), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1160), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(G378));
  INV_X1    g0973(.A(new_n1167), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n330), .A2(new_n662), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n356), .B(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n914), .B2(new_n920), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n909), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n919), .B1(new_n878), .B2(new_n890), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n915), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1182), .A2(new_n1185), .A3(new_n1179), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n904), .A2(new_n1181), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n914), .A2(new_n920), .A3(new_n1180), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1179), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1188), .A2(new_n1189), .B1(new_n900), .B2(G330), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1175), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT57), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n904), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1188), .A2(new_n1189), .A3(G330), .A4(new_n900), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(KEYINPUT57), .A3(new_n1175), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1193), .A2(new_n682), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n727), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1179), .A2(new_n731), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n292), .A2(new_n331), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n207), .B2(new_n775), .C1(new_n367), .C2(new_n749), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n823), .A2(new_n437), .B1(new_n824), .B2(new_n746), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1203), .B(new_n1045), .C1(G97), .C2(new_n810), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1057), .B2(new_n768), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1202), .B(new_n1205), .C1(G116), .C2(new_n812), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n778), .A2(new_n1136), .B1(G125), .B2(new_n812), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G128), .A2(new_n776), .B1(new_n750), .B2(G137), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n322), .C2(new_n823), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G132), .B2(new_n810), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT59), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G33), .B(G41), .C1(new_n769), .C2(G124), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n410), .C2(new_n746), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n234), .B1(G33), .B2(G41), .C1(new_n292), .C2(new_n331), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1207), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n741), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n830), .A2(new_n234), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1200), .A2(new_n728), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1199), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1198), .A2(new_n1222), .ZN(G375));
  NAND2_X1  g1023(.A1(new_n830), .A2(new_n437), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n728), .B(new_n1224), .C1(new_n845), .C2(new_n732), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n749), .A2(new_n207), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n331), .B1(new_n778), .B2(G97), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n254), .B2(new_n771), .C1(new_n1057), .C2(new_n775), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(G294), .C2(new_n812), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1048), .B1(G77), .B2(new_n747), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(new_n761), .C2(new_n768), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT125), .Z(new_n1232));
  NOR2_X1   g1032(.A1(new_n760), .A2(new_n410), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n769), .A2(G128), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n331), .C1(new_n234), .C2(new_n823), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n824), .A2(new_n746), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n749), .A2(new_n322), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n775), .A2(new_n820), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n812), .A2(G132), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(new_n771), .C2(new_n1137), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1232), .B1(new_n1233), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1225), .B1(new_n1242), .B2(new_n741), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1166), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(new_n727), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n965), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1245), .B1(new_n1247), .B2(new_n1168), .ZN(G381));
  INV_X1    g1048(.A(G390), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1010), .A2(new_n1038), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(G396), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1044), .A2(new_n1251), .A3(new_n1075), .ZN(new_n1252));
  OR4_X1    g1052(.A1(G384), .A2(new_n1250), .A3(G381), .A4(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1198), .A2(new_n1172), .A3(new_n1222), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1253), .A2(new_n1254), .ZN(G407));
  AND2_X1   g1055(.A1(new_n1253), .A2(G343), .ZN(new_n1256));
  OAI21_X1  g1056(.A(G213), .B1(new_n1256), .B2(new_n1254), .ZN(G409));
  AND3_X1   g1057(.A1(new_n1196), .A2(KEYINPUT57), .A3(new_n1175), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1175), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n683), .ZN(new_n1260));
  OAI21_X1  g1060(.A(G378), .B1(new_n1260), .B2(new_n1221), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n683), .B1(new_n1246), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1168), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(new_n1262), .C2(new_n1246), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1265), .A2(G384), .A3(new_n1245), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G384), .B1(new_n1265), .B2(new_n1245), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n658), .A2(G343), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1196), .A2(new_n965), .A3(new_n1175), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT126), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1196), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1194), .A2(KEYINPUT126), .A3(new_n1195), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n727), .A3(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1172), .A2(new_n1271), .A3(new_n1220), .A4(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1261), .A2(new_n1268), .A3(new_n1270), .A4(new_n1276), .ZN(new_n1277));
  XOR2_X1   g1077(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1261), .A2(new_n1270), .A3(new_n1276), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1269), .A2(G2897), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1268), .B(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1269), .B1(G375), .B2(G378), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n1286), .A3(new_n1268), .A4(new_n1276), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT61), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1279), .A2(new_n1284), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G387), .A2(G390), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G393), .A2(G396), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1290), .A2(new_n1250), .A3(new_n1252), .A4(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1252), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1010), .A2(new_n1038), .A3(new_n1249), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1249), .B1(new_n1010), .B2(new_n1038), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1293), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1292), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1289), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT61), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1268), .A4(new_n1276), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1277), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1300), .B(new_n1301), .C1(new_n1302), .C2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1299), .A2(new_n1305), .ZN(G405));
  NAND2_X1  g1106(.A1(new_n1261), .A2(new_n1254), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1268), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1261), .B(new_n1254), .C1(new_n1267), .C2(new_n1266), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1310), .B(new_n1297), .ZN(G402));
endmodule


