

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578;

  NOR2_X2 U323 ( .A1(n504), .A2(n503), .ZN(n505) );
  NOR2_X1 U324 ( .A1(n540), .A2(n539), .ZN(n561) );
  XOR2_X1 U325 ( .A(G64GAT), .B(G92GAT), .Z(n291) );
  INV_X1 U326 ( .A(n439), .ZN(n302) );
  XNOR2_X1 U327 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U328 ( .A(n305), .B(n304), .ZN(n306) );
  NOR2_X2 U329 ( .A1(n545), .A2(n544), .ZN(n556) );
  XOR2_X1 U330 ( .A(n343), .B(n342), .Z(n534) );
  XOR2_X1 U331 ( .A(n541), .B(KEYINPUT28), .Z(n493) );
  XOR2_X1 U332 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n449) );
  XOR2_X1 U333 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n293) );
  XNOR2_X1 U334 ( .A(KEYINPUT72), .B(KEYINPUT31), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n293), .B(n292), .ZN(n307) );
  XOR2_X1 U336 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n295) );
  NAND2_X1 U337 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U339 ( .A(n296), .B(KEYINPUT71), .Z(n300) );
  XNOR2_X1 U340 ( .A(G106GAT), .B(G78GAT), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n297), .B(G148GAT), .ZN(n345) );
  XNOR2_X1 U342 ( .A(G176GAT), .B(G204GAT), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n291), .B(n298), .ZN(n369) );
  XNOR2_X1 U344 ( .A(n345), .B(n369), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n305) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G71GAT), .Z(n335) );
  XOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .Z(n405) );
  XNOR2_X1 U348 ( .A(n335), .B(n405), .ZN(n303) );
  XNOR2_X1 U349 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n301), .B(KEYINPUT13), .ZN(n439) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n568) );
  XOR2_X1 U352 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n309) );
  XNOR2_X1 U353 ( .A(G197GAT), .B(G113GAT), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n318) );
  XOR2_X1 U355 ( .A(G141GAT), .B(G22GAT), .Z(n349) );
  XNOR2_X1 U356 ( .A(G15GAT), .B(G1GAT), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n310), .B(KEYINPUT68), .ZN(n440) );
  XOR2_X1 U358 ( .A(n349), .B(n440), .Z(n312) );
  NAND2_X1 U359 ( .A1(G229GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U361 ( .A(n313), .B(KEYINPUT29), .Z(n316) );
  XNOR2_X1 U362 ( .A(G169GAT), .B(G36GAT), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n314), .B(G8GAT), .ZN(n370) );
  XNOR2_X1 U364 ( .A(n370), .B(KEYINPUT67), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U367 ( .A(KEYINPUT7), .B(G50GAT), .Z(n320) );
  XNOR2_X1 U368 ( .A(G43GAT), .B(G29GAT), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U370 ( .A(KEYINPUT8), .B(n321), .Z(n410) );
  XOR2_X1 U371 ( .A(n322), .B(n410), .Z(n562) );
  XNOR2_X1 U372 ( .A(KEYINPUT69), .B(n562), .ZN(n546) );
  NAND2_X1 U373 ( .A1(n568), .A2(n546), .ZN(n323) );
  XOR2_X1 U374 ( .A(KEYINPUT75), .B(n323), .Z(n461) );
  XOR2_X1 U375 ( .A(G183GAT), .B(KEYINPUT19), .Z(n325) );
  XNOR2_X1 U376 ( .A(KEYINPUT85), .B(KEYINPUT17), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U378 ( .A(n326), .B(KEYINPUT18), .Z(n328) );
  XNOR2_X1 U379 ( .A(KEYINPUT86), .B(G190GAT), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n365) );
  XOR2_X1 U381 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n330) );
  XNOR2_X1 U382 ( .A(G15GAT), .B(G176GAT), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n365), .B(n331), .ZN(n343) );
  XOR2_X1 U385 ( .A(KEYINPUT20), .B(G99GAT), .Z(n333) );
  XNOR2_X1 U386 ( .A(G43GAT), .B(G134GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U388 ( .A(n335), .B(n334), .Z(n337) );
  NAND2_X1 U389 ( .A1(G227GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U391 ( .A(n338), .B(KEYINPUT87), .Z(n341) );
  XNOR2_X1 U392 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n339), .B(G127GAT), .ZN(n385) );
  XNOR2_X1 U394 ( .A(G169GAT), .B(n385), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U396 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n344), .B(KEYINPUT2), .ZN(n384) );
  XOR2_X1 U398 ( .A(KEYINPUT76), .B(G162GAT), .Z(n406) );
  XOR2_X1 U399 ( .A(n384), .B(n406), .Z(n351) );
  XOR2_X1 U400 ( .A(n345), .B(G204GAT), .Z(n347) );
  NAND2_X1 U401 ( .A1(G228GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U405 ( .A(KEYINPUT92), .B(KEYINPUT24), .Z(n353) );
  XNOR2_X1 U406 ( .A(G50GAT), .B(KEYINPUT89), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U408 ( .A(n355), .B(n354), .Z(n363) );
  XOR2_X1 U409 ( .A(KEYINPUT90), .B(G218GAT), .Z(n357) );
  XNOR2_X1 U410 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U412 ( .A(G197GAT), .B(n358), .Z(n364) );
  XOR2_X1 U413 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n360) );
  XNOR2_X1 U414 ( .A(KEYINPUT91), .B(KEYINPUT88), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n364), .B(n361), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n541) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n374) );
  XOR2_X1 U419 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n367) );
  NAND2_X1 U420 ( .A1(G226GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U422 ( .A(n368), .B(KEYINPUT96), .Z(n372) );
  XNOR2_X1 U423 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U425 ( .A(n374), .B(n373), .Z(n535) );
  XNOR2_X1 U426 ( .A(n535), .B(KEYINPUT27), .ZN(n398) );
  XOR2_X1 U427 ( .A(G85GAT), .B(G162GAT), .Z(n376) );
  XNOR2_X1 U428 ( .A(G141GAT), .B(G120GAT), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U430 ( .A(G134GAT), .B(KEYINPUT78), .Z(n414) );
  XOR2_X1 U431 ( .A(n377), .B(n414), .Z(n379) );
  XNOR2_X1 U432 ( .A(G29GAT), .B(G148GAT), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U434 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n381) );
  XNOR2_X1 U435 ( .A(G1GAT), .B(G57GAT), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U437 ( .A(n383), .B(n382), .Z(n387) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U439 ( .A(n387), .B(n386), .ZN(n392) );
  XOR2_X1 U440 ( .A(KEYINPUT1), .B(KEYINPUT93), .Z(n389) );
  NAND2_X1 U441 ( .A1(G225GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U443 ( .A(KEYINPUT6), .B(n390), .Z(n391) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n540) );
  NAND2_X1 U445 ( .A1(n398), .A2(n540), .ZN(n506) );
  NOR2_X1 U446 ( .A1(n493), .A2(n506), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n393), .B(KEYINPUT97), .ZN(n394) );
  NOR2_X1 U448 ( .A1(n534), .A2(n394), .ZN(n404) );
  NAND2_X1 U449 ( .A1(n534), .A2(n535), .ZN(n395) );
  NAND2_X1 U450 ( .A1(n541), .A2(n395), .ZN(n396) );
  XNOR2_X1 U451 ( .A(KEYINPUT25), .B(n396), .ZN(n401) );
  NOR2_X1 U452 ( .A1(n534), .A2(n541), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n397), .B(KEYINPUT26), .ZN(n560) );
  NAND2_X1 U454 ( .A1(n398), .A2(n560), .ZN(n399) );
  XOR2_X1 U455 ( .A(KEYINPUT98), .B(n399), .Z(n400) );
  NOR2_X1 U456 ( .A1(n401), .A2(n400), .ZN(n402) );
  NOR2_X1 U457 ( .A1(n402), .A2(n540), .ZN(n403) );
  NOR2_X1 U458 ( .A1(n404), .A2(n403), .ZN(n458) );
  XOR2_X1 U459 ( .A(KEYINPUT65), .B(KEYINPUT10), .Z(n408) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U461 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U462 ( .A(n409), .B(KEYINPUT9), .Z(n413) );
  INV_X1 U463 ( .A(n410), .ZN(n411) );
  XOR2_X1 U464 ( .A(n411), .B(G218GAT), .Z(n412) );
  XNOR2_X1 U465 ( .A(n413), .B(n412), .ZN(n418) );
  XOR2_X1 U466 ( .A(G92GAT), .B(n414), .Z(n416) );
  NAND2_X1 U467 ( .A1(G232GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U468 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U469 ( .A(n418), .B(n417), .Z(n423) );
  XOR2_X1 U470 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n420) );
  XNOR2_X1 U471 ( .A(G190GAT), .B(G106GAT), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U473 ( .A(G36GAT), .B(n421), .ZN(n422) );
  XOR2_X1 U474 ( .A(n423), .B(n422), .Z(n531) );
  INV_X1 U475 ( .A(n531), .ZN(n555) );
  XOR2_X1 U476 ( .A(G155GAT), .B(G78GAT), .Z(n425) );
  XNOR2_X1 U477 ( .A(G22GAT), .B(G211GAT), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U479 ( .A(G64GAT), .B(G71GAT), .Z(n427) );
  XNOR2_X1 U480 ( .A(G183GAT), .B(G127GAT), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U482 ( .A(n429), .B(n428), .Z(n434) );
  XOR2_X1 U483 ( .A(KEYINPUT79), .B(KEYINPUT81), .Z(n431) );
  NAND2_X1 U484 ( .A1(G231GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U486 ( .A(KEYINPUT80), .B(n432), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U488 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n436) );
  XNOR2_X1 U489 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U491 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U493 ( .A(n442), .B(n441), .Z(n552) );
  INV_X1 U494 ( .A(n552), .ZN(n571) );
  NOR2_X1 U495 ( .A1(n555), .A2(n571), .ZN(n443) );
  XOR2_X1 U496 ( .A(KEYINPUT82), .B(n443), .Z(n444) );
  XNOR2_X1 U497 ( .A(n444), .B(KEYINPUT16), .ZN(n445) );
  NOR2_X1 U498 ( .A1(n458), .A2(n445), .ZN(n446) );
  XNOR2_X1 U499 ( .A(KEYINPUT99), .B(n446), .ZN(n472) );
  NOR2_X1 U500 ( .A1(n461), .A2(n472), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n447), .B(KEYINPUT100), .ZN(n455) );
  NAND2_X1 U502 ( .A1(n455), .A2(n540), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U504 ( .A(G1GAT), .B(n450), .ZN(G1324GAT) );
  NAND2_X1 U505 ( .A1(n455), .A2(n535), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n451), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U507 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n453) );
  NAND2_X1 U508 ( .A1(n455), .A2(n534), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U510 ( .A(G15GAT), .B(n454), .ZN(G1326GAT) );
  XOR2_X1 U511 ( .A(G22GAT), .B(KEYINPUT103), .Z(n457) );
  NAND2_X1 U512 ( .A1(n493), .A2(n455), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n457), .B(n456), .ZN(G1327GAT) );
  XOR2_X1 U514 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n464) );
  XNOR2_X1 U515 ( .A(KEYINPUT36), .B(n531), .ZN(n575) );
  NOR2_X1 U516 ( .A1(n575), .A2(n458), .ZN(n459) );
  NAND2_X1 U517 ( .A1(n459), .A2(n571), .ZN(n460) );
  XOR2_X1 U518 ( .A(KEYINPUT37), .B(n460), .Z(n483) );
  NOR2_X1 U519 ( .A1(n483), .A2(n461), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(KEYINPUT38), .ZN(n469) );
  NAND2_X1 U521 ( .A1(n469), .A2(n540), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U523 ( .A(G29GAT), .B(n465), .ZN(G1328GAT) );
  NAND2_X1 U524 ( .A1(n469), .A2(n535), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n466), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U526 ( .A1(n469), .A2(n534), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT40), .ZN(n468) );
  XNOR2_X1 U528 ( .A(G43GAT), .B(n468), .ZN(G1330GAT) );
  NAND2_X1 U529 ( .A1(n469), .A2(n493), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n470), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U531 ( .A(n568), .B(KEYINPUT41), .Z(n525) );
  INV_X1 U532 ( .A(n525), .ZN(n548) );
  NAND2_X1 U533 ( .A1(n562), .A2(n548), .ZN(n471) );
  XOR2_X1 U534 ( .A(KEYINPUT105), .B(n471), .Z(n482) );
  NOR2_X1 U535 ( .A1(n472), .A2(n482), .ZN(n478) );
  NAND2_X1 U536 ( .A1(n478), .A2(n540), .ZN(n473) );
  XNOR2_X1 U537 ( .A(KEYINPUT42), .B(n473), .ZN(n474) );
  XNOR2_X1 U538 ( .A(G57GAT), .B(n474), .ZN(G1332GAT) );
  NAND2_X1 U539 ( .A1(n535), .A2(n478), .ZN(n475) );
  XNOR2_X1 U540 ( .A(n475), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U541 ( .A1(n534), .A2(n478), .ZN(n476) );
  XNOR2_X1 U542 ( .A(n476), .B(KEYINPUT106), .ZN(n477) );
  XNOR2_X1 U543 ( .A(G71GAT), .B(n477), .ZN(G1334GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n480) );
  NAND2_X1 U545 ( .A1(n478), .A2(n493), .ZN(n479) );
  XNOR2_X1 U546 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U547 ( .A(G78GAT), .B(n481), .Z(G1335GAT) );
  XNOR2_X1 U548 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n485) );
  NOR2_X1 U549 ( .A1(n483), .A2(n482), .ZN(n489) );
  NAND2_X1 U550 ( .A1(n489), .A2(n540), .ZN(n484) );
  XNOR2_X1 U551 ( .A(n485), .B(n484), .ZN(G1336GAT) );
  NAND2_X1 U552 ( .A1(n535), .A2(n489), .ZN(n486) );
  XNOR2_X1 U553 ( .A(n486), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U554 ( .A(G99GAT), .B(KEYINPUT109), .Z(n488) );
  NAND2_X1 U555 ( .A1(n489), .A2(n534), .ZN(n487) );
  XNOR2_X1 U556 ( .A(n488), .B(n487), .ZN(G1338GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n491) );
  NAND2_X1 U558 ( .A1(n489), .A2(n493), .ZN(n490) );
  XNOR2_X1 U559 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U560 ( .A(G106GAT), .B(n492), .Z(G1339GAT) );
  INV_X1 U561 ( .A(n493), .ZN(n509) );
  NOR2_X1 U562 ( .A1(n562), .A2(n525), .ZN(n494) );
  XNOR2_X1 U563 ( .A(n494), .B(KEYINPUT46), .ZN(n495) );
  NOR2_X1 U564 ( .A1(n555), .A2(n495), .ZN(n496) );
  NAND2_X1 U565 ( .A1(n571), .A2(n496), .ZN(n497) );
  XNOR2_X1 U566 ( .A(n497), .B(KEYINPUT47), .ZN(n504) );
  XNOR2_X1 U567 ( .A(KEYINPUT111), .B(KEYINPUT45), .ZN(n498) );
  XNOR2_X1 U568 ( .A(n498), .B(KEYINPUT64), .ZN(n500) );
  NOR2_X1 U569 ( .A1(n575), .A2(n571), .ZN(n499) );
  XOR2_X1 U570 ( .A(n500), .B(n499), .Z(n501) );
  NAND2_X1 U571 ( .A1(n568), .A2(n501), .ZN(n502) );
  NOR2_X1 U572 ( .A1(n502), .A2(n546), .ZN(n503) );
  XNOR2_X1 U573 ( .A(KEYINPUT48), .B(n505), .ZN(n537) );
  NOR2_X1 U574 ( .A1(n537), .A2(n506), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n522), .A2(n534), .ZN(n507) );
  XOR2_X1 U576 ( .A(KEYINPUT112), .B(n507), .Z(n508) );
  NAND2_X1 U577 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n510), .B(KEYINPUT113), .ZN(n517) );
  NAND2_X1 U579 ( .A1(n546), .A2(n517), .ZN(n511) );
  XNOR2_X1 U580 ( .A(G113GAT), .B(n511), .ZN(G1340GAT) );
  XOR2_X1 U581 ( .A(G120GAT), .B(KEYINPUT49), .Z(n513) );
  NAND2_X1 U582 ( .A1(n517), .A2(n548), .ZN(n512) );
  XNOR2_X1 U583 ( .A(n513), .B(n512), .ZN(G1341GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n515) );
  NAND2_X1 U585 ( .A1(n517), .A2(n552), .ZN(n514) );
  XNOR2_X1 U586 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U587 ( .A(G127GAT), .B(n516), .Z(G1342GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n519) );
  NAND2_X1 U589 ( .A1(n517), .A2(n555), .ZN(n518) );
  XNOR2_X1 U590 ( .A(n519), .B(n518), .ZN(n521) );
  XOR2_X1 U591 ( .A(G134GAT), .B(KEYINPUT115), .Z(n520) );
  XNOR2_X1 U592 ( .A(n521), .B(n520), .ZN(G1343GAT) );
  NAND2_X1 U593 ( .A1(n522), .A2(n560), .ZN(n530) );
  NOR2_X1 U594 ( .A1(n562), .A2(n530), .ZN(n524) );
  XNOR2_X1 U595 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n523) );
  XNOR2_X1 U596 ( .A(n524), .B(n523), .ZN(G1344GAT) );
  NOR2_X1 U597 ( .A1(n525), .A2(n530), .ZN(n527) );
  XNOR2_X1 U598 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n526) );
  XNOR2_X1 U599 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U600 ( .A(G148GAT), .B(n528), .ZN(G1345GAT) );
  NOR2_X1 U601 ( .A1(n571), .A2(n530), .ZN(n529) );
  XOR2_X1 U602 ( .A(G155GAT), .B(n529), .Z(G1346GAT) );
  NOR2_X1 U603 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U604 ( .A(G162GAT), .B(n532), .Z(n533) );
  XNOR2_X1 U605 ( .A(KEYINPUT118), .B(n533), .ZN(G1347GAT) );
  INV_X1 U606 ( .A(n534), .ZN(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n543) );
  XNOR2_X1 U608 ( .A(KEYINPUT119), .B(n535), .ZN(n536) );
  NOR2_X1 U609 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U610 ( .A(KEYINPUT54), .B(n538), .Z(n539) );
  NAND2_X1 U611 ( .A1(n561), .A2(n541), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U613 ( .A1(n556), .A2(n546), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n550) );
  NAND2_X1 U616 ( .A1(n556), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(n551), .ZN(G1349GAT) );
  XOR2_X1 U619 ( .A(G183GAT), .B(KEYINPUT121), .Z(n554) );
  NAND2_X1 U620 ( .A1(n556), .A2(n552), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1350GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n558) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U625 ( .A(G190GAT), .B(n559), .Z(G1351GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n574) );
  NOR2_X1 U627 ( .A1(n562), .A2(n574), .ZN(n567) );
  XOR2_X1 U628 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n564) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  NOR2_X1 U633 ( .A1(n568), .A2(n574), .ZN(n570) );
  XNOR2_X1 U634 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1353GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n574), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1354GAT) );
  NOR2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U640 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U642 ( .A(G218GAT), .B(n578), .Z(G1355GAT) );
endmodule

