//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT24), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g004(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n221));
  OAI211_X1 g020(.A(KEYINPUT23), .B(new_n213), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n205), .A2(new_n209), .A3(new_n223), .A4(new_n206), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n211), .A2(new_n219), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT25), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(KEYINPUT67), .A3(new_n226), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT68), .B(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n207), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n205), .A2(new_n206), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT23), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n234), .A2(KEYINPUT25), .A3(new_n219), .A4(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n229), .A2(new_n230), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT27), .B(G183gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n231), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT28), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n214), .A2(new_n242), .A3(new_n215), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n243), .B(new_n203), .C1(new_n242), .C2(new_n214), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G226gat), .A2(G233gat), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n237), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(new_n237), .B2(new_n245), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT22), .ZN(new_n252));
  INV_X1    g051(.A(G211gat), .ZN(new_n253));
  INV_X1    g052(.A(G218gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT74), .ZN(new_n256));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT74), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n258), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G211gat), .B(G218gat), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n260), .B(new_n262), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n247), .A2(new_n251), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n260), .B(new_n261), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n225), .A2(KEYINPUT67), .A3(new_n226), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT67), .B1(new_n225), .B2(new_n226), .ZN(new_n267));
  INV_X1    g066(.A(new_n236), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n241), .A2(new_n244), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n249), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n237), .A2(new_n245), .A3(new_n246), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n265), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT37), .B1(new_n264), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT75), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G8gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n277), .B(G36gat), .Z(new_n278));
  OAI21_X1  g077(.A(new_n263), .B1(new_n247), .B2(new_n251), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT37), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n271), .A2(new_n265), .A3(new_n272), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n274), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT91), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT38), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(new_n283), .B2(KEYINPUT38), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G57gat), .B(G85gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n293));
  NAND2_X1  g092(.A1(G225gat), .A2(G233gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G113gat), .B(G120gat), .ZN(new_n296));
  OAI21_X1  g095(.A(G127gat), .B1(new_n296), .B2(KEYINPUT1), .ZN(new_n297));
  INV_X1    g096(.A(G120gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G113gat), .ZN(new_n299));
  INV_X1    g098(.A(G113gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G120gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303));
  INV_X1    g102(.A(G127gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n297), .A2(new_n305), .A3(G134gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  INV_X1    g106(.A(G155gat), .ZN(new_n308));
  INV_X1    g107(.A(G162gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n307), .B1(new_n310), .B2(KEYINPUT2), .ZN(new_n311));
  INV_X1    g110(.A(G148gat), .ZN(new_n312));
  INV_X1    g111(.A(G141gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT77), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G141gat), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n312), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n313), .A2(G148gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n311), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n310), .A2(new_n307), .ZN(new_n320));
  XNOR2_X1  g119(.A(G141gat), .B(G148gat), .ZN(new_n321));
  OR2_X1    g120(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n322));
  NAND2_X1  g121(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n320), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(G134gat), .B1(new_n297), .B2(new_n305), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n306), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G134gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n304), .B1(new_n302), .B2(new_n303), .ZN(new_n330));
  AOI211_X1 g129(.A(KEYINPUT1), .B(G127gat), .C1(new_n299), .C2(new_n301), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n297), .A2(new_n305), .A3(G134gat), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n332), .A2(new_n333), .B1(new_n319), .B2(new_n325), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n295), .B1(new_n328), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n326), .B1(new_n306), .B2(new_n327), .ZN(new_n338));
  INV_X1    g137(.A(new_n318), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT77), .B(G141gat), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n339), .B1(new_n340), .B2(new_n312), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n312), .A2(G141gat), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n322), .B(new_n323), .C1(new_n318), .C2(new_n342), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n341), .A2(new_n311), .B1(new_n343), .B2(new_n320), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n332), .A2(new_n344), .A3(new_n333), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n294), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT5), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n337), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n336), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n319), .A2(new_n325), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n350), .B1(new_n319), .B2(new_n325), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n332), .A2(new_n333), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n295), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n345), .A2(KEYINPUT4), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT4), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n332), .A2(new_n344), .A3(new_n357), .A4(new_n333), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n355), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n355), .B2(new_n359), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n349), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n306), .A2(new_n327), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n357), .A4(new_n344), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n358), .A2(KEYINPUT81), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n366), .A2(new_n367), .A3(new_n356), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n354), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n347), .A3(new_n294), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT82), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(new_n367), .A3(new_n356), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n347), .A4(new_n355), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n292), .B(new_n293), .C1(new_n363), .C2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT85), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n355), .A2(new_n359), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n355), .A2(new_n359), .A3(new_n360), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n380), .A2(new_n336), .A3(new_n348), .A4(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(new_n371), .A3(new_n374), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n383), .A2(KEYINPUT85), .A3(new_n292), .A4(new_n293), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n292), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n382), .A2(new_n386), .A3(new_n371), .A4(new_n374), .ZN(new_n387));
  INV_X1    g186(.A(new_n293), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n371), .A2(new_n374), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n386), .B1(new_n390), .B2(new_n382), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT90), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n383), .A2(new_n292), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n393), .A2(new_n394), .A3(new_n388), .A4(new_n387), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n283), .A2(KEYINPUT38), .ZN(new_n397));
  INV_X1    g196(.A(new_n278), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n279), .A2(new_n398), .A3(new_n281), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n287), .A2(new_n385), .A3(new_n396), .A4(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT92), .ZN(new_n403));
  XNOR2_X1  g202(.A(G78gat), .B(G106gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT31), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G50gat), .ZN(new_n406));
  INV_X1    g205(.A(G22gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(G228gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n260), .A2(new_n409), .A3(new_n261), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n248), .B(new_n410), .C1(new_n265), .C2(new_n409), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n344), .B1(new_n411), .B2(new_n350), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n263), .B1(KEYINPUT29), .B2(new_n351), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n408), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n408), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT3), .B1(new_n265), .B2(new_n248), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n416), .B(new_n413), .C1(new_n417), .C2(new_n344), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n407), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT87), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n406), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n260), .A2(new_n261), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n260), .A2(new_n261), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n422), .A2(new_n423), .A3(new_n409), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n410), .A2(new_n248), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n350), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n414), .B1(new_n426), .B2(new_n326), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n418), .B1(new_n427), .B2(new_n416), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(G22gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n415), .A2(new_n407), .A3(new_n418), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(KEYINPUT87), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n421), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(new_n430), .A3(new_n406), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT88), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT88), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n429), .A2(new_n435), .A3(new_n430), .A4(new_n406), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n432), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n372), .A2(new_n369), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n295), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n338), .A2(new_n345), .A3(new_n294), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(KEYINPUT39), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT39), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(new_n442), .A3(new_n295), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT89), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n443), .A2(new_n444), .A3(new_n386), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n443), .B2(new_n386), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT40), .B(new_n441), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  OR4_X1    g246(.A1(KEYINPUT30), .A2(new_n264), .A3(new_n273), .A4(new_n278), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n278), .B1(new_n264), .B2(new_n273), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(KEYINPUT30), .A3(new_n399), .ZN(new_n450));
  AND4_X1   g249(.A1(new_n393), .A2(new_n447), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n437), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n402), .A2(new_n403), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n354), .B1(new_n269), .B2(new_n270), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT34), .ZN(new_n458));
  INV_X1    g257(.A(G227gat), .ZN(new_n459));
  INV_X1    g258(.A(G233gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n237), .A2(new_n364), .A3(new_n245), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n457), .A2(new_n458), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT71), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n237), .A2(new_n364), .A3(new_n245), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n364), .B1(new_n237), .B2(new_n245), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT70), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT70), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n457), .A2(new_n469), .A3(new_n463), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n462), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT34), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT32), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G43gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(G71gat), .B(G99gat), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n478), .B(new_n479), .Z(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n480), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n474), .B(KEYINPUT32), .C1(new_n476), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n473), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n465), .A2(new_n481), .A3(new_n472), .A4(new_n483), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(KEYINPUT73), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT73), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n485), .A2(KEYINPUT36), .A3(new_n486), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n378), .A2(new_n384), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n387), .A2(KEYINPUT84), .A3(new_n388), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n495), .A2(new_n393), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n389), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n494), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n448), .A2(new_n450), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n437), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n403), .B1(new_n402), .B2(new_n455), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n456), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n501), .B1(new_n396), .B2(new_n385), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n489), .ZN(new_n507));
  INV_X1    g306(.A(new_n437), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT35), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n485), .A2(new_n486), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(new_n437), .ZN(new_n513));
  INV_X1    g312(.A(new_n499), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT35), .A4(new_n500), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n202), .B1(new_n505), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n402), .A2(new_n455), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT92), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n402), .A2(new_n455), .A3(new_n403), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n519), .A2(new_n502), .A3(new_n493), .A4(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n511), .A2(new_n515), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT93), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(G1gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT16), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G1gat), .B2(new_n525), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G43gat), .B(G50gat), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT95), .B1(new_n532), .B2(KEYINPUT15), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(KEYINPUT15), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n533), .B(new_n534), .Z(new_n535));
  NAND2_X1  g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT94), .ZN(new_n537));
  NOR2_X1   g336(.A1(G29gat), .A2(G36gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT14), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT96), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n537), .ZN(new_n542));
  OAI211_X1 g341(.A(KEYINPUT15), .B(new_n532), .C1(new_n542), .C2(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(KEYINPUT17), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n546), .B1(new_n541), .B2(new_n543), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n531), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n544), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n549), .A2(new_n531), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT18), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n544), .B(new_n531), .Z(new_n556));
  XOR2_X1   g355(.A(new_n551), .B(KEYINPUT13), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n554), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n548), .A2(new_n550), .A3(new_n551), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n555), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT11), .B(G169gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G197gat), .ZN(new_n563));
  XOR2_X1   g362(.A(G113gat), .B(G141gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT12), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n555), .A2(new_n566), .A3(new_n558), .A4(new_n560), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G57gat), .B(G64gat), .Z(new_n571));
  INV_X1    g370(.A(KEYINPUT9), .ZN(new_n572));
  INV_X1    g371(.A(G71gat), .ZN(new_n573));
  INV_X1    g372(.A(G78gat), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G71gat), .B(G78gat), .Z(new_n577));
  OR2_X1    g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  INV_X1    g381(.A(G85gat), .ZN(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(KEYINPUT8), .A2(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(new_n583), .B2(new_n584), .ZN(new_n587));
  NAND4_X1  g386(.A1(KEYINPUT100), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G99gat), .B(G106gat), .Z(new_n590));
  OR2_X1    g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n581), .A2(KEYINPUT10), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n580), .B(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n595), .B2(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n595), .A2(G230gat), .A3(G233gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(new_n213), .ZN(new_n602));
  INV_X1    g401(.A(G204gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n600), .B(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n570), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n524), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT21), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n531), .B1(new_n609), .B2(new_n580), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n610), .A2(G211gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(G211gat), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n611), .B2(new_n613), .ZN(new_n615));
  XOR2_X1   g414(.A(G127gat), .B(G155gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT20), .ZN(new_n617));
  OR3_X1    g416(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT19), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT98), .B(G183gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n617), .B1(new_n614), .B2(new_n615), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n618), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n618), .B2(new_n623), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n594), .B1(new_n545), .B2(new_n547), .ZN(new_n630));
  NAND3_X1  g429(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n544), .A2(new_n591), .A3(new_n592), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G190gat), .B(G218gat), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n635), .A2(new_n636), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT99), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n639), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n633), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n643), .B1(new_n633), .B2(new_n638), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n629), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n628), .A3(new_n644), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n627), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n608), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n514), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n526), .ZN(G1324gat));
  NAND3_X1  g453(.A1(new_n608), .A2(new_n651), .A3(new_n501), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT16), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(new_n656), .B2(new_n530), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT42), .ZN(new_n658));
  NAND2_X1  g457(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n658), .B1(new_n657), .B2(new_n659), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT102), .B1(new_n655), .B2(G8gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n655), .A2(KEYINPUT102), .A3(G8gat), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI22_X1  g463(.A1(new_n660), .A2(new_n661), .B1(new_n662), .B2(new_n664), .ZN(G1325gat));
  INV_X1    g464(.A(G15gat), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n652), .A2(new_n666), .A3(new_n493), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n608), .A2(new_n651), .A3(new_n507), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n666), .B2(new_n668), .ZN(G1326gat));
  NOR2_X1   g468(.A1(new_n652), .A2(new_n508), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  NAND2_X1  g471(.A1(new_n607), .A2(new_n627), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n524), .A2(new_n650), .A3(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n675), .A2(G29gat), .A3(new_n514), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT45), .Z(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n524), .B2(new_n650), .ZN(new_n679));
  INV_X1    g478(.A(new_n650), .ZN(new_n680));
  AOI211_X1 g479(.A(KEYINPUT44), .B(new_n680), .C1(new_n521), .C2(new_n522), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n674), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G29gat), .B1(new_n682), .B2(new_n514), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n683), .ZN(G1328gat));
  NOR3_X1   g483(.A1(new_n675), .A2(G36gat), .A3(new_n500), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT46), .ZN(new_n686));
  OAI21_X1  g485(.A(G36gat), .B1(new_n682), .B2(new_n500), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(G1329gat));
  INV_X1    g487(.A(KEYINPUT47), .ZN(new_n689));
  INV_X1    g488(.A(G43gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n493), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n674), .B(new_n691), .C1(new_n679), .C2(new_n681), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693));
  INV_X1    g492(.A(new_n507), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n690), .B1(new_n675), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n693), .B1(new_n692), .B2(new_n695), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n689), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n698), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(KEYINPUT47), .A3(new_n696), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(G1330gat));
  INV_X1    g501(.A(G50gat), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n682), .A2(new_n703), .A3(new_n508), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n675), .B2(new_n508), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n704), .A2(KEYINPUT48), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT48), .B1(new_n704), .B2(new_n705), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(G1331gat));
  NAND2_X1  g507(.A1(new_n521), .A2(new_n522), .ZN(new_n709));
  INV_X1    g508(.A(new_n570), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n710), .A2(new_n627), .A3(new_n650), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n606), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n514), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT104), .B(G57gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1332gat));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n712), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n500), .B(KEYINPUT106), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT49), .B(G64gat), .Z(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(G1333gat));
  NOR2_X1   g521(.A1(new_n712), .A2(new_n694), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n573), .ZN(new_n726));
  INV_X1    g525(.A(new_n493), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n717), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G71gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n437), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g533(.A1(new_n679), .A2(new_n681), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n710), .A2(new_n626), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n606), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n514), .A2(new_n583), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n709), .A2(new_n650), .A3(new_n736), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n740), .B2(new_n742), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n499), .A3(new_n606), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n738), .A2(new_n739), .B1(new_n745), .B2(new_n583), .ZN(G1336gat));
  NAND3_X1  g545(.A1(new_n740), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT51), .B1(new_n740), .B2(KEYINPUT109), .ZN(new_n749));
  INV_X1    g548(.A(new_n606), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n752));
  INV_X1    g551(.A(new_n718), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(G92gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n749), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n756), .A2(new_n606), .A3(new_n754), .A4(new_n747), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT110), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n584), .B1(new_n738), .B2(new_n501), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT52), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n744), .A2(new_n606), .A3(new_n754), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n735), .A2(new_n753), .A3(new_n737), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n584), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n761), .A2(new_n765), .ZN(G1337gat));
  INV_X1    g565(.A(G99gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n507), .A2(new_n767), .A3(new_n606), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT111), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n744), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n735), .A2(new_n493), .A3(new_n737), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n767), .ZN(G1338gat));
  INV_X1    g571(.A(new_n737), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n437), .B(new_n773), .C1(new_n679), .C2(new_n681), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G106gat), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n508), .A2(G106gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n744), .A2(new_n606), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n774), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT112), .B1(new_n774), .B2(G106gat), .ZN(new_n781));
  AND4_X1   g580(.A1(new_n606), .A2(new_n756), .A3(new_n747), .A4(new_n777), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n779), .B1(new_n783), .B2(new_n776), .ZN(G1339gat));
  AND2_X1   g583(.A1(new_n548), .A2(new_n550), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n785), .A2(new_n551), .B1(new_n556), .B2(new_n557), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n565), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n569), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT54), .B1(new_n596), .B2(new_n597), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n598), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n605), .B1(new_n598), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(KEYINPUT55), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n598), .A2(new_n789), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n596), .A2(new_n597), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n604), .B1(new_n796), .B2(KEYINPUT54), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n600), .A2(new_n605), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n793), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n650), .A2(new_n788), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n800), .B1(new_n568), .B2(new_n569), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n606), .A2(new_n787), .A3(new_n569), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n680), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n650), .A2(new_n788), .A3(KEYINPUT113), .A4(new_n801), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n627), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n711), .A2(new_n750), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n507), .A3(new_n508), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n514), .A2(new_n718), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G113gat), .B1(new_n816), .B2(new_n570), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n514), .B1(new_n810), .B2(new_n811), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n513), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n753), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n710), .A2(new_n300), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(G1340gat));
  OAI21_X1  g621(.A(G120gat), .B1(new_n816), .B2(new_n750), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n606), .A2(new_n298), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n820), .B2(new_n824), .ZN(G1341gat));
  NOR3_X1   g624(.A1(new_n816), .A2(new_n304), .A3(new_n627), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n819), .A2(new_n626), .A3(new_n753), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n826), .B1(new_n304), .B2(new_n827), .ZN(G1342gat));
  NOR2_X1   g627(.A1(new_n680), .A2(new_n501), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n819), .A2(new_n329), .A3(new_n829), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT56), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n831), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(KEYINPUT115), .B2(KEYINPUT56), .ZN(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n816), .B2(new_n680), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT116), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n831), .A2(new_n833), .A3(new_n834), .A4(new_n832), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(new_n838), .A3(new_n839), .ZN(G1343gat));
  NOR2_X1   g639(.A1(new_n727), .A2(new_n508), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n818), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n753), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(G141gat), .A3(new_n570), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n812), .A2(new_n437), .ZN(new_n845));
  XNOR2_X1  g644(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n812), .A2(new_n848), .A3(new_n437), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n815), .A2(new_n493), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n710), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n844), .B1(new_n340), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n855), .B(new_n856), .ZN(G1344gat));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858));
  AOI211_X1 g657(.A(KEYINPUT59), .B(new_n312), .C1(new_n851), .C2(new_n606), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n807), .A2(new_n802), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n860), .A2(new_n627), .B1(new_n711), .B2(new_n750), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n848), .B1(new_n861), .B2(new_n508), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n812), .A2(new_n437), .A3(new_n846), .ZN(new_n865));
  OAI211_X1 g664(.A(KEYINPUT119), .B(new_n848), .C1(new_n861), .C2(new_n508), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n606), .A3(new_n850), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n867), .A2(KEYINPUT120), .A3(new_n606), .A4(new_n850), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(G148gat), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n859), .B1(new_n872), .B2(KEYINPUT59), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n842), .A2(new_n312), .A3(new_n606), .A4(new_n753), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n858), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n312), .B1(new_n868), .B2(new_n869), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n871), .ZN(new_n879));
  OAI211_X1 g678(.A(KEYINPUT121), .B(new_n874), .C1(new_n879), .C2(new_n859), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n876), .A2(new_n880), .ZN(G1345gat));
  NAND3_X1  g680(.A1(new_n851), .A2(G155gat), .A3(new_n626), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n308), .B1(new_n843), .B2(new_n627), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(G1346gat));
  NAND3_X1  g684(.A1(new_n842), .A2(new_n309), .A3(new_n829), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n851), .A2(new_n650), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n309), .ZN(G1347gat));
  AOI211_X1 g687(.A(new_n499), .B(new_n753), .C1(new_n810), .C2(new_n811), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n513), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n891), .B(new_n710), .C1(new_n220), .C2(new_n221), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n499), .A2(new_n500), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT122), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n814), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n710), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n897), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT123), .B1(new_n897), .B2(G169gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n892), .B1(new_n898), .B2(new_n899), .ZN(G1348gat));
  NOR3_X1   g699(.A1(new_n895), .A2(new_n213), .A3(new_n750), .ZN(new_n901));
  AOI21_X1  g700(.A(G176gat), .B1(new_n891), .B2(new_n606), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(G1349gat));
  OAI21_X1  g702(.A(G183gat), .B1(new_n895), .B2(new_n627), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n891), .A2(new_n626), .A3(new_n239), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT60), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n906), .A2(KEYINPUT60), .ZN(new_n909));
  XOR2_X1   g708(.A(new_n908), .B(new_n909), .Z(G1350gat));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n650), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(G190gat), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT125), .B(new_n208), .C1(new_n896), .C2(new_n650), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  OR3_X1    g714(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n891), .A2(new_n650), .A3(new_n231), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n915), .B1(new_n913), .B2(new_n914), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G1351gat));
  NAND2_X1  g718(.A1(new_n894), .A2(new_n493), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT126), .Z(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n867), .ZN(new_n922));
  OAI21_X1  g721(.A(G197gat), .B1(new_n922), .B2(new_n570), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n889), .A2(new_n841), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(G197gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n923), .B1(new_n570), .B2(new_n925), .ZN(G1352gat));
  NOR3_X1   g725(.A1(new_n924), .A2(G204gat), .A3(new_n750), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT62), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n921), .A2(new_n867), .A3(new_n606), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n603), .B2(new_n929), .ZN(G1353gat));
  OAI21_X1  g729(.A(G211gat), .B1(new_n922), .B2(new_n627), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n931), .A2(KEYINPUT63), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(KEYINPUT63), .ZN(new_n933));
  INV_X1    g732(.A(new_n924), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n253), .A3(new_n626), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT127), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n932), .A2(new_n933), .A3(new_n936), .ZN(G1354gat));
  OAI21_X1  g736(.A(G218gat), .B1(new_n922), .B2(new_n680), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n934), .A2(new_n254), .A3(new_n650), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1355gat));
endmodule


