//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT69), .A2(G116), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT69), .A2(G116), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G119), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(KEYINPUT5), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G113), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT5), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n192), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(KEYINPUT2), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G113), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n190), .A2(new_n193), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G104), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(KEYINPUT77), .A3(G104), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n205), .B1(KEYINPUT3), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT78), .B(G101), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n209), .A2(new_n204), .A3(KEYINPUT77), .A4(G104), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  OAI21_X1  g027(.A(G101), .B1(new_n213), .B2(new_n205), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n198), .A2(new_n203), .A3(new_n211), .A4(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G110), .B(G122), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n206), .A2(KEYINPUT3), .ZN(new_n217));
  INV_X1    g031(.A(new_n205), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n210), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G101), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n211), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n222), .A3(G101), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n202), .B1(new_n190), .B2(new_n193), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n190), .A2(new_n193), .A3(new_n202), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n215), .B(new_n216), .C1(new_n221), .C2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n216), .B(KEYINPUT8), .ZN(new_n228));
  INV_X1    g042(.A(new_n215), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n198), .A2(new_n203), .B1(new_n211), .B2(new_n214), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G224), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(G953), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(KEYINPUT86), .ZN(new_n234));
  XNOR2_X1  g048(.A(G143), .B(G146), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G128), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(G125), .ZN(new_n239));
  INV_X1    g053(.A(G143), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT1), .B1(new_n240), .B2(G146), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT67), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G128), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n241), .A2(KEYINPUT66), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G143), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT1), .ZN(new_n250));
  AOI211_X1 g064(.A(KEYINPUT68), .B(new_n235), .C1(new_n246), .C2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n241), .A2(KEYINPUT66), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n243), .A2(new_n245), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n250), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n240), .A2(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n248), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n252), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n239), .B1(new_n251), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  OR2_X1    g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n257), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n248), .A2(new_n256), .A3(KEYINPUT0), .A4(G128), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G125), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n234), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT7), .B1(new_n232), .B2(G953), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n227), .B(new_n231), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n267), .ZN(new_n269));
  AOI211_X1 g083(.A(new_n269), .B(new_n234), .C1(new_n259), .C2(new_n265), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n187), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n259), .A2(new_n265), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n233), .B(KEYINPUT84), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n259), .A2(new_n265), .A3(new_n273), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n215), .B1(new_n221), .B2(new_n226), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n216), .B(KEYINPUT83), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n227), .A2(KEYINPUT6), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n281));
  INV_X1    g095(.A(new_n279), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n211), .ZN(new_n283));
  INV_X1    g097(.A(new_n224), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n203), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n285), .A3(new_n223), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n281), .B(new_n282), .C1(new_n286), .C2(new_n215), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n277), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT85), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n277), .B(new_n290), .C1(new_n280), .C2(new_n287), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n271), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n293), .B(KEYINPUT87), .Z(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n294), .B(KEYINPUT88), .Z(new_n297));
  OAI21_X1  g111(.A(new_n296), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G214), .B1(G237), .B2(G902), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n188), .A2(G122), .A3(new_n189), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n191), .A2(G122), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT14), .ZN(new_n303));
  OAI21_X1  g117(.A(G107), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n302), .B(new_n304), .Z(new_n305));
  INV_X1    g119(.A(KEYINPUT92), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n243), .A2(new_n245), .A3(G143), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n240), .A2(G128), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n306), .A3(new_n308), .ZN(new_n311));
  AOI21_X1  g125(.A(G134), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n311), .ZN(new_n313));
  INV_X1    g127(.A(G134), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n313), .A2(new_n314), .A3(new_n309), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n305), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT93), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n314), .B1(new_n313), .B2(new_n309), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT93), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n302), .A2(new_n204), .ZN(new_n321));
  OAI21_X1  g135(.A(G107), .B1(new_n300), .B2(new_n301), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT13), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n308), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n240), .A2(KEYINPUT13), .A3(G128), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n307), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n321), .A2(new_n322), .B1(G134), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n318), .A2(new_n320), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT9), .B(G234), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(G217), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n316), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n316), .B2(new_n328), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n187), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT15), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G478), .ZN(new_n338));
  INV_X1    g152(.A(G478), .ZN(new_n339));
  OAI221_X1 g153(.A(new_n187), .B1(KEYINPUT15), .B2(new_n339), .C1(new_n334), .C2(new_n335), .ZN(new_n340));
  INV_X1    g154(.A(G952), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(G953), .ZN(new_n342));
  INV_X1    g156(.A(G234), .ZN(new_n343));
  INV_X1    g157(.A(G237), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n187), .B(new_n331), .C1(G234), .C2(G237), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT21), .B(G898), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n338), .A2(new_n340), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n344), .A2(new_n331), .A3(G214), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n240), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n344), .A2(new_n331), .A3(G143), .A4(G214), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT18), .A3(G131), .ZN(new_n356));
  XOR2_X1   g170(.A(G125), .B(G140), .Z(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G146), .ZN(new_n358));
  XNOR2_X1  g172(.A(G125), .B(G140), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n247), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n355), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT18), .A2(G131), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT89), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT90), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  AND4_X1   g179(.A1(KEYINPUT90), .A2(new_n364), .A3(new_n353), .A4(new_n354), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n356), .B(new_n361), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G113), .B(G122), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(new_n212), .ZN(new_n369));
  INV_X1    g183(.A(G125), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n370), .A2(KEYINPUT16), .A3(G140), .ZN(new_n371));
  AOI211_X1 g185(.A(new_n247), .B(new_n371), .C1(KEYINPUT16), .C2(new_n359), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n371), .B1(new_n359), .B2(KEYINPUT16), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G146), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT73), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n375), .A2(G146), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n355), .A2(G131), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT17), .ZN(new_n382));
  INV_X1    g196(.A(G131), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n353), .A2(new_n383), .A3(new_n354), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n355), .A2(KEYINPUT17), .A3(G131), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n367), .B(new_n369), .C1(new_n380), .C2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n378), .B1(new_n373), .B2(new_n372), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n390), .A2(new_n377), .A3(new_n385), .A4(new_n386), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n369), .B1(new_n391), .B2(new_n367), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n187), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G475), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n359), .A2(KEYINPUT19), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n359), .A2(KEYINPUT19), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n247), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT91), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(new_n376), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT19), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n357), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(G146), .B1(new_n403), .B2(new_n396), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT91), .B1(new_n404), .B2(new_n372), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n381), .A2(new_n384), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n407), .A2(new_n367), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n388), .B1(new_n408), .B2(new_n369), .ZN(new_n409));
  NOR2_X1   g223(.A1(G475), .A2(G902), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n395), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n369), .B1(new_n407), .B2(new_n367), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n395), .B(new_n410), .C1(new_n389), .C2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n394), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n351), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n298), .A2(new_n299), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n262), .A2(KEYINPUT70), .A3(new_n263), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT70), .B1(new_n262), .B2(new_n263), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n223), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT79), .B1(new_n421), .B2(new_n221), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT70), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n264), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n262), .A2(KEYINPUT70), .A3(new_n263), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT79), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n283), .A4(new_n223), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G137), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G134), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT11), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(KEYINPUT11), .A3(G134), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n314), .A2(G137), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n383), .A2(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT10), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n237), .B1(new_n251), .B2(new_n258), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n211), .A2(new_n214), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n440), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n237), .A2(KEYINPUT80), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n241), .A2(G128), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n237), .A2(KEYINPUT80), .B1(new_n257), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n440), .A3(new_n443), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n429), .B(new_n439), .C1(new_n444), .C2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G140), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n331), .A2(G227), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n429), .B1(new_n444), .B2(new_n450), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT81), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n438), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n255), .A2(new_n257), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT68), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n255), .A2(new_n252), .A3(new_n257), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n238), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT10), .B1(new_n463), .B2(new_n442), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n464), .A2(new_n449), .B1(new_n422), .B2(new_n428), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT81), .B1(new_n465), .B2(new_n439), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n456), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n448), .A2(new_n443), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n441), .B2(new_n443), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n438), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT12), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(KEYINPUT12), .A3(new_n438), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n455), .B1(new_n474), .B2(new_n451), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT82), .B1(new_n467), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n454), .B1(new_n465), .B2(new_n439), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n465), .A2(KEYINPUT81), .A3(new_n439), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n458), .B1(new_n457), .B2(new_n438), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT82), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n474), .A2(new_n451), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n454), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n476), .A2(new_n484), .A3(G469), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n477), .A2(new_n474), .ZN(new_n486));
  INV_X1    g300(.A(new_n451), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n466), .B2(new_n459), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n488), .B2(new_n455), .ZN(new_n489));
  INV_X1    g303(.A(G469), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(new_n187), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n187), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n485), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G221), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(new_n330), .B2(new_n187), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n418), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n426), .A2(new_n438), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n435), .A2(G131), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(KEYINPUT65), .B2(new_n431), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(KEYINPUT65), .B2(new_n431), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n436), .A2(new_n383), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n499), .B(KEYINPUT30), .C1(new_n463), .C2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n264), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n441), .A2(new_n504), .B1(new_n438), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n506), .B(new_n285), .C1(KEYINPUT30), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n344), .A2(new_n331), .A3(G210), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n510), .B(KEYINPUT27), .Z(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G101), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n441), .A2(new_n504), .B1(new_n438), .B2(new_n426), .ZN(new_n515));
  INV_X1    g329(.A(new_n285), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n509), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT31), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT28), .ZN(new_n520));
  OAI22_X1  g334(.A1(new_n517), .A2(new_n520), .B1(new_n516), .B2(new_n508), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT28), .B1(new_n515), .B2(new_n516), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n513), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT31), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n509), .A2(new_n524), .A3(new_n514), .A4(new_n517), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(G472), .A2(G902), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT32), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n441), .A2(new_n504), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n499), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n285), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n517), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT28), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT71), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n522), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n522), .A2(new_n536), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n514), .A2(KEYINPUT29), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n535), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n187), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n514), .B1(new_n521), .B2(new_n522), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n509), .A2(new_n513), .A3(new_n517), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT29), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G472), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n526), .A2(KEYINPUT32), .A3(new_n527), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n530), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n548));
  INV_X1    g362(.A(G110), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT67), .B(G128), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT23), .A3(G119), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT23), .B1(new_n242), .B2(G119), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n242), .A2(G119), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n549), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n550), .B2(G119), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT24), .B(G110), .Z(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n380), .A2(new_n558), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n551), .A2(new_n554), .A3(new_n549), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n556), .A2(new_n557), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n376), .B(new_n360), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT22), .B(G137), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n495), .A2(new_n343), .A3(G953), .ZN(new_n565));
  XOR2_X1   g379(.A(new_n564), .B(new_n565), .Z(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(KEYINPUT74), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n559), .A2(new_n570), .A3(new_n562), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n566), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n548), .B1(new_n574), .B2(G902), .ZN(new_n575));
  INV_X1    g389(.A(new_n571), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n570), .B1(new_n559), .B2(new_n562), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n567), .ZN(new_n579));
  INV_X1    g393(.A(new_n548), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n187), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(G217), .B1(new_n343), .B2(G902), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n583), .B(KEYINPUT72), .Z(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n187), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n582), .A2(new_n585), .B1(new_n579), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n547), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT76), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n547), .A2(KEYINPUT76), .A3(new_n588), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n498), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n208), .ZN(G3));
  NAND2_X1  g408(.A1(new_n289), .A2(new_n291), .ZN(new_n595));
  INV_X1    g409(.A(new_n271), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n295), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI211_X1 g411(.A(new_n294), .B(new_n271), .C1(new_n289), .C2(new_n291), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n299), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT94), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n187), .A2(G478), .ZN(new_n601));
  INV_X1    g415(.A(new_n335), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n316), .A2(new_n328), .A3(new_n333), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT33), .B1(new_n334), .B2(new_n335), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT95), .B(G478), .Z(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n336), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n415), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n613), .B(new_n299), .C1(new_n597), .C2(new_n598), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n600), .A2(new_n350), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n494), .A2(new_n497), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n526), .A2(new_n187), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G472), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n588), .A2(new_n528), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NOR2_X1   g437(.A1(new_n394), .A2(KEYINPUT96), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n393), .B2(G475), .ZN(new_n626));
  OAI22_X1  g440(.A1(new_n624), .A2(new_n626), .B1(new_n411), .B2(new_n414), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n338), .A2(new_n340), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n600), .A2(new_n350), .A3(new_n614), .A4(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(KEYINPUT97), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(KEYINPUT97), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n617), .B(new_n620), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  AOI21_X1  g450(.A(new_n580), .B1(new_n579), .B2(new_n187), .ZN(new_n637));
  AOI211_X1 g451(.A(G902), .B(new_n548), .C1(new_n578), .C2(new_n567), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n585), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n572), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT98), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n640), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n587), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n645), .A2(new_n619), .A3(new_n528), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n646), .A2(new_n418), .A3(new_n497), .A4(new_n494), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT37), .B(G110), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(G12));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n346), .B1(new_n347), .B2(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n627), .A2(new_n629), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n600), .A2(new_n614), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT100), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n547), .A2(new_n645), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n600), .A2(new_n657), .A3(new_n614), .A4(new_n653), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n655), .A2(new_n617), .A3(new_n656), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XOR2_X1   g474(.A(new_n652), .B(KEYINPUT39), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n617), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n298), .B(KEYINPUT38), .ZN(new_n665));
  INV_X1    g479(.A(new_n299), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n410), .B1(new_n389), .B2(new_n412), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT20), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n668), .A2(new_n413), .B1(G475), .B2(new_n393), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n645), .A2(new_n666), .A3(new_n669), .A4(new_n629), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n509), .A2(new_n517), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n514), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n672), .B(new_n187), .C1(new_n514), .C2(new_n534), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n528), .A2(new_n529), .B1(G472), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n546), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n665), .A2(new_n670), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n663), .A2(new_n664), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  NOR2_X1   g492(.A1(new_n611), .A2(new_n652), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n600), .A2(new_n614), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n617), .A3(KEYINPUT101), .A4(new_n656), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n494), .A2(new_n547), .A3(new_n497), .A4(new_n645), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n683), .B1(new_n684), .B2(new_n680), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  INV_X1    g501(.A(new_n589), .ZN(new_n688));
  INV_X1    g502(.A(new_n491), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n490), .B1(new_n489), .B2(new_n187), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n689), .A2(new_n690), .A3(new_n496), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT102), .B1(new_n692), .B2(new_n615), .ZN(new_n693));
  INV_X1    g507(.A(new_n690), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n497), .A3(new_n491), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n589), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n616), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT103), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n699), .B(new_n701), .ZN(G15));
  OAI21_X1  g516(.A(new_n696), .B1(new_n632), .B2(new_n633), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  NAND3_X1  g520(.A1(new_n691), .A2(new_n614), .A3(new_n600), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n547), .A2(new_n416), .A3(new_n645), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(G119), .Z(G21));
  XOR2_X1   g524(.A(new_n527), .B(KEYINPUT105), .Z(new_n711));
  AND2_X1   g525(.A1(new_n535), .A2(new_n538), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n514), .B1(new_n712), .B2(new_n537), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n519), .A2(new_n525), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(new_n619), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n691), .A2(new_n588), .A3(new_n350), .A4(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n629), .A2(new_n669), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n600), .A2(new_n614), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT106), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n588), .A2(new_n715), .A3(new_n619), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n695), .A2(new_n721), .A3(new_n349), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n600), .A2(new_n614), .A3(new_n718), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  AND4_X1   g541(.A1(new_n619), .A2(new_n679), .A3(new_n715), .A4(new_n645), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n691), .A3(new_n614), .A4(new_n600), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  NAND2_X1  g544(.A1(new_n530), .A2(KEYINPUT108), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n546), .A3(new_n545), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n530), .A2(KEYINPUT108), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n588), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OR3_X1    g548(.A1(new_n298), .A2(KEYINPUT107), .A3(new_n666), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n467), .A2(new_n475), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n492), .B1(new_n736), .B2(G469), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n496), .B1(new_n737), .B2(new_n491), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT107), .B1(new_n298), .B2(new_n666), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n735), .A2(new_n679), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT42), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n735), .A2(new_n739), .A3(new_n738), .ZN(new_n742));
  INV_X1    g556(.A(new_n679), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(KEYINPUT42), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n688), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n383), .ZN(G33));
  NAND3_X1  g561(.A1(new_n742), .A2(new_n688), .A3(new_n653), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  NAND2_X1  g563(.A1(new_n735), .A2(new_n739), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n619), .A2(new_n528), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n645), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT110), .Z(new_n754));
  OR2_X1    g568(.A1(new_n607), .A2(new_n610), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n669), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT43), .Z(new_n757));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n751), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n759), .B2(new_n758), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n736), .A2(KEYINPUT45), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(G469), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT45), .B1(new_n476), .B2(new_n484), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n762), .B1(new_n766), .B2(new_n492), .ZN(new_n767));
  OAI211_X1 g581(.A(KEYINPUT46), .B(new_n493), .C1(new_n764), .C2(new_n765), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n491), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n497), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n771), .A2(new_n772), .A3(new_n661), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n772), .B1(new_n771), .B2(new_n661), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n761), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT111), .B(G137), .Z(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G39));
  NOR4_X1   g591(.A1(new_n750), .A2(new_n547), .A3(new_n588), .A4(new_n743), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n771), .A2(KEYINPUT47), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n771), .A2(KEYINPUT47), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n617), .A2(new_n656), .A3(new_n658), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n654), .A2(KEYINPUT100), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n716), .A2(new_n645), .A3(new_n679), .ZN(new_n787));
  INV_X1    g601(.A(new_n652), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n639), .A2(new_n644), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n674), .B2(new_n546), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n738), .ZN(new_n791));
  OAI22_X1  g605(.A1(new_n707), .A2(new_n787), .B1(new_n791), .B2(new_n719), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n786), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT114), .B1(new_n793), .B2(new_n686), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n599), .A2(KEYINPUT94), .ZN(new_n795));
  INV_X1    g609(.A(new_n614), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n695), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n789), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n738), .A2(new_n675), .A3(new_n798), .ZN(new_n799));
  AOI22_X1  g613(.A1(new_n797), .A2(new_n728), .B1(new_n799), .B2(new_n724), .ZN(new_n800));
  AND4_X1   g614(.A1(KEYINPUT114), .A2(new_n686), .A3(new_n659), .A4(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n783), .B1(new_n794), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n682), .A2(new_n685), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n724), .A2(new_n738), .A3(new_n790), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n729), .B(new_n805), .C1(new_n784), .C2(new_n785), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n686), .A2(new_n800), .A3(KEYINPUT114), .A4(new_n659), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(KEYINPUT52), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n802), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n628), .A2(new_n669), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n611), .A2(new_n811), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n299), .A2(new_n812), .A3(new_n298), .A4(new_n350), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(new_n620), .A3(new_n497), .A4(new_n494), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n814), .B(new_n647), .C1(new_n707), .C2(new_n708), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n593), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n816), .A2(new_n699), .A3(new_n726), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n741), .A2(new_n745), .A3(new_n748), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n742), .A2(new_n728), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n627), .A2(new_n628), .A3(new_n652), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT113), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n751), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n819), .B1(new_n822), .B2(new_n684), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n817), .A2(new_n705), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n810), .A2(KEYINPUT53), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT117), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n817), .A2(new_n705), .A3(new_n824), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n802), .B2(new_n809), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT53), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n659), .A2(new_n729), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(new_n686), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(KEYINPUT52), .A3(new_n805), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(new_n807), .B2(new_n808), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g651(.A(KEYINPUT115), .B(KEYINPUT52), .C1(new_n807), .C2(new_n808), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT116), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n802), .A2(KEYINPUT115), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n835), .A2(new_n836), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n834), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n828), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n827), .B(new_n831), .C1(new_n844), .C2(KEYINPUT53), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT54), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n828), .A2(new_n847), .ZN(new_n848));
  AND4_X1   g662(.A1(KEYINPUT52), .A2(new_n832), .A3(new_n686), .A4(new_n805), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n802), .B2(KEYINPUT115), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n841), .B1(new_n850), .B2(new_n842), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n837), .A2(KEYINPUT116), .A3(new_n838), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n829), .A2(KEYINPUT53), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n853), .A2(KEYINPUT118), .A3(new_n854), .A4(new_n856), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n750), .A2(new_n695), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n346), .A3(new_n757), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n734), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT48), .ZN(new_n864));
  INV_X1    g678(.A(new_n588), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n675), .A2(new_n865), .A3(new_n345), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n611), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n757), .A2(new_n346), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n721), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n342), .B1(new_n871), .B2(new_n707), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n864), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  OR3_X1    g687(.A1(new_n867), .A2(new_n415), .A3(new_n755), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n716), .A2(new_n645), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n665), .A2(new_n695), .A3(new_n299), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n870), .A2(KEYINPUT50), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT50), .B1(new_n870), .B2(new_n876), .ZN(new_n878));
  OAI221_X1 g692(.A(new_n874), .B1(new_n875), .B2(new_n862), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n779), .A2(new_n780), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n689), .A2(new_n690), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n497), .B2(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n869), .A2(new_n721), .A3(new_n750), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n879), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n873), .B1(new_n885), .B2(KEYINPUT51), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(KEYINPUT51), .B2(new_n885), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n846), .A2(new_n859), .A3(new_n860), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n341), .A2(new_n331), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n755), .A2(new_n497), .A3(new_n299), .A4(new_n669), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n865), .B(new_n891), .C1(new_n882), .C2(KEYINPUT49), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT112), .Z(new_n893));
  NOR2_X1   g707(.A1(new_n665), .A2(new_n675), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n893), .B(new_n894), .C1(KEYINPUT49), .C2(new_n882), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n890), .A2(new_n895), .ZN(G75));
  AOI21_X1  g710(.A(new_n282), .B1(new_n286), .B2(new_n215), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT6), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n227), .A2(KEYINPUT6), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(new_n897), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n277), .ZN(new_n901));
  XOR2_X1   g715(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n187), .B1(new_n853), .B2(new_n856), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n294), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n331), .A2(G952), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n903), .A2(new_n906), .ZN(new_n909));
  INV_X1    g723(.A(new_n297), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(G51));
  XNOR2_X1  g726(.A(new_n492), .B(KEYINPUT57), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n854), .B1(new_n853), .B2(new_n856), .ZN(new_n914));
  INV_X1    g728(.A(new_n848), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n839), .B2(new_n843), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n916), .A2(KEYINPUT54), .A3(new_n855), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n913), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n489), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n904), .A2(new_n766), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n908), .B1(new_n919), .B2(new_n920), .ZN(G54));
  NAND3_X1  g735(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  INV_X1    g736(.A(new_n409), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n908), .ZN(G60));
  AND2_X1   g740(.A1(new_n605), .A2(new_n606), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n914), .B2(new_n917), .ZN(new_n931));
  INV_X1    g745(.A(new_n908), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n929), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n827), .A2(new_n831), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n825), .B1(new_n851), .B2(new_n852), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n847), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n860), .B1(new_n937), .B2(new_n854), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n917), .A2(KEYINPUT118), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n933), .B1(new_n940), .B2(new_n927), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n643), .B(new_n944), .C1(new_n916), .C2(new_n855), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n853), .B2(new_n856), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n932), .B(new_n945), .C1(new_n946), .C2(new_n579), .ZN(new_n947));
  NAND2_X1  g761(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n947), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n944), .B1(new_n916), .B2(new_n855), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n908), .B1(new_n953), .B2(new_n574), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(new_n949), .A3(new_n950), .A4(new_n945), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n952), .A2(new_n955), .ZN(G66));
  OAI21_X1  g770(.A(G953), .B1(new_n348), .B2(new_n232), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n817), .A2(new_n705), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT121), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n959), .B2(G953), .ZN(new_n960));
  INV_X1    g774(.A(new_n900), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(G898), .B2(new_n331), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n960), .B(new_n962), .ZN(G69));
  OAI21_X1  g777(.A(new_n506), .B1(new_n508), .B2(KEYINPUT30), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n403), .A2(new_n396), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT122), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n833), .A2(new_n677), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT123), .Z(new_n970));
  INV_X1    g784(.A(new_n662), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n591), .A2(new_n592), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n971), .A2(new_n972), .A3(new_n751), .A4(new_n812), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n974));
  AND4_X1   g788(.A1(new_n775), .A2(new_n781), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n967), .B1(new_n976), .B2(new_n331), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n734), .A2(new_n719), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n773), .B2(new_n774), .ZN(new_n979));
  INV_X1    g793(.A(new_n833), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(new_n818), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n775), .A2(new_n979), .A3(new_n781), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n331), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n966), .B1(G900), .B2(G953), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT124), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n977), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n331), .B1(G227), .B2(G900), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n987), .B(new_n989), .ZN(G72));
  NAND3_X1  g804(.A1(new_n970), .A2(new_n959), .A3(new_n975), .ZN(new_n991));
  XNOR2_X1  g805(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n992));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n672), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n994), .B1(new_n982), .B2(new_n959), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n932), .B1(new_n997), .B2(new_n543), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(KEYINPUT126), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n1000), .B(new_n932), .C1(new_n997), .C2(new_n543), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n996), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n845), .A2(new_n543), .A3(new_n672), .A4(new_n995), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n1002), .A2(new_n1003), .ZN(G57));
endmodule


