//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932;
  NOR2_X1   g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT14), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G43gat), .B(G50gat), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  OAI221_X1 g006(.A(new_n204), .B1(KEYINPUT15), .B2(new_n205), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(KEYINPUT15), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n208), .B(new_n209), .Z(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT17), .ZN(new_n211));
  XNOR2_X1  g010(.A(G15gat), .B(G22gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(G1gat), .ZN(new_n213));
  AOI21_X1  g012(.A(G8gat), .B1(new_n213), .B2(KEYINPUT96), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n215), .A2(KEYINPUT95), .A3(G1gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT95), .B1(new_n215), .B2(G1gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n213), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n219), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT97), .ZN(new_n223));
  INV_X1    g022(.A(new_n222), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n211), .A2(new_n223), .B1(new_n224), .B2(new_n210), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT18), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT99), .ZN(new_n230));
  XNOR2_X1  g029(.A(G113gat), .B(G141gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT11), .ZN(new_n232));
  INV_X1    g031(.A(G169gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(G197gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT12), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n225), .A2(KEYINPUT18), .A3(new_n226), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT98), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n224), .B(new_n210), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n226), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n239), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n237), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n236), .ZN(new_n247));
  INV_X1    g046(.A(new_n229), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT94), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT74), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  INV_X1    g053(.A(G113gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(G120gat), .ZN(new_n256));
  INV_X1    g055(.A(G120gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(G113gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n254), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G127gat), .B(G134gat), .Z(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(KEYINPUT67), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(G113gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(G120gat), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G127gat), .B(G134gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n261), .A2(new_n267), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n274), .B1(new_n275), .B2(KEYINPUT24), .ZN(new_n276));
  INV_X1    g075(.A(G183gat), .ZN(new_n277));
  INV_X1    g076(.A(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n275), .A2(KEYINPUT24), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT23), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(KEYINPUT64), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n281), .A2(KEYINPUT25), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT25), .B1(new_n281), .B2(new_n286), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n277), .A2(KEYINPUT27), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G183gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n293), .A3(new_n278), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT28), .B1(new_n294), .B2(KEYINPUT65), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n291), .A2(new_n293), .A3(new_n296), .A4(new_n278), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n295), .A2(KEYINPUT66), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT66), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n274), .ZN(new_n304));
  NOR3_X1   g103(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n275), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n273), .B(new_n290), .C1(new_n302), .C2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT65), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(new_n300), .A3(new_n297), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT66), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n295), .A2(KEYINPUT66), .A3(new_n297), .ZN(new_n314));
  INV_X1    g113(.A(new_n301), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n306), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n289), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(KEYINPUT69), .A3(new_n273), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n317), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n290), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n261), .A2(new_n267), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n268), .A2(new_n272), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n319), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G227gat), .ZN(new_n327));
  INV_X1    g126(.A(G233gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n253), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT34), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n326), .A2(new_n329), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT32), .ZN(new_n333));
  XNOR2_X1  g132(.A(G15gat), .B(G43gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G71gat), .B(G99gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT33), .B1(new_n337), .B2(KEYINPUT72), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(KEYINPUT72), .B2(new_n337), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT71), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT70), .ZN(new_n343));
  INV_X1    g142(.A(new_n329), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT69), .B1(new_n318), .B2(new_n273), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n318), .A2(new_n273), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n344), .B1(new_n347), .B2(new_n319), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT32), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n343), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n332), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT33), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n336), .B1(new_n332), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n342), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT70), .B1(new_n332), .B2(KEYINPUT32), .ZN(new_n356));
  AOI211_X1 g155(.A(new_n343), .B(new_n349), .C1(new_n326), .C2(new_n329), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n342), .B(new_n354), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n341), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT71), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n340), .B1(new_n364), .B2(new_n358), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT73), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n331), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n331), .B(new_n341), .C1(new_n355), .C2(new_n359), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n369), .A2(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(new_n369), .B2(KEYINPUT22), .ZN(new_n371));
  XNOR2_X1  g170(.A(G197gat), .B(G204gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G211gat), .B(G218gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT2), .ZN(new_n377));
  INV_X1    g176(.A(G148gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G141gat), .ZN(new_n379));
  INV_X1    g178(.A(G141gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(G148gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383));
  OR3_X1    g182(.A1(KEYINPUT81), .A2(G155gat), .A3(G162gat), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n378), .B2(G141gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n378), .A2(G141gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n380), .A2(KEYINPUT82), .A3(G148gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G155gat), .B(G162gat), .ZN(new_n392));
  INV_X1    g191(.A(G155gat), .ZN(new_n393));
  INV_X1    g192(.A(G162gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT83), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G162gat), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n393), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n391), .B(new_n392), .C1(new_n398), .C2(new_n377), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n386), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n376), .B1(new_n404), .B2(KEYINPUT88), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(KEYINPUT88), .B2(new_n404), .ZN(new_n406));
  INV_X1    g205(.A(G228gat), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n401), .B1(new_n375), .B2(KEYINPUT29), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n386), .A2(new_n399), .ZN(new_n409));
  AOI211_X1 g208(.A(new_n407), .B(new_n328), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n374), .B1(new_n371), .B2(new_n372), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT29), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n414), .B1(new_n376), .B2(new_n413), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n409), .A2(KEYINPUT84), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT84), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n386), .A2(new_n399), .A3(new_n417), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n415), .A2(new_n401), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n376), .B1(new_n403), .B2(new_n402), .ZN(new_n420));
  OAI22_X1  g219(.A1(new_n419), .A2(new_n420), .B1(new_n407), .B2(new_n328), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT31), .B(G50gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n411), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n421), .B2(new_n411), .ZN(new_n425));
  XNOR2_X1  g224(.A(G78gat), .B(G106gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(G22gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  OR3_X1    g227(.A1(new_n424), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n428), .B1(new_n424), .B2(new_n425), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n368), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n252), .B1(new_n367), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G226gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(new_n328), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n321), .B2(new_n403), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n301), .B1(new_n311), .B2(new_n312), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n306), .B1(new_n437), .B2(new_n314), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n435), .B1(new_n438), .B2(new_n289), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n375), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT29), .B1(new_n320), .B2(new_n290), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n376), .B(new_n439), .C1(new_n443), .C2(new_n435), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G8gat), .B(G36gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(G64gat), .ZN(new_n447));
  INV_X1    g246(.A(G92gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n449), .B(KEYINPUT79), .Z(new_n450));
  OAI211_X1 g249(.A(KEYINPUT78), .B(new_n375), .C1(new_n436), .C2(new_n440), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n445), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT80), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n444), .A2(new_n442), .ZN(new_n455));
  OAI22_X1  g254(.A1(new_n318), .A2(KEYINPUT29), .B1(new_n434), .B2(new_n328), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n376), .B1(new_n456), .B2(new_n439), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n451), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n449), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT30), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n451), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(KEYINPUT30), .A3(new_n449), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n454), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G225gat), .A2(G233gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n324), .A2(new_n409), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n400), .A2(new_n273), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT5), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT86), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n466), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n324), .A2(new_n409), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n400), .A2(new_n273), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT86), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n416), .A2(new_n418), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT4), .B1(new_n478), .B2(new_n324), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT4), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n473), .A2(KEYINPUT85), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n468), .B2(KEYINPUT4), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n409), .A2(KEYINPUT3), .B1(new_n322), .B2(new_n323), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n472), .B1(new_n485), .B2(new_n402), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n471), .A2(new_n477), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n416), .A2(new_n480), .A3(new_n273), .A4(new_n418), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT4), .B1(new_n324), .B2(new_n409), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(new_n470), .A3(new_n486), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G1gat), .B(G29gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(KEYINPUT0), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(G57gat), .ZN(new_n496));
  INV_X1    g295(.A(G85gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT6), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(new_n498), .B2(new_n493), .ZN(new_n500));
  INV_X1    g299(.A(new_n498), .ZN(new_n501));
  OAI211_X1 g300(.A(KEYINPUT6), .B(new_n501), .C1(new_n487), .C2(new_n492), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n465), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n331), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n365), .A2(KEYINPUT73), .ZN(new_n507));
  AOI211_X1 g306(.A(new_n361), .B(new_n340), .C1(new_n364), .C2(new_n358), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n432), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(KEYINPUT94), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n433), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n368), .A2(KEYINPUT75), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT75), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n365), .A2(new_n515), .A3(new_n331), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT76), .B1(new_n365), .B2(new_n331), .ZN(new_n518));
  OR3_X1    g317(.A1(new_n365), .A2(KEYINPUT76), .A3(new_n331), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n487), .A2(KEYINPUT91), .A3(new_n492), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n477), .A2(new_n471), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n484), .A2(new_n486), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n522), .B1(new_n525), .B2(new_n491), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n501), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n499), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n528), .A2(new_n502), .ZN(new_n529));
  INV_X1    g328(.A(new_n431), .ZN(new_n530));
  NOR4_X1   g329(.A1(new_n465), .A2(new_n529), .A3(new_n530), .A4(KEYINPUT35), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n520), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n530), .B1(new_n465), .B2(new_n504), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT37), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n463), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT38), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n450), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n441), .A2(new_n444), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(KEYINPUT37), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n528), .A2(new_n502), .A3(new_n541), .A4(new_n460), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n458), .A2(new_n459), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n449), .B1(new_n543), .B2(KEYINPUT37), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n537), .B1(new_n544), .B2(new_n536), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n431), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n485), .A2(new_n402), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n490), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(KEYINPUT89), .A3(new_n472), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT89), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n488), .A2(new_n489), .B1(new_n402), .B2(new_n485), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(new_n466), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT39), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n473), .A2(new_n474), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n554), .B1(new_n555), .B2(new_n466), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n550), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n498), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT39), .B1(new_n550), .B2(new_n553), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n547), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT40), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n547), .B(KEYINPUT40), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n452), .B(KEYINPUT80), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n462), .A2(new_n464), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n527), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT92), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n465), .A2(KEYINPUT92), .A3(new_n527), .A4(new_n564), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n546), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n534), .B1(new_n571), .B2(KEYINPUT93), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT93), .ZN(new_n573));
  AOI211_X1 g372(.A(new_n573), .B(new_n546), .C1(new_n569), .C2(new_n570), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n368), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT36), .B1(new_n367), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT36), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n517), .A2(new_n578), .A3(new_n519), .A4(new_n518), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n251), .B1(new_n533), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT7), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n497), .B2(new_n448), .ZN(new_n587));
  XNOR2_X1  g386(.A(G99gat), .B(G106gat), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n585), .B(new_n587), .C1(KEYINPUT103), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(KEYINPUT103), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n211), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G190gat), .B(G218gat), .Z(new_n594));
  INV_X1    g393(.A(KEYINPUT104), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT41), .ZN(new_n596));
  NAND2_X1  g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597));
  OAI22_X1  g396(.A1(new_n594), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n598), .B1(new_n210), .B2(new_n591), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n595), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G134gat), .B(G162gat), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n596), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT21), .ZN(new_n609));
  INV_X1    g408(.A(G71gat), .ZN(new_n610));
  INV_X1    g409(.A(G78gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(G71gat), .B2(G78gat), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT100), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  XOR2_X1   g418(.A(G57gat), .B(G64gat), .Z(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(KEYINPUT9), .B2(new_n612), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT9), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n623), .A2(G71gat), .A3(G78gat), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n620), .B1(new_n612), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n222), .B1(new_n609), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G183gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT102), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n628), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n626), .A2(new_n609), .ZN(new_n634));
  XOR2_X1   g433(.A(G127gat), .B(G155gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(G211gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n608), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n591), .B(new_n626), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n646), .B2(KEYINPUT10), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(KEYINPUT105), .A3(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n591), .A2(KEYINPUT10), .A3(new_n625), .A4(new_n622), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n652), .B2(new_n645), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G176gat), .ZN(new_n656));
  INV_X1    g455(.A(G204gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n654), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n643), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n583), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n503), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(G1gat), .Z(G1324gat));
  INV_X1    g465(.A(new_n465), .ZN(new_n667));
  OAI21_X1  g466(.A(G8gat), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT106), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  NAND4_X1  g469(.A1(new_n583), .A2(new_n465), .A3(new_n663), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT42), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n664), .B2(new_n581), .ZN(new_n674));
  INV_X1    g473(.A(G15gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n520), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n664), .B2(new_n676), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n664), .A2(new_n431), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  NOR2_X1   g479(.A1(new_n662), .A2(new_n642), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n608), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n583), .A2(new_n206), .A3(new_n504), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n533), .A2(KEYINPUT107), .A3(new_n582), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n512), .A2(KEYINPUT35), .B1(new_n520), .B2(new_n531), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n580), .A2(new_n572), .A3(new_n574), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n608), .A2(KEYINPUT44), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n686), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n608), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n688), .B2(new_n689), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT44), .ZN(new_n695));
  AOI211_X1 g494(.A(new_n251), .B(new_n682), .C1(new_n692), .C2(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(new_n504), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n685), .B1(new_n697), .B2(new_n206), .ZN(G1328gat));
  AOI21_X1  g497(.A(new_n207), .B1(new_n696), .B2(new_n465), .ZN(new_n699));
  AOI21_X1  g498(.A(G36gat), .B1(KEYINPUT108), .B2(KEYINPUT46), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n583), .A2(new_n465), .A3(new_n683), .A4(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n701), .B(new_n702), .Z(new_n703));
  NOR2_X1   g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1329gat));
  INV_X1    g505(.A(G43gat), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n583), .A2(new_n707), .A3(new_n520), .A4(new_n683), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n696), .A2(new_n580), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(G43gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n711), .B(new_n712), .Z(G1330gat));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n530), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n431), .A2(G50gat), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(KEYINPUT111), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(KEYINPUT111), .ZN(new_n717));
  NOR4_X1   g516(.A1(new_n682), .A2(new_n716), .A3(new_n717), .A4(new_n608), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n714), .A2(G50gat), .B1(new_n583), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g519(.A1(new_n686), .A2(new_n690), .ZN(new_n721));
  INV_X1    g520(.A(new_n662), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n250), .A2(new_n643), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n504), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g526(.A1(new_n724), .A2(new_n667), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  AND2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n728), .B2(new_n729), .ZN(G1333gat));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733));
  OAI21_X1  g532(.A(G71gat), .B1(new_n724), .B2(new_n581), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n721), .A2(new_n610), .A3(new_n520), .A4(new_n723), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n734), .A2(new_n733), .A3(new_n735), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT50), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n738), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n740), .A2(new_n736), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n739), .A2(new_n742), .ZN(G1334gat));
  NOR2_X1   g542(.A1(new_n724), .A2(new_n431), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(new_n611), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n503), .A2(G85gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n251), .A2(new_n641), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT113), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n694), .B2(KEYINPUT115), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n693), .C1(new_n688), .C2(new_n689), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n750), .A2(KEYINPUT51), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT51), .B1(new_n750), .B2(new_n752), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n662), .B(new_n746), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n692), .A2(new_n695), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n748), .A2(new_n662), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n756), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  AOI211_X1 g559(.A(KEYINPUT114), .B(new_n758), .C1(new_n692), .C2(new_n695), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n760), .A2(new_n761), .A3(new_n503), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n755), .B1(new_n762), .B2(new_n497), .ZN(G1336gat));
  NOR2_X1   g562(.A1(new_n667), .A2(G92gat), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n662), .B(new_n764), .C1(new_n753), .C2(new_n754), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n757), .A2(new_n759), .ZN(new_n766));
  OAI21_X1  g565(.A(G92gat), .B1(new_n766), .B2(new_n667), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n760), .A2(new_n761), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n465), .ZN(new_n771));
  NOR2_X1   g570(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n750), .A2(new_n752), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n750), .B2(new_n752), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n722), .A2(G92gat), .A3(new_n667), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n771), .A2(G92gat), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n769), .B1(new_n778), .B2(new_n768), .ZN(G1337gat));
  INV_X1    g578(.A(G99gat), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n581), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n520), .B(new_n662), .C1(new_n753), .C2(new_n754), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n770), .A2(new_n781), .B1(new_n782), .B2(new_n780), .ZN(G1338gat));
  NOR3_X1   g582(.A1(new_n722), .A2(G106gat), .A3(new_n431), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n774), .B2(new_n775), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(KEYINPUT118), .B(new_n784), .C1(new_n774), .C2(new_n775), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT117), .B(G106gat), .Z(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n770), .B2(new_n530), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT53), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n784), .B1(new_n753), .B2(new_n754), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n766), .A2(new_n431), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n793), .B(new_n794), .C1(new_n795), .C2(new_n790), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(G1339gat));
  NOR2_X1   g596(.A1(new_n653), .A2(KEYINPUT54), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(new_n658), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n651), .A2(new_n652), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(KEYINPUT54), .A3(new_n653), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT55), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n804), .A2(new_n660), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n805), .B(new_n250), .C1(KEYINPUT55), .C2(new_n803), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n225), .A2(new_n226), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n241), .A2(new_n242), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n235), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n246), .A2(new_n662), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n693), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n246), .A2(new_n693), .A3(new_n809), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n803), .A2(KEYINPUT55), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n804), .A2(new_n660), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n641), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n251), .A2(new_n663), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n433), .A2(new_n511), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n465), .A2(new_n503), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n250), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n431), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n520), .A2(new_n820), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n251), .A2(new_n255), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(G1340gat));
  AOI21_X1  g626(.A(G120gat), .B1(new_n821), .B2(new_n662), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n722), .A2(new_n257), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n825), .B2(new_n829), .ZN(G1341gat));
  INV_X1    g629(.A(G127gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n821), .A2(new_n831), .A3(new_n642), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n823), .A2(new_n641), .A3(new_n824), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n831), .B2(new_n833), .ZN(G1342gat));
  INV_X1    g633(.A(G134gat), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n825), .B2(new_n693), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT119), .Z(new_n837));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n835), .A3(new_n693), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT56), .Z(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(G1343gat));
  NAND2_X1  g639(.A1(new_n818), .A2(new_n530), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n581), .A2(new_n820), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n380), .A3(new_n250), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT55), .B1(new_n802), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n845), .B2(new_n802), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n805), .A2(new_n250), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n693), .B1(new_n848), .B2(new_n810), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n641), .B1(new_n849), .B2(new_n815), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n850), .A2(new_n851), .B1(new_n251), .B2(new_n663), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n431), .A2(new_n854), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n853), .A2(new_n855), .B1(new_n841), .B2(new_n854), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(new_n251), .A3(new_n842), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n844), .B1(new_n857), .B2(new_n380), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT58), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(new_n844), .C1(new_n857), .C2(new_n380), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1344gat));
  NAND3_X1  g661(.A1(new_n843), .A2(new_n378), .A3(new_n662), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n856), .A2(new_n722), .A3(new_n842), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(KEYINPUT59), .A3(new_n378), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  AOI211_X1 g665(.A(KEYINPUT57), .B(new_n431), .C1(new_n850), .C2(new_n817), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(KEYINPUT57), .B2(new_n841), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n868), .A2(new_n581), .A3(new_n662), .A4(new_n820), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n866), .B1(new_n869), .B2(G148gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n863), .B1(new_n865), .B2(new_n870), .ZN(G1345gat));
  NAND3_X1  g670(.A1(new_n843), .A2(new_n393), .A3(new_n642), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n856), .A2(new_n641), .A3(new_n842), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n393), .ZN(G1346gat));
  AND2_X1   g673(.A1(new_n395), .A2(new_n397), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n843), .A2(new_n875), .A3(new_n693), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n856), .A2(new_n608), .A3(new_n842), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n875), .ZN(G1347gat));
  AND4_X1   g677(.A1(new_n503), .A2(new_n818), .A3(new_n465), .A4(new_n819), .ZN(new_n879));
  AOI21_X1  g678(.A(G169gat), .B1(new_n879), .B2(new_n250), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n520), .A2(new_n503), .A3(new_n465), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n823), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n251), .A2(new_n233), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(G1348gat));
  INV_X1    g683(.A(G176gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n879), .A2(new_n885), .A3(new_n662), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n823), .A2(new_n722), .A3(new_n881), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n885), .B2(new_n887), .ZN(G1349gat));
  AOI21_X1  g687(.A(new_n277), .B1(new_n882), .B2(new_n642), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n642), .A2(new_n291), .A3(new_n293), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n879), .B2(new_n890), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g691(.A(new_n278), .B1(new_n882), .B2(new_n693), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT61), .Z(new_n894));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n278), .A3(new_n693), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1351gat));
  NOR2_X1   g695(.A1(new_n580), .A2(new_n667), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n503), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT124), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n868), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G197gat), .B1(new_n900), .B2(new_n251), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n818), .A2(new_n503), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n897), .A2(new_n530), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(KEYINPUT122), .B2(new_n903), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n903), .A2(KEYINPUT122), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n251), .A2(G197gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(KEYINPUT123), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(KEYINPUT123), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n901), .B1(new_n909), .B2(new_n910), .ZN(G1352gat));
  INV_X1    g710(.A(new_n906), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n657), .A3(new_n662), .ZN(new_n913));
  XOR2_X1   g712(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n868), .A2(new_n662), .A3(new_n899), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n657), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n918), .B2(new_n917), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n913), .A2(new_n915), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n916), .A2(new_n920), .A3(new_n921), .ZN(G1353gat));
  NAND3_X1  g721(.A1(new_n912), .A2(new_n637), .A3(new_n642), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n868), .A2(new_n642), .A3(new_n899), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n924), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT63), .B1(new_n924), .B2(G211gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1354gat));
  INV_X1    g726(.A(G218gat), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n900), .A2(new_n928), .A3(new_n608), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n906), .B2(new_n608), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT127), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(KEYINPUT127), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1355gat));
endmodule


