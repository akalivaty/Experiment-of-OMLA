

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U547 ( .A(n534), .Z(n514) );
  NOR2_X2 U548 ( .A1(n540), .A2(n539), .ZN(G160) );
  BUF_X1 U549 ( .A(n532), .Z(n515) );
  NOR2_X1 U550 ( .A1(G2105), .A2(n524), .ZN(n532) );
  XNOR2_X2 U551 ( .A(n525), .B(KEYINPUT65), .ZN(n543) );
  XNOR2_X1 U552 ( .A(n714), .B(KEYINPUT95), .ZN(n715) );
  XNOR2_X1 U553 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U554 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n720) );
  XNOR2_X1 U555 ( .A(n721), .B(n720), .ZN(n722) );
  INV_X1 U556 ( .A(KEYINPUT32), .ZN(n735) );
  NOR2_X1 U557 ( .A1(G651), .A2(n634), .ZN(n649) );
  INV_X1 U558 ( .A(G2104), .ZN(n516) );
  NAND2_X1 U559 ( .A1(n516), .A2(KEYINPUT64), .ZN(n519) );
  INV_X1 U560 ( .A(KEYINPUT64), .ZN(n517) );
  NAND2_X1 U561 ( .A1(n517), .A2(G2104), .ZN(n518) );
  NAND2_X1 U562 ( .A1(n519), .A2(n518), .ZN(n524) );
  NAND2_X1 U563 ( .A1(n515), .A2(G102), .ZN(n523) );
  NOR2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XOR2_X1 U565 ( .A(KEYINPUT66), .B(n520), .Z(n521) );
  XNOR2_X1 U566 ( .A(n521), .B(KEYINPUT17), .ZN(n534) );
  NAND2_X1 U567 ( .A1(G138), .A2(n514), .ZN(n522) );
  NAND2_X1 U568 ( .A1(n523), .A2(n522), .ZN(n531) );
  NAND2_X1 U569 ( .A1(n524), .A2(G2105), .ZN(n525) );
  NAND2_X1 U570 ( .A1(G126), .A2(n543), .ZN(n528) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U572 ( .A1(n888), .A2(G114), .ZN(n526) );
  XNOR2_X1 U573 ( .A(n526), .B(KEYINPUT82), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U575 ( .A(KEYINPUT83), .B(n529), .Z(n530) );
  NOR2_X1 U576 ( .A1(n531), .A2(n530), .ZN(G164) );
  NAND2_X1 U577 ( .A1(G101), .A2(n532), .ZN(n533) );
  XOR2_X1 U578 ( .A(n533), .B(KEYINPUT23), .Z(n536) );
  NAND2_X1 U579 ( .A1(G137), .A2(n534), .ZN(n535) );
  NAND2_X1 U580 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U581 ( .A1(G113), .A2(n888), .ZN(n538) );
  NAND2_X1 U582 ( .A1(G125), .A2(n543), .ZN(n537) );
  NAND2_X1 U583 ( .A1(n538), .A2(n537), .ZN(n539) );
  AND2_X1 U584 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U585 ( .A1(G111), .A2(n888), .ZN(n542) );
  NAND2_X1 U586 ( .A1(G135), .A2(n514), .ZN(n541) );
  NAND2_X1 U587 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U588 ( .A1(n543), .A2(G123), .ZN(n544) );
  XOR2_X1 U589 ( .A(KEYINPUT18), .B(n544), .Z(n545) );
  NOR2_X1 U590 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X1 U591 ( .A1(n515), .A2(G99), .ZN(n547) );
  NAND2_X1 U592 ( .A1(n548), .A2(n547), .ZN(n948) );
  XNOR2_X1 U593 ( .A(G2096), .B(n948), .ZN(n549) );
  OR2_X1 U594 ( .A1(G2100), .A2(n549), .ZN(G156) );
  INV_X1 U595 ( .A(G57), .ZN(G237) );
  INV_X1 U596 ( .A(G132), .ZN(G219) );
  INV_X1 U597 ( .A(G82), .ZN(G220) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n641) );
  NAND2_X1 U599 ( .A1(n641), .A2(G89), .ZN(n550) );
  XNOR2_X1 U600 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  XOR2_X1 U601 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  INV_X1 U602 ( .A(G651), .ZN(n555) );
  NOR2_X1 U603 ( .A1(n634), .A2(n555), .ZN(n645) );
  NAND2_X1 U604 ( .A1(G76), .A2(n645), .ZN(n551) );
  NAND2_X1 U605 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U606 ( .A(n553), .B(KEYINPUT5), .ZN(n561) );
  NAND2_X1 U607 ( .A1(n649), .A2(G51), .ZN(n554) );
  XNOR2_X1 U608 ( .A(n554), .B(KEYINPUT74), .ZN(n558) );
  NOR2_X1 U609 ( .A1(G543), .A2(n555), .ZN(n556) );
  XOR2_X1 U610 ( .A(KEYINPUT1), .B(n556), .Z(n642) );
  NAND2_X1 U611 ( .A1(G63), .A2(n642), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U613 ( .A(KEYINPUT6), .B(n559), .Z(n560) );
  NAND2_X1 U614 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U615 ( .A(n562), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .ZN(n563) );
  XNOR2_X1 U617 ( .A(n563), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U618 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U619 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U620 ( .A(G223), .ZN(n828) );
  NAND2_X1 U621 ( .A1(n828), .A2(G567), .ZN(n565) );
  XNOR2_X1 U622 ( .A(n565), .B(KEYINPUT11), .ZN(n566) );
  XNOR2_X1 U623 ( .A(KEYINPUT71), .B(n566), .ZN(G234) );
  NAND2_X1 U624 ( .A1(n641), .A2(G81), .ZN(n567) );
  XNOR2_X1 U625 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G68), .A2(n645), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n571) );
  XOR2_X1 U628 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n570) );
  XNOR2_X1 U629 ( .A(n571), .B(n570), .ZN(n574) );
  NAND2_X1 U630 ( .A1(n642), .A2(G56), .ZN(n572) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n572), .Z(n573) );
  NOR2_X1 U632 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n649), .A2(G43), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n934) );
  INV_X1 U635 ( .A(G860), .ZN(n602) );
  OR2_X1 U636 ( .A1(n934), .A2(n602), .ZN(G153) );
  NAND2_X1 U637 ( .A1(G90), .A2(n641), .ZN(n578) );
  NAND2_X1 U638 ( .A1(G77), .A2(n645), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U640 ( .A(KEYINPUT9), .B(n579), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G64), .A2(n642), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G52), .A2(n649), .ZN(n580) );
  AND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n583), .A2(n582), .ZN(G301) );
  NAND2_X1 U645 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U646 ( .A1(n649), .A2(G54), .ZN(n590) );
  NAND2_X1 U647 ( .A1(G92), .A2(n641), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G66), .A2(n642), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U650 ( .A1(G79), .A2(n645), .ZN(n586) );
  XNOR2_X1 U651 ( .A(KEYINPUT73), .B(n586), .ZN(n587) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U653 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U654 ( .A(KEYINPUT15), .B(n591), .Z(n936) );
  INV_X1 U655 ( .A(G868), .ZN(n659) );
  NAND2_X1 U656 ( .A1(n936), .A2(n659), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G65), .A2(n642), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G53), .A2(n649), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G91), .A2(n641), .ZN(n597) );
  NAND2_X1 U662 ( .A1(G78), .A2(n645), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U664 ( .A1(n599), .A2(n598), .ZN(n925) );
  XOR2_X1 U665 ( .A(n925), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U666 ( .A1(G299), .A2(G868), .ZN(n601) );
  NOR2_X1 U667 ( .A1(G286), .A2(n659), .ZN(n600) );
  NOR2_X1 U668 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n602), .A2(G559), .ZN(n603) );
  INV_X1 U670 ( .A(n936), .ZN(n609) );
  NAND2_X1 U671 ( .A1(n603), .A2(n609), .ZN(n604) );
  XNOR2_X1 U672 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U673 ( .A1(n609), .A2(G868), .ZN(n605) );
  NOR2_X1 U674 ( .A1(G559), .A2(n605), .ZN(n606) );
  XNOR2_X1 U675 ( .A(n606), .B(KEYINPUT76), .ZN(n608) );
  NOR2_X1 U676 ( .A1(n934), .A2(G868), .ZN(n607) );
  NOR2_X1 U677 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U678 ( .A1(G559), .A2(n609), .ZN(n610) );
  XOR2_X1 U679 ( .A(KEYINPUT77), .B(n610), .Z(n611) );
  XNOR2_X1 U680 ( .A(n934), .B(n611), .ZN(n657) );
  NOR2_X1 U681 ( .A1(n657), .A2(G860), .ZN(n618) );
  NAND2_X1 U682 ( .A1(G67), .A2(n642), .ZN(n613) );
  NAND2_X1 U683 ( .A1(G55), .A2(n649), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U685 ( .A1(G93), .A2(n641), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G80), .A2(n645), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n616) );
  OR2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n660) );
  XOR2_X1 U689 ( .A(n618), .B(n660), .Z(G145) );
  NAND2_X1 U690 ( .A1(G85), .A2(n641), .ZN(n620) );
  NAND2_X1 U691 ( .A1(G72), .A2(n645), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n621), .B(KEYINPUT67), .ZN(n623) );
  NAND2_X1 U694 ( .A1(G47), .A2(n649), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U696 ( .A1(G60), .A2(n642), .ZN(n624) );
  XOR2_X1 U697 ( .A(KEYINPUT68), .B(n624), .Z(n625) );
  NOR2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U699 ( .A(KEYINPUT69), .B(n627), .ZN(G290) );
  NAND2_X1 U700 ( .A1(G88), .A2(n641), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G75), .A2(n645), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U703 ( .A1(G62), .A2(n642), .ZN(n631) );
  NAND2_X1 U704 ( .A1(G50), .A2(n649), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U706 ( .A1(n633), .A2(n632), .ZN(G166) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U708 ( .A1(G49), .A2(n649), .ZN(n636) );
  NAND2_X1 U709 ( .A1(G87), .A2(n634), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U711 ( .A1(n642), .A2(n637), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n640), .B(KEYINPUT78), .ZN(G288) );
  NAND2_X1 U714 ( .A1(G86), .A2(n641), .ZN(n644) );
  NAND2_X1 U715 ( .A1(G61), .A2(n642), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n645), .A2(G73), .ZN(n646) );
  XOR2_X1 U718 ( .A(KEYINPUT2), .B(n646), .Z(n647) );
  NOR2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U720 ( .A1(n649), .A2(G48), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(G305) );
  XOR2_X1 U722 ( .A(G299), .B(KEYINPUT19), .Z(n653) );
  XNOR2_X1 U723 ( .A(G166), .B(G288), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n653), .B(n652), .ZN(n654) );
  XOR2_X1 U725 ( .A(n660), .B(n654), .Z(n655) );
  XNOR2_X1 U726 ( .A(n655), .B(G305), .ZN(n656) );
  XNOR2_X1 U727 ( .A(G290), .B(n656), .ZN(n898) );
  XNOR2_X1 U728 ( .A(n657), .B(n898), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n658), .A2(G868), .ZN(n662) );
  NAND2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U731 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT20), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(KEYINPUT79), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n665), .A2(G2090), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n666), .B(KEYINPUT21), .ZN(n667) );
  XNOR2_X1 U737 ( .A(n667), .B(KEYINPUT80), .ZN(n668) );
  NAND2_X1 U738 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U740 ( .A1(G220), .A2(G219), .ZN(n669) );
  XNOR2_X1 U741 ( .A(KEYINPUT22), .B(n669), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n670), .A2(G96), .ZN(n671) );
  NOR2_X1 U743 ( .A1(n671), .A2(G218), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n672), .B(KEYINPUT81), .ZN(n834) );
  NAND2_X1 U745 ( .A1(n834), .A2(G2106), .ZN(n676) );
  NAND2_X1 U746 ( .A1(G108), .A2(G120), .ZN(n673) );
  NOR2_X1 U747 ( .A1(G237), .A2(n673), .ZN(n674) );
  NAND2_X1 U748 ( .A1(G69), .A2(n674), .ZN(n835) );
  NAND2_X1 U749 ( .A1(n835), .A2(G567), .ZN(n675) );
  NAND2_X1 U750 ( .A1(n676), .A2(n675), .ZN(n856) );
  NAND2_X1 U751 ( .A1(G661), .A2(G483), .ZN(n677) );
  NOR2_X1 U752 ( .A1(n856), .A2(n677), .ZN(n831) );
  NAND2_X1 U753 ( .A1(n831), .A2(G36), .ZN(G176) );
  INV_X1 U754 ( .A(G166), .ZN(G303) );
  NOR2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U756 ( .A1(G1971), .A2(G303), .ZN(n678) );
  NOR2_X1 U757 ( .A1(n749), .A2(n678), .ZN(n939) );
  NOR2_X1 U758 ( .A1(G164), .A2(G1384), .ZN(n753) );
  NAND2_X1 U759 ( .A1(G160), .A2(G40), .ZN(n752) );
  XOR2_X1 U760 ( .A(n752), .B(KEYINPUT88), .Z(n680) );
  NAND2_X1 U761 ( .A1(n753), .A2(n680), .ZN(n709) );
  INV_X1 U762 ( .A(n709), .ZN(n703) );
  NAND2_X1 U763 ( .A1(n703), .A2(G2072), .ZN(n681) );
  XNOR2_X1 U764 ( .A(n681), .B(KEYINPUT27), .ZN(n683) );
  XOR2_X1 U765 ( .A(G1956), .B(KEYINPUT92), .Z(n996) );
  NOR2_X1 U766 ( .A1(n703), .A2(n996), .ZN(n682) );
  NOR2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n685) );
  NOR2_X1 U768 ( .A1(n925), .A2(n685), .ZN(n684) );
  XOR2_X1 U769 ( .A(n684), .B(KEYINPUT28), .Z(n700) );
  NAND2_X1 U770 ( .A1(n925), .A2(n685), .ZN(n698) );
  INV_X1 U771 ( .A(G1996), .ZN(n971) );
  NOR2_X1 U772 ( .A1(n709), .A2(n971), .ZN(n686) );
  XOR2_X1 U773 ( .A(n686), .B(KEYINPUT26), .Z(n688) );
  NAND2_X1 U774 ( .A1(n709), .A2(G1341), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U776 ( .A1(n934), .A2(n689), .ZN(n693) );
  NAND2_X1 U777 ( .A1(G1348), .A2(n709), .ZN(n691) );
  NAND2_X1 U778 ( .A1(G2067), .A2(n703), .ZN(n690) );
  NAND2_X1 U779 ( .A1(n691), .A2(n690), .ZN(n694) );
  NOR2_X1 U780 ( .A1(n936), .A2(n694), .ZN(n692) );
  OR2_X1 U781 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U782 ( .A1(n936), .A2(n694), .ZN(n695) );
  NAND2_X1 U783 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U785 ( .A1(n700), .A2(n699), .ZN(n702) );
  XOR2_X1 U786 ( .A(KEYINPUT93), .B(KEYINPUT29), .Z(n701) );
  XNOR2_X1 U787 ( .A(n702), .B(n701), .ZN(n707) );
  NAND2_X1 U788 ( .A1(G1961), .A2(n709), .ZN(n705) );
  XOR2_X1 U789 ( .A(KEYINPUT25), .B(G2078), .Z(n975) );
  NAND2_X1 U790 ( .A1(n703), .A2(n975), .ZN(n704) );
  NAND2_X1 U791 ( .A1(n705), .A2(n704), .ZN(n708) );
  NOR2_X1 U792 ( .A1(n708), .A2(G301), .ZN(n706) );
  NOR2_X1 U793 ( .A1(n707), .A2(n706), .ZN(n723) );
  AND2_X1 U794 ( .A1(G301), .A2(n708), .ZN(n719) );
  INV_X1 U795 ( .A(KEYINPUT91), .ZN(n711) );
  NAND2_X1 U796 ( .A1(G8), .A2(n709), .ZN(n813) );
  NOR2_X1 U797 ( .A1(G1966), .A2(n813), .ZN(n710) );
  XNOR2_X1 U798 ( .A(n711), .B(n710), .ZN(n742) );
  NOR2_X1 U799 ( .A1(G2084), .A2(n709), .ZN(n738) );
  NOR2_X1 U800 ( .A1(n742), .A2(n738), .ZN(n712) );
  XNOR2_X1 U801 ( .A(KEYINPUT94), .B(n712), .ZN(n713) );
  NAND2_X1 U802 ( .A1(n713), .A2(G8), .ZN(n716) );
  INV_X1 U803 ( .A(KEYINPUT30), .ZN(n714) );
  NOR2_X1 U804 ( .A1(G168), .A2(n717), .ZN(n718) );
  NOR2_X1 U805 ( .A1(n719), .A2(n718), .ZN(n721) );
  NOR2_X1 U806 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U807 ( .A(KEYINPUT97), .B(n724), .ZN(n737) );
  AND2_X1 U808 ( .A1(G286), .A2(G8), .ZN(n725) );
  NAND2_X1 U809 ( .A1(n737), .A2(n725), .ZN(n734) );
  INV_X1 U810 ( .A(G8), .ZN(n732) );
  NOR2_X1 U811 ( .A1(G1971), .A2(n813), .ZN(n726) );
  XOR2_X1 U812 ( .A(KEYINPUT98), .B(n726), .Z(n727) );
  NAND2_X1 U813 ( .A1(n727), .A2(G303), .ZN(n729) );
  NOR2_X1 U814 ( .A1(G2090), .A2(n709), .ZN(n728) );
  NOR2_X1 U815 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U816 ( .A(n730), .B(KEYINPUT99), .ZN(n731) );
  OR2_X1 U817 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U818 ( .A1(n734), .A2(n733), .ZN(n736) );
  XNOR2_X1 U819 ( .A(n736), .B(n735), .ZN(n746) );
  INV_X1 U820 ( .A(n737), .ZN(n741) );
  NAND2_X1 U821 ( .A1(G8), .A2(n738), .ZN(n739) );
  XOR2_X1 U822 ( .A(KEYINPUT90), .B(n739), .Z(n740) );
  NOR2_X1 U823 ( .A1(n741), .A2(n740), .ZN(n744) );
  INV_X1 U824 ( .A(n742), .ZN(n743) );
  NAND2_X1 U825 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U826 ( .A1(n746), .A2(n745), .ZN(n807) );
  NAND2_X1 U827 ( .A1(n939), .A2(n807), .ZN(n747) );
  NAND2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n928) );
  NAND2_X1 U829 ( .A1(n747), .A2(n928), .ZN(n748) );
  XNOR2_X1 U830 ( .A(KEYINPUT100), .B(n748), .ZN(n789) );
  NAND2_X1 U831 ( .A1(n749), .A2(KEYINPUT33), .ZN(n750) );
  OR2_X1 U832 ( .A1(n750), .A2(n813), .ZN(n751) );
  XOR2_X1 U833 ( .A(G1981), .B(G305), .Z(n920) );
  NAND2_X1 U834 ( .A1(n751), .A2(n920), .ZN(n784) );
  NOR2_X1 U835 ( .A1(n753), .A2(n752), .ZN(n801) );
  NAND2_X1 U836 ( .A1(G116), .A2(n888), .ZN(n755) );
  NAND2_X1 U837 ( .A1(G128), .A2(n543), .ZN(n754) );
  NAND2_X1 U838 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U839 ( .A(n756), .B(KEYINPUT35), .ZN(n761) );
  NAND2_X1 U840 ( .A1(n515), .A2(G104), .ZN(n758) );
  NAND2_X1 U841 ( .A1(G140), .A2(n514), .ZN(n757) );
  NAND2_X1 U842 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U843 ( .A(KEYINPUT34), .B(n759), .Z(n760) );
  NAND2_X1 U844 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U845 ( .A(n762), .B(KEYINPUT36), .Z(n894) );
  XNOR2_X1 U846 ( .A(G2067), .B(KEYINPUT37), .ZN(n790) );
  NOR2_X1 U847 ( .A1(n894), .A2(n790), .ZN(n960) );
  NAND2_X1 U848 ( .A1(n801), .A2(n960), .ZN(n797) );
  XNOR2_X1 U849 ( .A(n801), .B(KEYINPUT86), .ZN(n780) );
  NAND2_X1 U850 ( .A1(n543), .A2(G119), .ZN(n763) );
  XOR2_X1 U851 ( .A(KEYINPUT84), .B(n763), .Z(n768) );
  NAND2_X1 U852 ( .A1(n515), .A2(G95), .ZN(n765) );
  NAND2_X1 U853 ( .A1(G131), .A2(n514), .ZN(n764) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U855 ( .A(KEYINPUT85), .B(n766), .Z(n767) );
  NOR2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n888), .A2(G107), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n882) );
  NAND2_X1 U859 ( .A1(G1991), .A2(n882), .ZN(n779) );
  NAND2_X1 U860 ( .A1(G117), .A2(n888), .ZN(n772) );
  NAND2_X1 U861 ( .A1(G141), .A2(n514), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n515), .A2(G105), .ZN(n773) );
  XOR2_X1 U864 ( .A(KEYINPUT38), .B(n773), .Z(n774) );
  NOR2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n543), .A2(G129), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n867) );
  NAND2_X1 U868 ( .A1(G1996), .A2(n867), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n959) );
  NAND2_X1 U870 ( .A1(n780), .A2(n959), .ZN(n781) );
  XNOR2_X1 U871 ( .A(n781), .B(KEYINPUT87), .ZN(n794) );
  INV_X1 U872 ( .A(n794), .ZN(n782) );
  AND2_X1 U873 ( .A1(n797), .A2(n782), .ZN(n816) );
  INV_X1 U874 ( .A(n816), .ZN(n783) );
  OR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n786) );
  XNOR2_X1 U876 ( .A(G1986), .B(G290), .ZN(n931) );
  NAND2_X1 U877 ( .A1(n931), .A2(n801), .ZN(n818) );
  INV_X1 U878 ( .A(n818), .ZN(n785) );
  NOR2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n821) );
  INV_X1 U880 ( .A(n821), .ZN(n787) );
  OR2_X1 U881 ( .A1(n813), .A2(n787), .ZN(n788) );
  NOR2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n804) );
  AND2_X1 U883 ( .A1(n894), .A2(n790), .ZN(n791) );
  XOR2_X1 U884 ( .A(KEYINPUT102), .B(n791), .Z(n965) );
  NOR2_X1 U885 ( .A1(G1996), .A2(n867), .ZN(n946) );
  NOR2_X1 U886 ( .A1(G1986), .A2(G290), .ZN(n792) );
  NOR2_X1 U887 ( .A1(G1991), .A2(n882), .ZN(n950) );
  NOR2_X1 U888 ( .A1(n792), .A2(n950), .ZN(n793) );
  NOR2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U890 ( .A1(n946), .A2(n795), .ZN(n796) );
  XNOR2_X1 U891 ( .A(n796), .B(KEYINPUT39), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U893 ( .A(KEYINPUT101), .B(n799), .Z(n800) );
  NAND2_X1 U894 ( .A1(n965), .A2(n800), .ZN(n802) );
  AND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n825) );
  NOR2_X1 U897 ( .A1(G2090), .A2(G303), .ZN(n805) );
  NAND2_X1 U898 ( .A1(G8), .A2(n805), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n810) );
  AND2_X1 U900 ( .A1(n813), .A2(n816), .ZN(n808) );
  AND2_X1 U901 ( .A1(n808), .A2(n818), .ZN(n809) );
  AND2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n820) );
  NOR2_X1 U903 ( .A1(G1981), .A2(G305), .ZN(n811) );
  XNOR2_X1 U904 ( .A(n811), .B(KEYINPUT24), .ZN(n812) );
  XNOR2_X1 U905 ( .A(n812), .B(KEYINPUT89), .ZN(n814) );
  NOR2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n817) );
  AND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U909 ( .A1(n820), .A2(n819), .ZN(n823) );
  NAND2_X1 U910 ( .A1(n821), .A2(KEYINPUT33), .ZN(n822) );
  AND2_X1 U911 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U912 ( .A1(n825), .A2(n824), .ZN(n827) );
  XOR2_X1 U913 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n826) );
  XNOR2_X1 U914 ( .A(n827), .B(n826), .ZN(G329) );
  INV_X1 U915 ( .A(G301), .ZN(G171) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n828), .ZN(G217) );
  NAND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n829) );
  XNOR2_X1 U918 ( .A(KEYINPUT105), .B(n829), .ZN(n830) );
  NAND2_X1 U919 ( .A1(n830), .A2(G661), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G1), .A2(G3), .ZN(n832) );
  NAND2_X1 U921 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U922 ( .A(n833), .B(KEYINPUT106), .ZN(G188) );
  XNOR2_X1 U923 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  INV_X1 U925 ( .A(G108), .ZN(G238) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  NOR2_X1 U927 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  XOR2_X1 U929 ( .A(G2474), .B(G1986), .Z(n837) );
  XNOR2_X1 U930 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U932 ( .A(n838), .B(KEYINPUT109), .Z(n840) );
  XNOR2_X1 U933 ( .A(G1966), .B(G1981), .ZN(n839) );
  XNOR2_X1 U934 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U935 ( .A(G1976), .B(G1971), .Z(n842) );
  XNOR2_X1 U936 ( .A(G1961), .B(G1956), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U938 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U939 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n845) );
  XNOR2_X1 U940 ( .A(n846), .B(n845), .ZN(G229) );
  XOR2_X1 U941 ( .A(G2096), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U942 ( .A(G2090), .B(KEYINPUT42), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U944 ( .A(n849), .B(G2678), .Z(n851) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U946 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U947 ( .A(KEYINPUT108), .B(G2100), .Z(n853) );
  XNOR2_X1 U948 ( .A(G2084), .B(G2078), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U950 ( .A(n855), .B(n854), .ZN(G227) );
  INV_X1 U951 ( .A(n856), .ZN(G319) );
  NAND2_X1 U952 ( .A1(n514), .A2(G136), .ZN(n857) );
  XNOR2_X1 U953 ( .A(n857), .B(KEYINPUT112), .ZN(n860) );
  NAND2_X1 U954 ( .A1(G100), .A2(n515), .ZN(n858) );
  XOR2_X1 U955 ( .A(KEYINPUT113), .B(n858), .Z(n859) );
  NAND2_X1 U956 ( .A1(n860), .A2(n859), .ZN(n866) );
  NAND2_X1 U957 ( .A1(G124), .A2(n543), .ZN(n861) );
  XOR2_X1 U958 ( .A(KEYINPUT44), .B(n861), .Z(n862) );
  XNOR2_X1 U959 ( .A(n862), .B(KEYINPUT111), .ZN(n864) );
  NAND2_X1 U960 ( .A1(G112), .A2(n888), .ZN(n863) );
  NAND2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U962 ( .A1(n866), .A2(n865), .ZN(G162) );
  XNOR2_X1 U963 ( .A(G164), .B(n867), .ZN(n868) );
  XNOR2_X1 U964 ( .A(n868), .B(n948), .ZN(n881) );
  XOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n879) );
  NAND2_X1 U966 ( .A1(G118), .A2(n888), .ZN(n870) );
  NAND2_X1 U967 ( .A1(G130), .A2(n543), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U969 ( .A1(n515), .A2(G106), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G142), .A2(n514), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(KEYINPUT45), .B(n873), .Z(n874) );
  XNOR2_X1 U973 ( .A(KEYINPUT114), .B(n874), .ZN(n875) );
  NOR2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U975 ( .A(G160), .B(n877), .ZN(n878) );
  XNOR2_X1 U976 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n881), .B(n880), .ZN(n884) );
  XNOR2_X1 U978 ( .A(n882), .B(G162), .ZN(n883) );
  XNOR2_X1 U979 ( .A(n884), .B(n883), .ZN(n896) );
  NAND2_X1 U980 ( .A1(n515), .A2(G103), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G139), .A2(n514), .ZN(n885) );
  NAND2_X1 U982 ( .A1(n886), .A2(n885), .ZN(n893) );
  NAND2_X1 U983 ( .A1(n543), .A2(G127), .ZN(n887) );
  XOR2_X1 U984 ( .A(KEYINPUT115), .B(n887), .Z(n890) );
  NAND2_X1 U985 ( .A1(n888), .A2(G115), .ZN(n889) );
  NAND2_X1 U986 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U987 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n955) );
  XNOR2_X1 U989 ( .A(n955), .B(n894), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U991 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U992 ( .A(G286), .B(n936), .ZN(n899) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n934), .B(G171), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G397) );
  NOR2_X1 U997 ( .A1(G229), .A2(G227), .ZN(n904) );
  XNOR2_X1 U998 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n916) );
  XOR2_X1 U1000 ( .A(G2443), .B(G2427), .Z(n906) );
  XNOR2_X1 U1001 ( .A(G2438), .B(G2454), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1003 ( .A(n907), .B(G2435), .Z(n909) );
  XNOR2_X1 U1004 ( .A(G1341), .B(G1348), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n913) );
  XOR2_X1 U1006 ( .A(G2430), .B(G2446), .Z(n911) );
  XNOR2_X1 U1007 ( .A(KEYINPUT104), .B(G2451), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1009 ( .A(n913), .B(n912), .Z(n914) );
  NAND2_X1 U1010 ( .A1(G14), .A2(n914), .ZN(n919) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n919), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G69), .ZN(G235) );
  INV_X1 U1017 ( .A(n919), .ZN(G401) );
  XOR2_X1 U1018 ( .A(KEYINPUT56), .B(G16), .Z(n944) );
  XNOR2_X1 U1019 ( .A(G1966), .B(G168), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n922), .B(KEYINPUT57), .ZN(n933) );
  XNOR2_X1 U1022 ( .A(G171), .B(G1961), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(G1971), .A2(G303), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1025 ( .A(n925), .B(G1956), .Z(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n942) );
  XNOR2_X1 U1030 ( .A(G1341), .B(KEYINPUT124), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(n935), .B(n934), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(G1348), .B(n936), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n1024) );
  XOR2_X1 U1037 ( .A(G2090), .B(G162), .Z(n945) );
  NOR2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1039 ( .A(KEYINPUT51), .B(n947), .Z(n954) );
  XNOR2_X1 U1040 ( .A(G160), .B(G2084), .ZN(n949) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n951) );
  NOR2_X1 U1042 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1043 ( .A(KEYINPUT117), .B(n952), .Z(n953) );
  NAND2_X1 U1044 ( .A1(n954), .A2(n953), .ZN(n964) );
  XOR2_X1 U1045 ( .A(G2072), .B(n955), .Z(n957) );
  XOR2_X1 U1046 ( .A(G164), .B(G2078), .Z(n956) );
  NOR2_X1 U1047 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1048 ( .A(KEYINPUT50), .B(n958), .ZN(n962) );
  NOR2_X1 U1049 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1050 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1051 ( .A1(n964), .A2(n963), .ZN(n966) );
  NAND2_X1 U1052 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1053 ( .A(n967), .B(KEYINPUT118), .ZN(n968) );
  XNOR2_X1 U1054 ( .A(KEYINPUT52), .B(n968), .ZN(n969) );
  NAND2_X1 U1055 ( .A1(n969), .A2(G29), .ZN(n1022) );
  XOR2_X1 U1056 ( .A(G1991), .B(G25), .Z(n970) );
  NAND2_X1 U1057 ( .A1(G28), .A2(n970), .ZN(n974) );
  XOR2_X1 U1058 ( .A(G32), .B(n971), .Z(n972) );
  XNOR2_X1 U1059 ( .A(KEYINPUT122), .B(n972), .ZN(n973) );
  NOR2_X1 U1060 ( .A1(n974), .A2(n973), .ZN(n983) );
  XNOR2_X1 U1061 ( .A(n975), .B(G27), .ZN(n981) );
  XNOR2_X1 U1062 ( .A(G2067), .B(KEYINPUT120), .ZN(n976) );
  XNOR2_X1 U1063 ( .A(n976), .B(G26), .ZN(n978) );
  XNOR2_X1 U1064 ( .A(G33), .B(G2072), .ZN(n977) );
  NOR2_X1 U1065 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1066 ( .A(KEYINPUT121), .B(n979), .ZN(n980) );
  NOR2_X1 U1067 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1068 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1069 ( .A(n984), .B(KEYINPUT53), .ZN(n987) );
  XOR2_X1 U1070 ( .A(G2084), .B(G34), .Z(n985) );
  XNOR2_X1 U1071 ( .A(KEYINPUT54), .B(n985), .ZN(n986) );
  NAND2_X1 U1072 ( .A1(n987), .A2(n986), .ZN(n990) );
  XOR2_X1 U1073 ( .A(KEYINPUT119), .B(G2090), .Z(n988) );
  XNOR2_X1 U1074 ( .A(G35), .B(n988), .ZN(n989) );
  NOR2_X1 U1075 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1076 ( .A(KEYINPUT123), .B(n991), .Z(n992) );
  NOR2_X1 U1077 ( .A1(G29), .A2(n992), .ZN(n993) );
  XOR2_X1 U1078 ( .A(KEYINPUT55), .B(n993), .Z(n1020) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G21), .ZN(n995) );
  XNOR2_X1 U1080 ( .A(G1961), .B(G5), .ZN(n994) );
  NOR2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n1007) );
  XOR2_X1 U1082 ( .A(G1341), .B(G19), .Z(n998) );
  XNOR2_X1 U1083 ( .A(n996), .B(G20), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1004) );
  XOR2_X1 U1085 ( .A(G1981), .B(G6), .Z(n1002) );
  XOR2_X1 U1086 ( .A(G1348), .B(G4), .Z(n999) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(n999), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(KEYINPUT59), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1005), .B(KEYINPUT60), .ZN(n1006) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1014) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G23), .B(G1976), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XOR2_X1 U1096 ( .A(G1986), .B(G24), .Z(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(KEYINPUT61), .B(n1015), .Z(n1016) );
  NOR2_X1 U1101 ( .A1(G16), .A2(n1016), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(KEYINPUT126), .B(n1017), .Z(n1018) );
  NAND2_X1 U1103 ( .A1(G11), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1106 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1025), .Z(n1026) );
  XNOR2_X1 U1108 ( .A(KEYINPUT127), .B(n1026), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

