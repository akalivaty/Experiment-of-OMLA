

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591;

  XNOR2_X1 U322 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U323 ( .A(n332), .B(n331), .ZN(n338) );
  XNOR2_X1 U324 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n393) );
  XNOR2_X1 U325 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U326 ( .A(n394), .B(n393), .ZN(n533) );
  XNOR2_X1 U327 ( .A(n345), .B(n344), .ZN(n562) );
  XOR2_X1 U328 ( .A(n365), .B(n364), .Z(n585) );
  XNOR2_X1 U329 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U330 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT71), .B(G92GAT), .Z(n291) );
  XNOR2_X1 U332 ( .A(G99GAT), .B(G85GAT), .ZN(n290) );
  XNOR2_X1 U333 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U334 ( .A(G106GAT), .B(n292), .Z(n343) );
  XOR2_X1 U335 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n295) );
  XOR2_X1 U336 ( .A(G176GAT), .B(G71GAT), .Z(n310) );
  XNOR2_X1 U337 ( .A(G120GAT), .B(G148GAT), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n293), .B(G57GAT), .ZN(n427) );
  XNOR2_X1 U339 ( .A(n310), .B(n427), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n343), .B(n296), .ZN(n305) );
  XOR2_X1 U342 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n298) );
  NAND2_X1 U343 ( .A1(G230GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U345 ( .A(n299), .B(KEYINPUT33), .Z(n303) );
  XNOR2_X1 U346 ( .A(G78GAT), .B(KEYINPUT70), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n300), .B(G204GAT), .ZN(n446) );
  XNOR2_X1 U348 ( .A(G64GAT), .B(KEYINPUT13), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n301), .B(KEYINPUT69), .ZN(n357) );
  XNOR2_X1 U350 ( .A(n446), .B(n357), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n582) );
  XNOR2_X1 U353 ( .A(n582), .B(KEYINPUT41), .ZN(n556) );
  XOR2_X1 U354 ( .A(KEYINPUT111), .B(n556), .Z(n539) );
  INV_X1 U355 ( .A(KEYINPUT122), .ZN(n457) );
  XOR2_X1 U356 ( .A(G120GAT), .B(KEYINPUT82), .Z(n307) );
  XNOR2_X1 U357 ( .A(G15GAT), .B(G99GAT), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n318) );
  XOR2_X1 U359 ( .A(G127GAT), .B(KEYINPUT80), .Z(n309) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n421) );
  XOR2_X1 U362 ( .A(n310), .B(n421), .Z(n312) );
  NAND2_X1 U363 ( .A1(G227GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U365 ( .A(n313), .B(KEYINPUT20), .Z(n316) );
  XNOR2_X1 U366 ( .A(G43GAT), .B(G190GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n314), .B(G134GAT), .ZN(n325) );
  XNOR2_X1 U368 ( .A(n325), .B(KEYINPUT83), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n323) );
  XNOR2_X1 U371 ( .A(KEYINPUT17), .B(KEYINPUT81), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n319), .B(KEYINPUT19), .ZN(n320) );
  XOR2_X1 U373 ( .A(n320), .B(KEYINPUT18), .Z(n322) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(G183GAT), .ZN(n321) );
  XOR2_X1 U375 ( .A(n322), .B(n321), .Z(n410) );
  XNOR2_X1 U376 ( .A(n323), .B(n410), .ZN(n535) );
  INV_X1 U377 ( .A(KEYINPUT75), .ZN(n346) );
  INV_X1 U378 ( .A(n325), .ZN(n324) );
  XOR2_X1 U379 ( .A(G36GAT), .B(G218GAT), .Z(n395) );
  NAND2_X1 U380 ( .A1(n324), .A2(n395), .ZN(n328) );
  INV_X1 U381 ( .A(n395), .ZN(n326) );
  NAND2_X1 U382 ( .A1(n326), .A2(n325), .ZN(n327) );
  NAND2_X1 U383 ( .A1(n328), .A2(n327), .ZN(n332) );
  NAND2_X1 U384 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  INV_X1 U385 ( .A(KEYINPUT11), .ZN(n329) );
  INV_X1 U386 ( .A(n338), .ZN(n336) );
  XOR2_X1 U387 ( .A(G29GAT), .B(KEYINPUT7), .Z(n334) );
  XNOR2_X1 U388 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n370) );
  XNOR2_X1 U390 ( .A(n370), .B(KEYINPUT74), .ZN(n337) );
  INV_X1 U391 ( .A(n337), .ZN(n335) );
  NAND2_X1 U392 ( .A1(n336), .A2(n335), .ZN(n340) );
  NAND2_X1 U393 ( .A1(n338), .A2(n337), .ZN(n339) );
  NAND2_X1 U394 ( .A1(n340), .A2(n339), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n341), .B(KEYINPUT9), .ZN(n345) );
  XOR2_X1 U396 ( .A(G50GAT), .B(G162GAT), .Z(n442) );
  XOR2_X1 U397 ( .A(n442), .B(KEYINPUT10), .Z(n342) );
  XNOR2_X1 U398 ( .A(n346), .B(n562), .ZN(n462) );
  XNOR2_X1 U399 ( .A(n462), .B(KEYINPUT36), .ZN(n493) );
  XOR2_X1 U400 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n348) );
  XNOR2_X1 U401 ( .A(G57GAT), .B(KEYINPUT76), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n365) );
  XOR2_X1 U403 ( .A(G211GAT), .B(G78GAT), .Z(n350) );
  XNOR2_X1 U404 ( .A(G71GAT), .B(G155GAT), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n352) );
  XOR2_X1 U406 ( .A(G183GAT), .B(G127GAT), .Z(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n361) );
  XNOR2_X1 U408 ( .A(KEYINPUT79), .B(KEYINPUT77), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n353), .B(KEYINPUT12), .ZN(n354) );
  XOR2_X1 U410 ( .A(n354), .B(KEYINPUT78), .Z(n359) );
  XOR2_X1 U411 ( .A(G1GAT), .B(G8GAT), .Z(n356) );
  XNOR2_X1 U412 ( .A(G15GAT), .B(G22GAT), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n369) );
  XNOR2_X1 U414 ( .A(n369), .B(n357), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n363) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n364) );
  INV_X1 U419 ( .A(n585), .ZN(n366) );
  NOR2_X1 U420 ( .A1(n493), .A2(n366), .ZN(n368) );
  INV_X1 U421 ( .A(KEYINPUT45), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n385) );
  XNOR2_X1 U423 ( .A(n370), .B(n369), .ZN(n383) );
  XOR2_X1 U424 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n372) );
  NAND2_X1 U425 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U426 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U427 ( .A(n373), .B(KEYINPUT29), .Z(n381) );
  XOR2_X1 U428 ( .A(G113GAT), .B(G50GAT), .Z(n375) );
  XNOR2_X1 U429 ( .A(G36GAT), .B(G43GAT), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U431 ( .A(KEYINPUT67), .B(G197GAT), .Z(n377) );
  XNOR2_X1 U432 ( .A(G169GAT), .B(G141GAT), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U435 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n383), .B(n382), .ZN(n577) );
  INV_X1 U437 ( .A(n577), .ZN(n537) );
  NAND2_X1 U438 ( .A1(n582), .A2(n537), .ZN(n384) );
  NOR2_X1 U439 ( .A1(n385), .A2(n384), .ZN(n392) );
  XOR2_X1 U440 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n387) );
  NAND2_X1 U441 ( .A1(n577), .A2(n556), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n388) );
  NOR2_X1 U443 ( .A1(n585), .A2(n388), .ZN(n389) );
  NAND2_X1 U444 ( .A1(n389), .A2(n562), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n390), .B(KEYINPUT47), .ZN(n391) );
  NOR2_X1 U446 ( .A1(n392), .A2(n391), .ZN(n394) );
  XOR2_X1 U447 ( .A(n395), .B(G92GAT), .Z(n399) );
  XOR2_X1 U448 ( .A(G211GAT), .B(KEYINPUT21), .Z(n397) );
  XNOR2_X1 U449 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n397), .B(n396), .ZN(n441) );
  XNOR2_X1 U451 ( .A(G190GAT), .B(n441), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U453 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n401) );
  NAND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U456 ( .A(n403), .B(n402), .Z(n408) );
  XOR2_X1 U457 ( .A(G64GAT), .B(G204GAT), .Z(n405) );
  XNOR2_X1 U458 ( .A(G8GAT), .B(G176GAT), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n406), .B(KEYINPUT97), .ZN(n407) );
  XNOR2_X1 U461 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U462 ( .A(n410), .B(n409), .ZN(n470) );
  INV_X1 U463 ( .A(n470), .ZN(n524) );
  NOR2_X1 U464 ( .A1(n533), .A2(n524), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n411), .B(KEYINPUT54), .ZN(n433) );
  XOR2_X1 U466 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n413) );
  XNOR2_X1 U467 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U469 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n415) );
  XNOR2_X1 U470 ( .A(KEYINPUT90), .B(KEYINPUT92), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U472 ( .A(n417), .B(n416), .Z(n426) );
  XOR2_X1 U473 ( .A(KEYINPUT88), .B(KEYINPUT3), .Z(n419) );
  XNOR2_X1 U474 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U476 ( .A(G141GAT), .B(n420), .Z(n452) );
  XOR2_X1 U477 ( .A(n421), .B(KEYINPUT1), .Z(n423) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n452), .B(n424), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n432) );
  XOR2_X1 U482 ( .A(n427), .B(G85GAT), .Z(n429) );
  XNOR2_X1 U483 ( .A(G29GAT), .B(G134GAT), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U485 ( .A(G162GAT), .B(n430), .Z(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n476) );
  XNOR2_X1 U487 ( .A(KEYINPUT94), .B(n476), .ZN(n522) );
  NAND2_X1 U488 ( .A1(n433), .A2(n522), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n434), .B(KEYINPUT65), .ZN(n575) );
  XOR2_X1 U490 ( .A(G148GAT), .B(KEYINPUT23), .Z(n436) );
  XNOR2_X1 U491 ( .A(KEYINPUT24), .B(KEYINPUT85), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U493 ( .A(KEYINPUT86), .B(G106GAT), .Z(n438) );
  XNOR2_X1 U494 ( .A(G22GAT), .B(G218GAT), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n450) );
  XOR2_X1 U497 ( .A(n442), .B(n441), .Z(n444) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U500 ( .A(n445), .B(KEYINPUT89), .Z(n448) );
  XNOR2_X1 U501 ( .A(n446), .B(KEYINPUT22), .ZN(n447) );
  XNOR2_X1 U502 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(n472) );
  NAND2_X1 U505 ( .A1(n575), .A2(n472), .ZN(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n455) );
  NAND2_X1 U508 ( .A1(n535), .A2(n455), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n457), .B(n456), .ZN(n569) );
  NAND2_X1 U510 ( .A1(n539), .A2(n569), .ZN(n461) );
  XOR2_X1 U511 ( .A(G176GAT), .B(KEYINPUT123), .Z(n459) );
  XOR2_X1 U512 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n458) );
  NAND2_X1 U513 ( .A1(n577), .A2(n582), .ZN(n498) );
  NAND2_X1 U514 ( .A1(n585), .A2(n462), .ZN(n463) );
  XOR2_X1 U515 ( .A(KEYINPUT16), .B(n463), .Z(n481) );
  XNOR2_X1 U516 ( .A(n535), .B(KEYINPUT84), .ZN(n466) );
  INV_X1 U517 ( .A(n522), .ZN(n553) );
  XNOR2_X1 U518 ( .A(KEYINPUT28), .B(n472), .ZN(n529) );
  AND2_X1 U519 ( .A1(n553), .A2(n529), .ZN(n464) );
  XOR2_X1 U520 ( .A(KEYINPUT27), .B(n524), .Z(n469) );
  NAND2_X1 U521 ( .A1(n464), .A2(n469), .ZN(n534) );
  XNOR2_X1 U522 ( .A(n534), .B(KEYINPUT98), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n467), .B(KEYINPUT99), .ZN(n479) );
  NOR2_X1 U525 ( .A1(n472), .A2(n535), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n468), .B(KEYINPUT26), .ZN(n576) );
  NAND2_X1 U527 ( .A1(n576), .A2(n469), .ZN(n551) );
  XNOR2_X1 U528 ( .A(KEYINPUT100), .B(n551), .ZN(n475) );
  NAND2_X1 U529 ( .A1(n470), .A2(n535), .ZN(n471) );
  NAND2_X1 U530 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U531 ( .A(KEYINPUT25), .B(n473), .Z(n474) );
  NAND2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n477) );
  NAND2_X1 U533 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n480) );
  XOR2_X1 U535 ( .A(KEYINPUT101), .B(n480), .Z(n495) );
  NAND2_X1 U536 ( .A1(n481), .A2(n495), .ZN(n511) );
  OR2_X1 U537 ( .A1(n498), .A2(n511), .ZN(n488) );
  NOR2_X1 U538 ( .A1(n522), .A2(n488), .ZN(n483) );
  XNOR2_X1 U539 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U541 ( .A(G1GAT), .B(n484), .Z(G1324GAT) );
  NOR2_X1 U542 ( .A1(n524), .A2(n488), .ZN(n485) );
  XOR2_X1 U543 ( .A(G8GAT), .B(n485), .Z(G1325GAT) );
  INV_X1 U544 ( .A(n535), .ZN(n526) );
  NOR2_X1 U545 ( .A1(n526), .A2(n488), .ZN(n487) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n529), .A2(n488), .ZN(n490) );
  XNOR2_X1 U549 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G22GAT), .B(n491), .ZN(G1327GAT) );
  XNOR2_X1 U552 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT37), .ZN(n497) );
  NOR2_X1 U554 ( .A1(n493), .A2(n585), .ZN(n494) );
  NAND2_X1 U555 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(n521) );
  NOR2_X1 U557 ( .A1(n521), .A2(n498), .ZN(n500) );
  XNOR2_X1 U558 ( .A(KEYINPUT38), .B(KEYINPUT107), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(n508) );
  NOR2_X1 U560 ( .A1(n508), .A2(n522), .ZN(n503) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(KEYINPUT108), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n508), .A2(n524), .ZN(n505) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(KEYINPUT109), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1329GAT) );
  NOR2_X1 U567 ( .A1(n526), .A2(n508), .ZN(n506) );
  XOR2_X1 U568 ( .A(n506), .B(KEYINPUT40), .Z(n507) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NOR2_X1 U570 ( .A1(n529), .A2(n508), .ZN(n509) );
  XOR2_X1 U571 ( .A(KEYINPUT110), .B(n509), .Z(n510) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(n510), .ZN(G1331GAT) );
  NAND2_X1 U573 ( .A1(n537), .A2(n539), .ZN(n520) );
  OR2_X1 U574 ( .A1(n520), .A2(n511), .ZN(n517) );
  NOR2_X1 U575 ( .A1(n522), .A2(n517), .ZN(n512) );
  XOR2_X1 U576 ( .A(n512), .B(KEYINPUT42), .Z(n513) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U578 ( .A1(n524), .A2(n517), .ZN(n514) );
  XOR2_X1 U579 ( .A(KEYINPUT112), .B(n514), .Z(n515) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NOR2_X1 U581 ( .A1(n526), .A2(n517), .ZN(n516) );
  XOR2_X1 U582 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U583 ( .A1(n529), .A2(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  OR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n528) );
  NOR2_X1 U587 ( .A1(n522), .A2(n528), .ZN(n523) );
  XOR2_X1 U588 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n528), .ZN(n525) );
  XOR2_X1 U590 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U591 ( .A1(n526), .A2(n528), .ZN(n527) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n527), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U594 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n533), .A2(n534), .ZN(n536) );
  NAND2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n548) );
  NOR2_X1 U599 ( .A1(n537), .A2(n548), .ZN(n538) );
  XOR2_X1 U600 ( .A(G113GAT), .B(n538), .Z(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  INV_X1 U602 ( .A(n548), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n545), .A2(n539), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n543) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U608 ( .A(KEYINPUT115), .B(n544), .Z(n547) );
  NAND2_X1 U609 ( .A1(n545), .A2(n585), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(G1342GAT) );
  NOR2_X1 U611 ( .A1(n462), .A2(n548), .ZN(n550) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NOR2_X1 U614 ( .A1(n533), .A2(n551), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U616 ( .A(KEYINPUT118), .B(n554), .Z(n564) );
  NAND2_X1 U617 ( .A1(n564), .A2(n577), .ZN(n555) );
  XNOR2_X1 U618 ( .A(n555), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n558) );
  NAND2_X1 U620 ( .A1(n564), .A2(n556), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n559), .ZN(G1345GAT) );
  XOR2_X1 U623 ( .A(G155GAT), .B(KEYINPUT119), .Z(n561) );
  NAND2_X1 U624 ( .A1(n585), .A2(n564), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(G1346GAT) );
  INV_X1 U626 ( .A(n562), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT120), .ZN(n566) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(n566), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n577), .A2(n569), .ZN(n567) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n567), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n569), .A2(n585), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U634 ( .A(n569), .ZN(n570) );
  NOR2_X1 U635 ( .A1(n570), .A2(n462), .ZN(n574) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT125), .B(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1351GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n576), .ZN(n589) );
  INV_X1 U641 ( .A(n589), .ZN(n586) );
  NAND2_X1 U642 ( .A1(n586), .A2(n577), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT59), .B(KEYINPUT126), .Z(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  OR2_X1 U648 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .Z(n588) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n493), .A2(n589), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

