

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716;

  INV_X1 U369 ( .A(G953), .ZN(n703) );
  INV_X1 U370 ( .A(n635), .ZN(n525) );
  OR2_X2 U371 ( .A1(n594), .A2(G902), .ZN(n441) );
  XOR2_X2 U372 ( .A(KEYINPUT38), .B(n559), .Z(n647) );
  INV_X2 U373 ( .A(n507), .ZN(n559) );
  XNOR2_X1 U374 ( .A(n371), .B(n370), .ZN(n506) );
  XNOR2_X1 U375 ( .A(n361), .B(n360), .ZN(n695) );
  XNOR2_X1 U376 ( .A(n355), .B(G110), .ZN(n425) );
  NAND2_X1 U377 ( .A1(n571), .A2(n354), .ZN(n575) );
  BUF_X1 U378 ( .A(n559), .Z(n349) );
  XNOR2_X1 U379 ( .A(n695), .B(n369), .ZN(n578) );
  XNOR2_X1 U380 ( .A(n356), .B(n351), .ZN(n361) );
  XOR2_X1 U381 ( .A(n425), .B(n384), .Z(n356) );
  XNOR2_X1 U382 ( .A(G143), .B(G128), .ZN(n386) );
  XOR2_X1 U383 ( .A(G146), .B(G125), .Z(n406) );
  AND2_X2 U384 ( .A1(n575), .A2(n574), .ZN(n348) );
  AND2_X1 U385 ( .A1(n575), .A2(n574), .ZN(n682) );
  NOR2_X1 U386 ( .A1(n489), .A2(n486), .ZN(n410) );
  XNOR2_X1 U387 ( .A(n488), .B(KEYINPUT101), .ZN(n539) );
  XNOR2_X1 U388 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U389 ( .A(n466), .B(n465), .ZN(n658) );
  AND2_X1 U390 ( .A1(n638), .A2(n637), .ZN(n478) );
  INV_X1 U391 ( .A(KEYINPUT98), .ZN(n401) );
  XNOR2_X1 U392 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U393 ( .A(n366), .B(KEYINPUT17), .ZN(n367) );
  INV_X1 U394 ( .A(KEYINPUT39), .ZN(n531) );
  XNOR2_X1 U395 ( .A(n417), .B(KEYINPUT22), .ZN(n458) );
  XNOR2_X1 U396 ( .A(n456), .B(n455), .ZN(n632) );
  INV_X1 U397 ( .A(KEYINPUT106), .ZN(n538) );
  XNOR2_X1 U398 ( .A(n684), .B(n683), .ZN(n685) );
  XOR2_X1 U399 ( .A(n519), .B(KEYINPUT76), .Z(n350) );
  XOR2_X1 U400 ( .A(KEYINPUT71), .B(KEYINPUT16), .Z(n351) );
  XOR2_X1 U401 ( .A(n553), .B(KEYINPUT47), .Z(n352) );
  XOR2_X1 U402 ( .A(n467), .B(KEYINPUT34), .Z(n353) );
  XNOR2_X1 U403 ( .A(n570), .B(KEYINPUT65), .ZN(n354) );
  XNOR2_X2 U404 ( .A(n550), .B(KEYINPUT1), .ZN(n638) );
  XOR2_X2 U405 ( .A(G116), .B(G107), .Z(n384) );
  INV_X1 U406 ( .A(KEYINPUT46), .ZN(n535) );
  INV_X1 U407 ( .A(KEYINPUT78), .ZN(n504) );
  XNOR2_X1 U408 ( .A(n502), .B(KEYINPUT45), .ZN(n572) );
  XNOR2_X1 U409 ( .A(n402), .B(n401), .ZN(n403) );
  NOR2_X1 U410 ( .A1(n349), .A2(n557), .ZN(n546) );
  XNOR2_X1 U411 ( .A(n450), .B(n449), .ZN(n451) );
  INV_X1 U412 ( .A(KEYINPUT2), .ZN(n628) );
  INV_X1 U413 ( .A(KEYINPUT123), .ZN(n683) );
  INV_X1 U414 ( .A(n458), .ZN(n462) );
  NAND2_X1 U415 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U416 ( .A(n539), .B(n538), .ZN(n614) );
  XNOR2_X1 U417 ( .A(n686), .B(n685), .ZN(n687) );
  INV_X1 U418 ( .A(KEYINPUT87), .ZN(n355) );
  XOR2_X1 U419 ( .A(G101), .B(G119), .Z(n358) );
  XNOR2_X1 U420 ( .A(KEYINPUT69), .B(KEYINPUT3), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n438) );
  XNOR2_X1 U422 ( .A(G113), .B(G104), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n359), .B(G122), .ZN(n399) );
  XNOR2_X1 U424 ( .A(n438), .B(n399), .ZN(n360) );
  XOR2_X1 U425 ( .A(KEYINPUT18), .B(KEYINPUT75), .Z(n362) );
  XNOR2_X1 U426 ( .A(n406), .B(n362), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n386), .B(KEYINPUT4), .ZN(n422) );
  XNOR2_X1 U428 ( .A(n363), .B(n422), .ZN(n368) );
  XOR2_X1 U429 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n365) );
  NAND2_X1 U430 ( .A1(G224), .A2(n703), .ZN(n364) );
  XNOR2_X1 U431 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U432 ( .A(G902), .B(KEYINPUT15), .ZN(n568) );
  AND2_X2 U433 ( .A1(n578), .A2(n568), .ZN(n371) );
  OR2_X1 U434 ( .A1(G237), .A2(G902), .ZN(n372) );
  AND2_X1 U435 ( .A1(n372), .A2(G210), .ZN(n370) );
  NAND2_X1 U436 ( .A1(G214), .A2(n372), .ZN(n373) );
  XNOR2_X1 U437 ( .A(KEYINPUT90), .B(n373), .ZN(n544) );
  INV_X1 U438 ( .A(n544), .ZN(n648) );
  NOR2_X1 U439 ( .A1(n506), .A2(n648), .ZN(n375) );
  XOR2_X1 U440 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n549) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n376) );
  XNOR2_X1 U443 ( .A(n376), .B(KEYINPUT14), .ZN(n378) );
  NAND2_X1 U444 ( .A1(n378), .A2(G902), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n377), .B(KEYINPUT91), .ZN(n508) );
  NOR2_X1 U446 ( .A1(G898), .A2(n703), .ZN(n696) );
  NAND2_X1 U447 ( .A1(n508), .A2(n696), .ZN(n380) );
  NAND2_X1 U448 ( .A1(G952), .A2(n378), .ZN(n664) );
  NOR2_X1 U449 ( .A1(G953), .A2(n664), .ZN(n511) );
  INV_X1 U450 ( .A(n511), .ZN(n379) );
  NAND2_X1 U451 ( .A1(n380), .A2(n379), .ZN(n381) );
  NAND2_X1 U452 ( .A1(n549), .A2(n381), .ZN(n383) );
  INV_X1 U453 ( .A(KEYINPUT0), .ZN(n382) );
  XNOR2_X2 U454 ( .A(n383), .B(n382), .ZN(n483) );
  XNOR2_X1 U455 ( .A(G134), .B(n384), .ZN(n388) );
  XOR2_X1 U456 ( .A(G122), .B(KEYINPUT7), .Z(n385) );
  XNOR2_X1 U457 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U458 ( .A(n388), .B(n387), .ZN(n394) );
  XOR2_X1 U459 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n392) );
  NAND2_X1 U460 ( .A1(n703), .A2(G234), .ZN(n390) );
  XNOR2_X1 U461 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n389) );
  XNOR2_X1 U462 ( .A(n390), .B(n389), .ZN(n444) );
  NAND2_X1 U463 ( .A1(G217), .A2(n444), .ZN(n391) );
  XNOR2_X1 U464 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U465 ( .A(n394), .B(n393), .ZN(n679) );
  NOR2_X1 U466 ( .A1(G902), .A2(n679), .ZN(n396) );
  XNOR2_X1 U467 ( .A(KEYINPUT100), .B(G478), .ZN(n395) );
  XOR2_X1 U468 ( .A(n396), .B(n395), .Z(n489) );
  XNOR2_X1 U469 ( .A(KEYINPUT13), .B(G475), .ZN(n469) );
  XOR2_X1 U470 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n398) );
  XNOR2_X1 U471 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n397) );
  XNOR2_X1 U472 ( .A(n398), .B(n397), .ZN(n400) );
  XOR2_X1 U473 ( .A(n400), .B(n399), .Z(n404) );
  NOR2_X1 U474 ( .A1(G953), .A2(G237), .ZN(n434) );
  NAND2_X1 U475 ( .A1(G214), .A2(n434), .ZN(n402) );
  XNOR2_X1 U476 ( .A(n404), .B(n403), .ZN(n409) );
  XNOR2_X1 U477 ( .A(G140), .B(KEYINPUT10), .ZN(n405) );
  XOR2_X1 U478 ( .A(n406), .B(n405), .Z(n701) );
  XNOR2_X1 U479 ( .A(KEYINPUT68), .B(G131), .ZN(n420) );
  XOR2_X1 U480 ( .A(n420), .B(G143), .Z(n407) );
  XNOR2_X1 U481 ( .A(n701), .B(n407), .ZN(n408) );
  XNOR2_X1 U482 ( .A(n409), .B(n408), .ZN(n589) );
  NOR2_X1 U483 ( .A1(G902), .A2(n589), .ZN(n468) );
  XNOR2_X1 U484 ( .A(n469), .B(n468), .ZN(n486) );
  XOR2_X1 U485 ( .A(n410), .B(KEYINPUT103), .Z(n650) );
  XOR2_X1 U486 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n412) );
  NAND2_X1 U487 ( .A1(G234), .A2(n568), .ZN(n411) );
  XNOR2_X1 U488 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U489 ( .A(KEYINPUT92), .B(n413), .ZN(n454) );
  NAND2_X1 U490 ( .A1(G221), .A2(n454), .ZN(n414) );
  XNOR2_X1 U491 ( .A(n414), .B(KEYINPUT21), .ZN(n631) );
  INV_X1 U492 ( .A(n631), .ZN(n415) );
  AND2_X1 U493 ( .A1(n650), .A2(n415), .ZN(n416) );
  NAND2_X1 U494 ( .A1(n483), .A2(n416), .ZN(n417) );
  INV_X1 U495 ( .A(G137), .ZN(n418) );
  XNOR2_X1 U496 ( .A(n418), .B(G134), .ZN(n419) );
  XNOR2_X1 U497 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U498 ( .A(n422), .B(n421), .ZN(n700) );
  XNOR2_X1 U499 ( .A(n700), .B(G146), .ZN(n440) );
  NAND2_X1 U500 ( .A1(n703), .A2(G227), .ZN(n423) );
  XNOR2_X1 U501 ( .A(n423), .B(KEYINPUT74), .ZN(n424) );
  XNOR2_X1 U502 ( .A(n425), .B(n424), .ZN(n429) );
  XNOR2_X1 U503 ( .A(G104), .B(G101), .ZN(n427) );
  XNOR2_X1 U504 ( .A(G140), .B(G107), .ZN(n426) );
  XNOR2_X1 U505 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U506 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U507 ( .A(n440), .B(n430), .ZN(n675) );
  OR2_X1 U508 ( .A1(n675), .A2(G902), .ZN(n431) );
  XNOR2_X2 U509 ( .A(n431), .B(G469), .ZN(n550) );
  NOR2_X2 U510 ( .A1(n458), .A2(n638), .ZN(n497) );
  XOR2_X1 U511 ( .A(KEYINPUT72), .B(KEYINPUT5), .Z(n433) );
  XNOR2_X1 U512 ( .A(G113), .B(G116), .ZN(n432) );
  XNOR2_X1 U513 ( .A(n433), .B(n432), .ZN(n436) );
  NAND2_X1 U514 ( .A1(n434), .A2(G210), .ZN(n435) );
  XNOR2_X1 U515 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U516 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U517 ( .A(n440), .B(n439), .ZN(n594) );
  XNOR2_X2 U518 ( .A(n441), .B(G472), .ZN(n635) );
  NAND2_X1 U519 ( .A1(n497), .A2(n525), .ZN(n443) );
  INV_X1 U520 ( .A(KEYINPUT64), .ZN(n442) );
  XNOR2_X1 U521 ( .A(n443), .B(n442), .ZN(n457) );
  NAND2_X1 U522 ( .A1(G221), .A2(n444), .ZN(n450) );
  XOR2_X1 U523 ( .A(G110), .B(G128), .Z(n446) );
  XNOR2_X1 U524 ( .A(G119), .B(G137), .ZN(n445) );
  XNOR2_X1 U525 ( .A(n446), .B(n445), .ZN(n448) );
  XOR2_X1 U526 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n447) );
  XNOR2_X1 U527 ( .A(n451), .B(n701), .ZN(n684) );
  NOR2_X1 U528 ( .A1(G902), .A2(n684), .ZN(n453) );
  XNOR2_X1 U529 ( .A(KEYINPUT25), .B(KEYINPUT73), .ZN(n452) );
  XNOR2_X1 U530 ( .A(n453), .B(n452), .ZN(n456) );
  NAND2_X1 U531 ( .A1(n454), .A2(G217), .ZN(n455) );
  AND2_X1 U532 ( .A1(n457), .A2(n632), .ZN(n607) );
  NAND2_X1 U533 ( .A1(n638), .A2(n632), .ZN(n460) );
  INV_X1 U534 ( .A(KEYINPUT6), .ZN(n459) );
  XNOR2_X1 U535 ( .A(n635), .B(n459), .ZN(n540) );
  NOR2_X1 U536 ( .A1(n460), .A2(n540), .ZN(n461) );
  XNOR2_X1 U537 ( .A(n463), .B(KEYINPUT32), .ZN(n715) );
  INV_X1 U538 ( .A(n715), .ZN(n464) );
  NOR2_X1 U539 ( .A1(n607), .A2(n464), .ZN(n474) );
  NOR2_X1 U540 ( .A1(n632), .A2(n631), .ZN(n637) );
  NAND2_X1 U541 ( .A1(n478), .A2(n540), .ZN(n466) );
  XNOR2_X1 U542 ( .A(KEYINPUT84), .B(KEYINPUT33), .ZN(n465) );
  NAND2_X1 U543 ( .A1(n483), .A2(n658), .ZN(n467) );
  XOR2_X1 U544 ( .A(n469), .B(n468), .Z(n490) );
  INV_X1 U545 ( .A(n489), .ZN(n487) );
  NOR2_X1 U546 ( .A1(n490), .A2(n487), .ZN(n470) );
  XNOR2_X1 U547 ( .A(n470), .B(KEYINPUT105), .ZN(n519) );
  NAND2_X1 U548 ( .A1(n353), .A2(n350), .ZN(n473) );
  INV_X1 U549 ( .A(KEYINPUT80), .ZN(n471) );
  XNOR2_X1 U550 ( .A(n471), .B(KEYINPUT35), .ZN(n472) );
  XNOR2_X1 U551 ( .A(n473), .B(n472), .ZN(n588) );
  NAND2_X1 U552 ( .A1(n474), .A2(n588), .ZN(n477) );
  INV_X1 U553 ( .A(KEYINPUT44), .ZN(n475) );
  AND2_X1 U554 ( .A1(n475), .A2(KEYINPUT70), .ZN(n476) );
  XNOR2_X1 U555 ( .A(n477), .B(n476), .ZN(n501) );
  XOR2_X1 U556 ( .A(KEYINPUT95), .B(KEYINPUT31), .Z(n481) );
  NAND2_X1 U557 ( .A1(n478), .A2(n635), .ZN(n479) );
  XOR2_X1 U558 ( .A(KEYINPUT94), .B(n479), .Z(n644) );
  NAND2_X1 U559 ( .A1(n644), .A2(n483), .ZN(n480) );
  XNOR2_X1 U560 ( .A(n481), .B(n480), .ZN(n620) );
  INV_X1 U561 ( .A(n620), .ZN(n485) );
  NAND2_X1 U562 ( .A1(n637), .A2(n550), .ZN(n514) );
  NOR2_X1 U563 ( .A1(n514), .A2(n635), .ZN(n482) );
  AND2_X1 U564 ( .A1(n483), .A2(n482), .ZN(n603) );
  INV_X1 U565 ( .A(n603), .ZN(n484) );
  NAND2_X1 U566 ( .A1(n485), .A2(n484), .ZN(n492) );
  NAND2_X1 U567 ( .A1(n487), .A2(n486), .ZN(n488) );
  NAND2_X1 U568 ( .A1(n490), .A2(n489), .ZN(n608) );
  XOR2_X1 U569 ( .A(KEYINPUT102), .B(n608), .Z(n562) );
  NOR2_X1 U570 ( .A1(n539), .A2(n562), .ZN(n653) );
  INV_X1 U571 ( .A(n653), .ZN(n491) );
  NAND2_X1 U572 ( .A1(n492), .A2(n491), .ZN(n495) );
  INV_X1 U573 ( .A(KEYINPUT70), .ZN(n493) );
  NAND2_X1 U574 ( .A1(n493), .A2(KEYINPUT44), .ZN(n494) );
  AND2_X1 U575 ( .A1(n495), .A2(n494), .ZN(n499) );
  NOR2_X1 U576 ( .A1(n540), .A2(n632), .ZN(n496) );
  NAND2_X1 U577 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U578 ( .A(n498), .B(KEYINPUT104), .ZN(n714) );
  AND2_X1 U579 ( .A1(n499), .A2(n714), .ZN(n500) );
  NAND2_X1 U580 ( .A1(n501), .A2(n500), .ZN(n502) );
  INV_X1 U581 ( .A(n568), .ZN(n503) );
  NAND2_X1 U582 ( .A1(n572), .A2(n503), .ZN(n505) );
  XNOR2_X1 U583 ( .A(n505), .B(n504), .ZN(n567) );
  INV_X1 U584 ( .A(n506), .ZN(n507) );
  NAND2_X1 U585 ( .A1(G953), .A2(n508), .ZN(n509) );
  NOR2_X1 U586 ( .A1(G900), .A2(n509), .ZN(n510) );
  NOR2_X1 U587 ( .A1(n511), .A2(n510), .ZN(n523) );
  NOR2_X1 U588 ( .A1(n648), .A2(n525), .ZN(n512) );
  XOR2_X1 U589 ( .A(KEYINPUT30), .B(n512), .Z(n513) );
  NOR2_X1 U590 ( .A1(n523), .A2(n513), .ZN(n516) );
  INV_X1 U591 ( .A(n514), .ZN(n515) );
  NAND2_X1 U592 ( .A1(n516), .A2(n515), .ZN(n530) );
  NOR2_X1 U593 ( .A1(n349), .A2(n530), .ZN(n517) );
  XNOR2_X1 U594 ( .A(n517), .B(KEYINPUT107), .ZN(n518) );
  NOR2_X1 U595 ( .A1(n519), .A2(n518), .ZN(n612) );
  NOR2_X1 U596 ( .A1(n647), .A2(n648), .ZN(n520) );
  XNOR2_X1 U597 ( .A(n520), .B(KEYINPUT109), .ZN(n652) );
  INV_X1 U598 ( .A(n650), .ZN(n521) );
  NOR2_X1 U599 ( .A1(n652), .A2(n521), .ZN(n522) );
  XNOR2_X1 U600 ( .A(n522), .B(KEYINPUT41), .ZN(n630) );
  NOR2_X1 U601 ( .A1(n523), .A2(n631), .ZN(n524) );
  NAND2_X1 U602 ( .A1(n632), .A2(n524), .ZN(n542) );
  NOR2_X1 U603 ( .A1(n542), .A2(n525), .ZN(n526) );
  XOR2_X1 U604 ( .A(KEYINPUT28), .B(n526), .Z(n552) );
  INV_X1 U605 ( .A(n552), .ZN(n527) );
  NAND2_X1 U606 ( .A1(n527), .A2(n550), .ZN(n528) );
  NOR2_X1 U607 ( .A1(n630), .A2(n528), .ZN(n529) );
  XNOR2_X1 U608 ( .A(n529), .B(KEYINPUT42), .ZN(n716) );
  XOR2_X1 U609 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n534) );
  NOR2_X1 U610 ( .A1(n530), .A2(n647), .ZN(n532) );
  XNOR2_X1 U611 ( .A(n532), .B(n531), .ZN(n561) );
  NAND2_X1 U612 ( .A1(n561), .A2(n539), .ZN(n533) );
  XNOR2_X1 U613 ( .A(n534), .B(n533), .ZN(n711) );
  NOR2_X1 U614 ( .A1(n716), .A2(n711), .ZN(n536) );
  XNOR2_X1 U615 ( .A(n536), .B(n535), .ZN(n537) );
  NOR2_X1 U616 ( .A1(n612), .A2(n537), .ZN(n555) );
  INV_X1 U617 ( .A(n614), .ZN(n617) );
  NAND2_X1 U618 ( .A1(n540), .A2(n617), .ZN(n541) );
  NOR2_X1 U619 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U620 ( .A1(n544), .A2(n543), .ZN(n557) );
  XNOR2_X1 U621 ( .A(KEYINPUT110), .B(KEYINPUT36), .ZN(n545) );
  XNOR2_X1 U622 ( .A(n546), .B(n545), .ZN(n547) );
  NAND2_X1 U623 ( .A1(n547), .A2(n638), .ZN(n548) );
  XNOR2_X1 U624 ( .A(n548), .B(KEYINPUT111), .ZN(n712) );
  NAND2_X1 U625 ( .A1(n549), .A2(n550), .ZN(n551) );
  OR2_X1 U626 ( .A1(n552), .A2(n551), .ZN(n613) );
  NOR2_X1 U627 ( .A1(n653), .A2(n613), .ZN(n553) );
  NOR2_X1 U628 ( .A1(n712), .A2(n352), .ZN(n554) );
  AND2_X1 U629 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U630 ( .A(n556), .B(KEYINPUT48), .ZN(n565) );
  OR2_X1 U631 ( .A1(n557), .A2(n638), .ZN(n558) );
  XNOR2_X1 U632 ( .A(n558), .B(KEYINPUT43), .ZN(n560) );
  NAND2_X1 U633 ( .A1(n560), .A2(n349), .ZN(n623) );
  AND2_X1 U634 ( .A1(n562), .A2(n561), .ZN(n622) );
  INV_X1 U635 ( .A(n622), .ZN(n563) );
  AND2_X1 U636 ( .A1(n623), .A2(n563), .ZN(n564) );
  NAND2_X1 U637 ( .A1(n565), .A2(n564), .ZN(n702) );
  INV_X1 U638 ( .A(n702), .ZN(n566) );
  NAND2_X1 U639 ( .A1(n567), .A2(n566), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n568), .B(KEYINPUT79), .ZN(n569) );
  AND2_X1 U641 ( .A1(n569), .A2(KEYINPUT2), .ZN(n570) );
  NOR2_X1 U642 ( .A1(n702), .A2(n628), .ZN(n573) );
  BUF_X1 U643 ( .A(n572), .Z(n625) );
  NAND2_X1 U644 ( .A1(n573), .A2(n625), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n348), .A2(G210), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n576) );
  XNOR2_X1 U647 ( .A(n576), .B(KEYINPUT55), .ZN(n577) );
  XOR2_X1 U648 ( .A(n577), .B(KEYINPUT121), .Z(n580) );
  XNOR2_X1 U649 ( .A(n578), .B(KEYINPUT54), .ZN(n579) );
  XNOR2_X1 U650 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U651 ( .A(n582), .B(n581), .ZN(n585) );
  INV_X1 U652 ( .A(G952), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n583), .A2(G953), .ZN(n584) );
  XNOR2_X1 U654 ( .A(n584), .B(KEYINPUT86), .ZN(n597) );
  NAND2_X1 U655 ( .A1(n585), .A2(n597), .ZN(n587) );
  INV_X1 U656 ( .A(KEYINPUT56), .ZN(n586) );
  XNOR2_X1 U657 ( .A(n587), .B(n586), .ZN(G51) );
  XNOR2_X1 U658 ( .A(n588), .B(G122), .ZN(G24) );
  NAND2_X1 U659 ( .A1(n682), .A2(G475), .ZN(n591) );
  XOR2_X1 U660 ( .A(n589), .B(KEYINPUT59), .Z(n590) );
  XNOR2_X1 U661 ( .A(n591), .B(n590), .ZN(n592) );
  INV_X1 U662 ( .A(n597), .ZN(n688) );
  NOR2_X2 U663 ( .A1(n592), .A2(n688), .ZN(n593) );
  XNOR2_X1 U664 ( .A(n593), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U665 ( .A1(n348), .A2(G472), .ZN(n596) );
  XOR2_X1 U666 ( .A(KEYINPUT62), .B(n594), .Z(n595) );
  XNOR2_X1 U667 ( .A(n596), .B(n595), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n601) );
  XNOR2_X1 U669 ( .A(KEYINPUT85), .B(KEYINPUT63), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n599), .B(KEYINPUT81), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n601), .B(n600), .ZN(G57) );
  NAND2_X1 U672 ( .A1(n617), .A2(n603), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(G104), .ZN(G6) );
  XOR2_X1 U674 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n605) );
  INV_X1 U675 ( .A(n608), .ZN(n619) );
  NAND2_X1 U676 ( .A1(n603), .A2(n619), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n605), .B(n604), .ZN(n606) );
  XNOR2_X1 U678 ( .A(G107), .B(n606), .ZN(G9) );
  XOR2_X1 U679 ( .A(G110), .B(n607), .Z(G12) );
  NOR2_X1 U680 ( .A1(n608), .A2(n613), .ZN(n610) );
  XNOR2_X1 U681 ( .A(KEYINPUT112), .B(KEYINPUT29), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U683 ( .A(G128), .B(n611), .ZN(G30) );
  XOR2_X1 U684 ( .A(G143), .B(n612), .Z(G45) );
  NOR2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n616) );
  XNOR2_X1 U686 ( .A(G146), .B(KEYINPUT113), .ZN(n615) );
  XNOR2_X1 U687 ( .A(n616), .B(n615), .ZN(G48) );
  NAND2_X1 U688 ( .A1(n617), .A2(n620), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(G113), .ZN(G15) );
  NAND2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U691 ( .A(n621), .B(G116), .ZN(G18) );
  XOR2_X1 U692 ( .A(G134), .B(n622), .Z(G36) );
  XNOR2_X1 U693 ( .A(G140), .B(KEYINPUT114), .ZN(n624) );
  XNOR2_X1 U694 ( .A(n624), .B(n623), .ZN(G42) );
  INV_X1 U695 ( .A(n625), .ZN(n626) );
  NOR2_X1 U696 ( .A1(n626), .A2(n702), .ZN(n627) );
  NOR2_X1 U697 ( .A1(n627), .A2(KEYINPUT77), .ZN(n629) );
  XNOR2_X1 U698 ( .A(n629), .B(n628), .ZN(n669) );
  AND2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U700 ( .A(KEYINPUT49), .B(n633), .Z(n634) );
  NOR2_X1 U701 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U702 ( .A(KEYINPUT115), .B(n636), .ZN(n641) );
  NOR2_X1 U703 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U704 ( .A(n639), .B(KEYINPUT50), .ZN(n640) );
  NOR2_X1 U705 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U706 ( .A(n642), .B(KEYINPUT116), .ZN(n643) );
  NOR2_X1 U707 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U708 ( .A(KEYINPUT51), .B(n645), .Z(n646) );
  NOR2_X1 U709 ( .A1(n630), .A2(n646), .ZN(n661) );
  NAND2_X1 U710 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U711 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U712 ( .A(KEYINPUT117), .B(n651), .ZN(n656) );
  NOR2_X1 U713 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U714 ( .A(n654), .B(KEYINPUT118), .ZN(n655) );
  NOR2_X1 U715 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U716 ( .A(KEYINPUT119), .B(n657), .Z(n659) );
  INV_X1 U717 ( .A(n658), .ZN(n665) );
  NOR2_X1 U718 ( .A1(n659), .A2(n665), .ZN(n660) );
  NOR2_X1 U719 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U720 ( .A(n662), .B(KEYINPUT52), .ZN(n663) );
  NOR2_X1 U721 ( .A1(n664), .A2(n663), .ZN(n667) );
  NOR2_X1 U722 ( .A1(n630), .A2(n665), .ZN(n666) );
  NOR2_X1 U723 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U724 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U725 ( .A1(G953), .A2(n670), .ZN(n672) );
  XNOR2_X1 U726 ( .A(KEYINPUT53), .B(KEYINPUT120), .ZN(n671) );
  XNOR2_X1 U727 ( .A(n672), .B(n671), .ZN(G75) );
  NAND2_X1 U728 ( .A1(n348), .A2(G469), .ZN(n677) );
  XOR2_X1 U729 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n673) );
  XNOR2_X1 U730 ( .A(n673), .B(KEYINPUT122), .ZN(n674) );
  XNOR2_X1 U731 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U732 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U733 ( .A1(n688), .A2(n678), .ZN(G54) );
  NAND2_X1 U734 ( .A1(n348), .A2(G478), .ZN(n680) );
  XNOR2_X1 U735 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U736 ( .A1(n688), .A2(n681), .ZN(G63) );
  NAND2_X1 U737 ( .A1(n348), .A2(G217), .ZN(n686) );
  NOR2_X1 U738 ( .A1(n688), .A2(n687), .ZN(G66) );
  NAND2_X1 U739 ( .A1(n625), .A2(n703), .ZN(n694) );
  NAND2_X1 U740 ( .A1(G224), .A2(G953), .ZN(n689) );
  XNOR2_X1 U741 ( .A(n689), .B(KEYINPUT61), .ZN(n690) );
  XNOR2_X1 U742 ( .A(KEYINPUT124), .B(n690), .ZN(n691) );
  NAND2_X1 U743 ( .A1(n691), .A2(G898), .ZN(n692) );
  XOR2_X1 U744 ( .A(KEYINPUT125), .B(n692), .Z(n693) );
  NAND2_X1 U745 ( .A1(n694), .A2(n693), .ZN(n698) );
  NOR2_X1 U746 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U747 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U748 ( .A(KEYINPUT126), .B(n699), .ZN(G69) );
  XNOR2_X1 U749 ( .A(n701), .B(n700), .ZN(n705) );
  XNOR2_X1 U750 ( .A(n702), .B(n705), .ZN(n704) );
  NAND2_X1 U751 ( .A1(n704), .A2(n703), .ZN(n710) );
  XNOR2_X1 U752 ( .A(n705), .B(G227), .ZN(n706) );
  NAND2_X1 U753 ( .A1(n706), .A2(G900), .ZN(n707) );
  XOR2_X1 U754 ( .A(KEYINPUT127), .B(n707), .Z(n708) );
  NAND2_X1 U755 ( .A1(G953), .A2(n708), .ZN(n709) );
  NAND2_X1 U756 ( .A1(n710), .A2(n709), .ZN(G72) );
  XOR2_X1 U757 ( .A(G131), .B(n711), .Z(G33) );
  XNOR2_X1 U758 ( .A(G125), .B(n712), .ZN(n713) );
  XNOR2_X1 U759 ( .A(n713), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U760 ( .A(G101), .B(n714), .ZN(G3) );
  XNOR2_X1 U761 ( .A(n715), .B(G119), .ZN(G21) );
  XOR2_X1 U762 ( .A(G137), .B(n716), .Z(G39) );
endmodule

