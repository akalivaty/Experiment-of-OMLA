

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759;

  INV_X1 U365 ( .A(n601), .ZN(n348) );
  NOR2_X1 U366 ( .A1(n681), .A2(n588), .ZN(n405) );
  NOR2_X1 U367 ( .A1(n622), .A2(n516), .ZN(n430) );
  INV_X1 U368 ( .A(n464), .ZN(n346) );
  XNOR2_X1 U369 ( .A(n400), .B(n467), .ZN(n499) );
  XNOR2_X1 U370 ( .A(n466), .B(n468), .ZN(n400) );
  XNOR2_X1 U371 ( .A(n501), .B(n457), .ZN(n545) );
  XNOR2_X1 U372 ( .A(n435), .B(G131), .ZN(n531) );
  INV_X1 U373 ( .A(KEYINPUT71), .ZN(n435) );
  INV_X1 U374 ( .A(G143), .ZN(n456) );
  INV_X2 U375 ( .A(G953), .ZN(n747) );
  AND2_X2 U376 ( .A1(n376), .A2(KEYINPUT60), .ZN(n375) );
  XNOR2_X2 U377 ( .A(n347), .B(n346), .ZN(n385) );
  OR2_X2 U378 ( .A1(n715), .A2(G902), .ZN(n347) );
  INV_X1 U379 ( .A(n349), .ZN(n731) );
  NAND2_X1 U380 ( .A1(n380), .A2(n349), .ZN(n379) );
  XNOR2_X2 U381 ( .A(n602), .B(n348), .ZN(n349) );
  NOR2_X1 U382 ( .A1(n567), .A2(n616), .ZN(n568) );
  NAND2_X1 U383 ( .A1(n439), .A2(n597), .ZN(n598) );
  XNOR2_X1 U384 ( .A(n499), .B(n498), .ZN(n724) );
  INV_X2 U385 ( .A(n710), .ZN(n719) );
  XNOR2_X2 U386 ( .A(KEYINPUT99), .B(n571), .ZN(n627) );
  XNOR2_X2 U387 ( .A(n405), .B(KEYINPUT31), .ZN(n664) );
  NOR2_X1 U388 ( .A1(n684), .A2(n588), .ZN(n432) );
  XNOR2_X1 U389 ( .A(n385), .B(KEYINPUT1), .ZN(n577) );
  XNOR2_X1 U390 ( .A(n537), .B(n536), .ZN(n590) );
  INV_X1 U391 ( .A(KEYINPUT87), .ZN(n433) );
  NAND2_X1 U392 ( .A1(n383), .A2(n381), .ZN(n669) );
  NAND2_X1 U393 ( .A1(n360), .A2(n350), .ZN(n746) );
  NOR2_X1 U394 ( .A1(n388), .A2(n387), .ZN(n386) );
  XNOR2_X1 U395 ( .A(n615), .B(KEYINPUT42), .ZN(n758) );
  XNOR2_X1 U396 ( .A(n611), .B(n610), .ZN(n701) );
  NOR2_X1 U397 ( .A1(n629), .A2(n632), .ZN(n661) );
  NOR2_X1 U398 ( .A1(n633), .A2(n632), .ZN(n658) );
  XNOR2_X1 U399 ( .A(n550), .B(G478), .ZN(n570) );
  NOR2_X1 U400 ( .A1(n717), .A2(G902), .ZN(n550) );
  XNOR2_X1 U401 ( .A(n531), .B(G137), .ZN(n434) );
  XOR2_X1 U402 ( .A(KEYINPUT4), .B(KEYINPUT68), .Z(n745) );
  XNOR2_X1 U403 ( .A(G116), .B(G107), .ZN(n541) );
  XNOR2_X1 U404 ( .A(KEYINPUT16), .B(G122), .ZN(n497) );
  XNOR2_X2 U405 ( .A(n384), .B(KEYINPUT64), .ZN(n710) );
  XNOR2_X1 U406 ( .A(n361), .B(n637), .ZN(n360) );
  INV_X1 U407 ( .A(G107), .ZN(n454) );
  XNOR2_X1 U408 ( .A(G104), .B(G110), .ZN(n455) );
  NAND2_X1 U409 ( .A1(n409), .A2(KEYINPUT44), .ZN(n408) );
  XNOR2_X1 U410 ( .A(n404), .B(n353), .ZN(n614) );
  OR2_X1 U411 ( .A1(n613), .A2(n612), .ZN(n404) );
  NAND2_X1 U412 ( .A1(n689), .A2(n396), .ZN(n395) );
  XOR2_X1 U413 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n524) );
  NOR2_X1 U414 ( .A1(n664), .A2(n395), .ZN(n387) );
  NOR2_X1 U415 ( .A1(KEYINPUT67), .A2(n634), .ZN(n635) );
  INV_X1 U416 ( .A(G134), .ZN(n457) );
  XNOR2_X1 U417 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U418 ( .A(n495), .B(n494), .ZN(n674) );
  XNOR2_X1 U419 ( .A(n493), .B(KEYINPUT25), .ZN(n494) );
  NOR2_X1 U420 ( .A1(G902), .A2(n720), .ZN(n495) );
  INV_X1 U421 ( .A(G146), .ZN(n453) );
  INV_X1 U422 ( .A(G140), .ZN(n458) );
  XNOR2_X1 U423 ( .A(n397), .B(n511), .ZN(n713) );
  XNOR2_X1 U424 ( .A(n724), .B(n508), .ZN(n397) );
  INV_X1 U425 ( .A(n746), .ZN(n380) );
  NOR2_X1 U426 ( .A1(n746), .A2(KEYINPUT2), .ZN(n382) );
  BUF_X1 U427 ( .A(n684), .Z(n703) );
  XNOR2_X1 U428 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n610) );
  NOR2_X1 U429 ( .A1(n690), .A2(n688), .ZN(n611) );
  NOR2_X1 U430 ( .A1(n626), .A2(n618), .ZN(n619) );
  NOR2_X1 U431 ( .A1(n603), .A2(n407), .ZN(n605) );
  BUF_X1 U432 ( .A(n622), .Z(n407) );
  OR2_X1 U433 ( .A1(n649), .A2(G902), .ZN(n475) );
  INV_X1 U434 ( .A(n674), .ZN(n582) );
  NAND2_X1 U435 ( .A1(n428), .A2(n673), .ZN(n427) );
  NAND2_X1 U436 ( .A1(n417), .A2(n356), .ZN(n423) );
  OR2_X1 U437 ( .A1(n645), .A2(G475), .ZN(n424) );
  NOR2_X1 U438 ( .A1(n645), .A2(KEYINPUT60), .ZN(n420) );
  NOR2_X1 U439 ( .A1(n369), .A2(n723), .ZN(n368) );
  NAND2_X1 U440 ( .A1(n392), .A2(n390), .ZN(n388) );
  NAND2_X1 U441 ( .A1(n391), .A2(KEYINPUT100), .ZN(n390) );
  NAND2_X1 U442 ( .A1(n394), .A2(n393), .ZN(n392) );
  XNOR2_X1 U443 ( .A(G143), .B(G113), .ZN(n528) );
  XOR2_X1 U444 ( .A(G122), .B(G104), .Z(n529) );
  XNOR2_X1 U445 ( .A(n526), .B(n451), .ZN(n527) );
  XNOR2_X1 U446 ( .A(KEYINPUT92), .B(KEYINPUT12), .ZN(n523) );
  INV_X1 U447 ( .A(G237), .ZN(n512) );
  INV_X1 U448 ( .A(G902), .ZN(n535) );
  XNOR2_X1 U449 ( .A(n621), .B(n363), .ZN(n362) );
  AND2_X1 U450 ( .A1(n450), .A2(n636), .ZN(n364) );
  INV_X1 U451 ( .A(KEYINPUT46), .ZN(n363) );
  XNOR2_X1 U452 ( .A(KEYINPUT86), .B(KEYINPUT15), .ZN(n490) );
  XNOR2_X1 U453 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n504) );
  NAND2_X1 U454 ( .A1(n594), .A2(n372), .ZN(n409) );
  NAND2_X1 U455 ( .A1(G234), .A2(G237), .ZN(n517) );
  XNOR2_X1 U456 ( .A(n609), .B(KEYINPUT108), .ZN(n690) );
  NAND2_X1 U457 ( .A1(n686), .A2(n685), .ZN(n609) );
  XNOR2_X1 U458 ( .A(n552), .B(n551), .ZN(n688) );
  OR2_X1 U459 ( .A1(n590), .A2(n589), .ZN(n552) );
  INV_X1 U460 ( .A(KEYINPUT38), .ZN(n608) );
  INV_X1 U461 ( .A(KEYINPUT19), .ZN(n440) );
  INV_X1 U462 ( .A(n688), .ZN(n428) );
  XOR2_X1 U463 ( .A(KEYINPUT89), .B(KEYINPUT5), .Z(n470) );
  XNOR2_X1 U464 ( .A(G119), .B(G116), .ZN(n467) );
  XNOR2_X1 U465 ( .A(n479), .B(n478), .ZN(n540) );
  XOR2_X1 U466 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n478) );
  XNOR2_X1 U467 ( .A(n477), .B(n476), .ZN(n479) );
  INV_X1 U468 ( .A(KEYINPUT70), .ZN(n476) );
  XNOR2_X1 U469 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n483) );
  XNOR2_X1 U470 ( .A(G128), .B(G137), .ZN(n481) );
  XOR2_X1 U471 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n542) );
  AND2_X1 U472 ( .A1(n645), .A2(G475), .ZN(n425) );
  XNOR2_X1 U473 ( .A(n399), .B(n587), .ZN(n684) );
  XNOR2_X1 U474 ( .A(n446), .B(KEYINPUT30), .ZN(n445) );
  NOR2_X1 U475 ( .A1(n612), .A2(n516), .ZN(n446) );
  NOR2_X1 U476 ( .A1(n710), .A2(n648), .ZN(n443) );
  XNOR2_X1 U477 ( .A(n403), .B(n461), .ZN(n715) );
  XNOR2_X1 U478 ( .A(n741), .B(n460), .ZN(n403) );
  XNOR2_X1 U479 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U480 ( .A1(n349), .A2(n382), .ZN(n381) );
  NAND2_X1 U481 ( .A1(n701), .A2(n631), .ZN(n615) );
  XNOR2_X1 U482 ( .A(n398), .B(n620), .ZN(n757) );
  OR2_X1 U483 ( .A1(n638), .A2(n662), .ZN(n398) );
  XNOR2_X1 U484 ( .A(KEYINPUT83), .B(KEYINPUT36), .ZN(n604) );
  XNOR2_X1 U485 ( .A(n431), .B(KEYINPUT102), .ZN(n759) );
  AND2_X1 U486 ( .A1(n378), .A2(n419), .ZN(n377) );
  INV_X1 U487 ( .A(KEYINPUT56), .ZN(n447) );
  NAND2_X1 U488 ( .A1(n366), .A2(n714), .ZN(n365) );
  INV_X1 U489 ( .A(n645), .ZN(n421) );
  AND2_X1 U490 ( .A1(n640), .A2(n639), .ZN(n350) );
  AND2_X1 U491 ( .A1(n671), .A2(n583), .ZN(n351) );
  AND2_X1 U492 ( .A1(n652), .A2(KEYINPUT100), .ZN(n352) );
  XNOR2_X1 U493 ( .A(KEYINPUT28), .B(KEYINPUT106), .ZN(n353) );
  XNOR2_X1 U494 ( .A(KEYINPUT62), .B(n649), .ZN(n354) );
  AND2_X1 U495 ( .A1(n449), .A2(G210), .ZN(n355) );
  AND2_X1 U496 ( .A1(n424), .A2(n448), .ZN(n356) );
  NAND2_X1 U497 ( .A1(n596), .A2(KEYINPUT66), .ZN(n357) );
  INV_X1 U498 ( .A(n723), .ZN(n448) );
  XNOR2_X1 U499 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n358) );
  XOR2_X1 U500 ( .A(G122), .B(KEYINPUT126), .Z(n359) );
  NAND2_X1 U501 ( .A1(n585), .A2(n586), .ZN(n399) );
  NOR2_X1 U502 ( .A1(n414), .A2(n411), .ZN(n410) );
  NAND2_X1 U503 ( .A1(n364), .A2(n362), .ZN(n361) );
  NAND2_X1 U504 ( .A1(n367), .A2(n365), .ZN(n371) );
  INV_X1 U505 ( .A(n719), .ZN(n366) );
  AND2_X1 U506 ( .A1(n370), .A2(n368), .ZN(n367) );
  NOR2_X1 U507 ( .A1(n449), .A2(G210), .ZN(n369) );
  NAND2_X1 U508 ( .A1(n719), .A2(n355), .ZN(n370) );
  XNOR2_X1 U509 ( .A(n371), .B(n447), .ZN(G51) );
  NOR2_X1 U510 ( .A1(n413), .A2(n357), .ZN(n599) );
  INV_X1 U511 ( .A(n413), .ZN(n372) );
  XNOR2_X1 U512 ( .A(n413), .B(n359), .ZN(G24) );
  XNOR2_X2 U513 ( .A(n592), .B(KEYINPUT35), .ZN(n413) );
  NAND2_X1 U514 ( .A1(n373), .A2(n560), .ZN(n561) );
  NAND2_X1 U515 ( .A1(n373), .A2(n351), .ZN(n431) );
  NAND2_X1 U516 ( .A1(n373), .A2(n555), .ZN(n597) );
  XNOR2_X2 U517 ( .A(n426), .B(KEYINPUT22), .ZN(n373) );
  NAND2_X1 U518 ( .A1(n377), .A2(n374), .ZN(G60) );
  NAND2_X1 U519 ( .A1(n418), .A2(n375), .ZN(n374) );
  NAND2_X1 U520 ( .A1(n422), .A2(n421), .ZN(n376) );
  NAND2_X1 U521 ( .A1(n423), .A2(n647), .ZN(n378) );
  NAND2_X1 U522 ( .A1(n379), .A2(KEYINPUT2), .ZN(n383) );
  NAND2_X1 U523 ( .A1(n669), .A2(n642), .ZN(n384) );
  NOR2_X1 U524 ( .A1(n385), .A2(n670), .ZN(n617) );
  NOR2_X1 U525 ( .A1(n614), .A2(n385), .ZN(n631) );
  NAND2_X1 U526 ( .A1(n386), .A2(n389), .ZN(n584) );
  NAND2_X1 U527 ( .A1(n664), .A2(n352), .ZN(n389) );
  INV_X1 U528 ( .A(n689), .ZN(n391) );
  INV_X1 U529 ( .A(n395), .ZN(n393) );
  INV_X1 U530 ( .A(n652), .ZN(n394) );
  INV_X1 U531 ( .A(KEYINPUT100), .ZN(n396) );
  XNOR2_X2 U532 ( .A(n561), .B(KEYINPUT32), .ZN(n439) );
  NOR2_X2 U533 ( .A1(n577), .A2(n670), .ZN(n585) );
  XNOR2_X1 U534 ( .A(n430), .B(n440), .ZN(n628) );
  NAND2_X1 U535 ( .A1(n445), .A2(n401), .ZN(n626) );
  AND2_X1 U536 ( .A1(n617), .A2(n444), .ZN(n401) );
  XNOR2_X1 U537 ( .A(n402), .B(n472), .ZN(n649) );
  XNOR2_X1 U538 ( .A(n473), .B(n474), .ZN(n402) );
  NOR2_X1 U539 ( .A1(n755), .A2(n660), .ZN(n450) );
  XNOR2_X1 U540 ( .A(n607), .B(KEYINPUT110), .ZN(n755) );
  AND2_X1 U541 ( .A1(n627), .A2(n406), .ZN(n572) );
  NOR2_X1 U542 ( .A1(n613), .A2(n516), .ZN(n406) );
  NAND2_X1 U543 ( .A1(n413), .A2(n600), .ZN(n412) );
  NAND2_X1 U544 ( .A1(n410), .A2(n408), .ZN(n602) );
  NOR2_X1 U545 ( .A1(n598), .A2(n412), .ZN(n411) );
  NAND2_X1 U546 ( .A1(n415), .A2(n595), .ZN(n414) );
  NAND2_X1 U547 ( .A1(n416), .A2(n599), .ZN(n415) );
  INV_X1 U548 ( .A(n598), .ZN(n416) );
  NAND2_X1 U549 ( .A1(n719), .A2(n425), .ZN(n417) );
  INV_X1 U550 ( .A(n423), .ZN(n418) );
  NAND2_X1 U551 ( .A1(n422), .A2(n420), .ZN(n419) );
  INV_X1 U552 ( .A(n719), .ZN(n422) );
  NOR2_X2 U553 ( .A1(n588), .A2(n427), .ZN(n426) );
  XNOR2_X2 U554 ( .A(n429), .B(n522), .ZN(n588) );
  NAND2_X1 U555 ( .A1(n628), .A2(n520), .ZN(n429) );
  XNOR2_X2 U556 ( .A(n480), .B(KEYINPUT10), .ZN(n740) );
  XNOR2_X1 U557 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U558 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U559 ( .A(n432), .B(KEYINPUT34), .ZN(n591) );
  XNOR2_X2 U560 ( .A(n473), .B(n433), .ZN(n741) );
  XNOR2_X2 U561 ( .A(n545), .B(n434), .ZN(n473) );
  XNOR2_X2 U562 ( .A(n456), .B(G128), .ZN(n501) );
  AND2_X1 U563 ( .A1(n436), .A2(n448), .ZN(G54) );
  XNOR2_X1 U564 ( .A(n438), .B(n437), .ZN(n436) );
  XNOR2_X1 U565 ( .A(n715), .B(n358), .ZN(n437) );
  NAND2_X1 U566 ( .A1(n719), .A2(G469), .ZN(n438) );
  AND2_X1 U567 ( .A1(n593), .A2(n439), .ZN(n594) );
  XNOR2_X1 U568 ( .A(n439), .B(G119), .ZN(G21) );
  XNOR2_X2 U569 ( .A(n514), .B(n513), .ZN(n622) );
  XNOR2_X1 U570 ( .A(n441), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U571 ( .A1(n442), .A2(n448), .ZN(n441) );
  XNOR2_X1 U572 ( .A(n443), .B(n354), .ZN(n442) );
  INV_X1 U573 ( .A(n612), .ZN(n677) );
  INV_X1 U574 ( .A(n616), .ZN(n444) );
  INV_X1 U575 ( .A(n714), .ZN(n449) );
  AND2_X1 U576 ( .A1(G214), .A2(n525), .ZN(n451) );
  INV_X1 U577 ( .A(KEYINPUT48), .ZN(n637) );
  XNOR2_X1 U578 ( .A(n740), .B(n527), .ZN(n534) );
  BUF_X1 U579 ( .A(n724), .Z(n728) );
  XNOR2_X1 U580 ( .A(n605), .B(n604), .ZN(n606) );
  INV_X1 U581 ( .A(G101), .ZN(n452) );
  XNOR2_X1 U582 ( .A(n745), .B(n452), .ZN(n509) );
  XNOR2_X1 U583 ( .A(n509), .B(n453), .ZN(n474) );
  XNOR2_X1 U584 ( .A(n455), .B(n454), .ZN(n726) );
  XNOR2_X1 U585 ( .A(n726), .B(KEYINPUT78), .ZN(n510) );
  XNOR2_X1 U586 ( .A(n474), .B(n510), .ZN(n461) );
  NAND2_X1 U587 ( .A1(G227), .A2(n747), .ZN(n459) );
  XNOR2_X1 U588 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n463) );
  INV_X1 U589 ( .A(G469), .ZN(n462) );
  INV_X1 U590 ( .A(n577), .ZN(n573) );
  XNOR2_X2 U591 ( .A(G113), .B(KEYINPUT75), .ZN(n466) );
  XNOR2_X2 U592 ( .A(KEYINPUT76), .B(KEYINPUT3), .ZN(n468) );
  NOR2_X1 U593 ( .A1(G953), .A2(G237), .ZN(n525) );
  NAND2_X1 U594 ( .A1(n525), .A2(G210), .ZN(n469) );
  XNOR2_X1 U595 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U596 ( .A(n499), .B(n471), .ZN(n472) );
  INV_X1 U597 ( .A(G472), .ZN(n648) );
  XNOR2_X2 U598 ( .A(n475), .B(n648), .ZN(n612) );
  NAND2_X1 U599 ( .A1(G234), .A2(n747), .ZN(n477) );
  NAND2_X1 U600 ( .A1(G221), .A2(n540), .ZN(n489) );
  XOR2_X2 U601 ( .A(G146), .B(G125), .Z(n500) );
  XNOR2_X1 U602 ( .A(n500), .B(G140), .ZN(n480) );
  XOR2_X1 U603 ( .A(G110), .B(G119), .Z(n482) );
  XNOR2_X1 U604 ( .A(n482), .B(n481), .ZN(n486) );
  XOR2_X1 U605 ( .A(KEYINPUT82), .B(KEYINPUT77), .Z(n484) );
  XNOR2_X1 U606 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U607 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U608 ( .A(n740), .B(n487), .ZN(n488) );
  XNOR2_X1 U609 ( .A(n489), .B(n488), .ZN(n720) );
  XNOR2_X1 U610 ( .A(n490), .B(G902), .ZN(n641) );
  NAND2_X1 U611 ( .A1(G234), .A2(n641), .ZN(n492) );
  XNOR2_X1 U612 ( .A(KEYINPUT88), .B(KEYINPUT20), .ZN(n491) );
  XNOR2_X1 U613 ( .A(n492), .B(n491), .ZN(n553) );
  NAND2_X1 U614 ( .A1(G217), .A2(n553), .ZN(n493) );
  NAND2_X1 U615 ( .A1(n612), .A2(n582), .ZN(n496) );
  NOR2_X1 U616 ( .A1(n573), .A2(n496), .ZN(n555) );
  XNOR2_X1 U617 ( .A(n497), .B(KEYINPUT79), .ZN(n498) );
  XNOR2_X1 U618 ( .A(n501), .B(n500), .ZN(n507) );
  XNOR2_X1 U619 ( .A(KEYINPUT80), .B(KEYINPUT84), .ZN(n503) );
  NAND2_X1 U620 ( .A1(n747), .A2(G224), .ZN(n502) );
  XNOR2_X1 U621 ( .A(n503), .B(n502), .ZN(n505) );
  XNOR2_X1 U622 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U623 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U624 ( .A(n510), .B(n509), .ZN(n511) );
  NAND2_X1 U625 ( .A1(n713), .A2(n641), .ZN(n514) );
  NAND2_X1 U626 ( .A1(n535), .A2(n512), .ZN(n515) );
  NAND2_X1 U627 ( .A1(n515), .A2(G210), .ZN(n513) );
  NAND2_X1 U628 ( .A1(n515), .A2(G214), .ZN(n685) );
  INV_X1 U629 ( .A(n685), .ZN(n516) );
  XNOR2_X1 U630 ( .A(n517), .B(KEYINPUT14), .ZN(n518) );
  NAND2_X1 U631 ( .A1(G952), .A2(n518), .ZN(n700) );
  NOR2_X1 U632 ( .A1(n700), .A2(G953), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G902), .A2(n518), .ZN(n562) );
  OR2_X1 U634 ( .A1(n747), .A2(G898), .ZN(n730) );
  NOR2_X1 U635 ( .A1(n562), .A2(n730), .ZN(n519) );
  OR2_X1 U636 ( .A1(n566), .A2(n519), .ZN(n520) );
  INV_X1 U637 ( .A(KEYINPUT65), .ZN(n521) );
  XNOR2_X1 U638 ( .A(n521), .B(KEYINPUT0), .ZN(n522) );
  XNOR2_X1 U639 ( .A(n524), .B(n523), .ZN(n526) );
  XNOR2_X1 U640 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U641 ( .A(n530), .B(KEYINPUT11), .ZN(n532) );
  XNOR2_X1 U642 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U643 ( .A(n534), .B(n533), .ZN(n644) );
  NAND2_X1 U644 ( .A1(n644), .A2(n535), .ZN(n537) );
  XOR2_X1 U645 ( .A(KEYINPUT13), .B(G475), .Z(n536) );
  XOR2_X1 U646 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n539) );
  XNOR2_X1 U647 ( .A(G122), .B(KEYINPUT95), .ZN(n538) );
  XNOR2_X1 U648 ( .A(n539), .B(n538), .ZN(n549) );
  NAND2_X1 U649 ( .A1(G217), .A2(n540), .ZN(n547) );
  XNOR2_X1 U650 ( .A(n541), .B(KEYINPUT96), .ZN(n543) );
  XNOR2_X1 U651 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U652 ( .A(n549), .B(n548), .ZN(n717) );
  INV_X1 U653 ( .A(n570), .ZN(n589) );
  INV_X1 U654 ( .A(KEYINPUT101), .ZN(n551) );
  AND2_X1 U655 ( .A1(n553), .A2(G221), .ZN(n554) );
  XNOR2_X1 U656 ( .A(n554), .B(KEYINPUT21), .ZN(n673) );
  INV_X1 U657 ( .A(n673), .ZN(n567) );
  XNOR2_X1 U658 ( .A(G110), .B(KEYINPUT114), .ZN(n556) );
  XNOR2_X1 U659 ( .A(n597), .B(n556), .ZN(G12) );
  INV_X1 U660 ( .A(n573), .ZN(n671) );
  OR2_X1 U661 ( .A1(n671), .A2(n674), .ZN(n559) );
  XNOR2_X1 U662 ( .A(n612), .B(KEYINPUT6), .ZN(n586) );
  INV_X1 U663 ( .A(KEYINPUT81), .ZN(n557) );
  XNOR2_X1 U664 ( .A(n586), .B(n557), .ZN(n558) );
  NOR2_X1 U665 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U666 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n575) );
  OR2_X1 U667 ( .A1(n747), .A2(n562), .ZN(n563) );
  XNOR2_X1 U668 ( .A(KEYINPUT104), .B(n563), .ZN(n564) );
  NOR2_X1 U669 ( .A1(G900), .A2(n564), .ZN(n565) );
  NOR2_X1 U670 ( .A1(n566), .A2(n565), .ZN(n616) );
  XNOR2_X1 U671 ( .A(KEYINPUT72), .B(n568), .ZN(n569) );
  NAND2_X1 U672 ( .A1(n569), .A2(n582), .ZN(n613) );
  XNOR2_X1 U673 ( .A(n590), .B(KEYINPUT94), .ZN(n580) );
  NAND2_X1 U674 ( .A1(n570), .A2(n580), .ZN(n571) );
  NAND2_X1 U675 ( .A1(n572), .A2(n586), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n603), .A2(n573), .ZN(n574) );
  XNOR2_X1 U677 ( .A(n575), .B(n574), .ZN(n576) );
  NAND2_X1 U678 ( .A1(n576), .A2(n407), .ZN(n639) );
  XNOR2_X1 U679 ( .A(n639), .B(G140), .ZN(G42) );
  NAND2_X1 U680 ( .A1(n674), .A2(n673), .ZN(n670) );
  NAND2_X1 U681 ( .A1(n585), .A2(n677), .ZN(n578) );
  XNOR2_X1 U682 ( .A(n578), .B(KEYINPUT90), .ZN(n681) );
  NAND2_X1 U683 ( .A1(n617), .A2(n612), .ZN(n579) );
  OR2_X1 U684 ( .A1(n579), .A2(n588), .ZN(n652) );
  INV_X1 U685 ( .A(n627), .ZN(n662) );
  INV_X1 U686 ( .A(n580), .ZN(n581) );
  NAND2_X1 U687 ( .A1(n581), .A2(n589), .ZN(n665) );
  NAND2_X1 U688 ( .A1(n662), .A2(n665), .ZN(n689) );
  NOR2_X1 U689 ( .A1(n586), .A2(n582), .ZN(n583) );
  AND2_X1 U690 ( .A1(n584), .A2(n759), .ZN(n595) );
  XNOR2_X1 U691 ( .A(KEYINPUT103), .B(KEYINPUT33), .ZN(n587) );
  AND2_X1 U692 ( .A1(n590), .A2(n589), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n591), .A2(n624), .ZN(n592) );
  AND2_X1 U694 ( .A1(n597), .A2(KEYINPUT66), .ZN(n593) );
  INV_X1 U695 ( .A(KEYINPUT44), .ZN(n596) );
  INV_X1 U696 ( .A(KEYINPUT66), .ZN(n600) );
  INV_X1 U697 ( .A(KEYINPUT45), .ZN(n601) );
  NOR2_X1 U698 ( .A1(n671), .A2(n606), .ZN(n607) );
  XNOR2_X1 U699 ( .A(n622), .B(n608), .ZN(n618) );
  INV_X1 U700 ( .A(n618), .ZN(n686) );
  XOR2_X1 U701 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n620) );
  XNOR2_X1 U702 ( .A(n619), .B(KEYINPUT39), .ZN(n638) );
  NAND2_X1 U703 ( .A1(n758), .A2(n757), .ZN(n621) );
  INV_X1 U704 ( .A(n407), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n660) );
  NAND2_X1 U707 ( .A1(n631), .A2(n627), .ZN(n629) );
  INV_X1 U708 ( .A(n628), .ZN(n632) );
  INV_X1 U709 ( .A(n665), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n633) );
  NOR2_X1 U711 ( .A1(n661), .A2(n658), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n635), .B(KEYINPUT47), .ZN(n636) );
  NOR2_X1 U713 ( .A1(n638), .A2(n665), .ZN(n668) );
  INV_X1 U714 ( .A(n668), .ZN(n640) );
  INV_X1 U715 ( .A(n641), .ZN(n642) );
  XNOR2_X1 U716 ( .A(KEYINPUT85), .B(KEYINPUT59), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n644), .B(n643), .ZN(n645) );
  INV_X1 U718 ( .A(G952), .ZN(n646) );
  AND2_X1 U719 ( .A1(n646), .A2(G953), .ZN(n723) );
  INV_X1 U720 ( .A(KEYINPUT60), .ZN(n647) );
  NOR2_X1 U721 ( .A1(n662), .A2(n652), .ZN(n651) );
  XNOR2_X1 U722 ( .A(G104), .B(KEYINPUT111), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n651), .B(n650), .ZN(G6) );
  NOR2_X1 U724 ( .A1(n665), .A2(n652), .ZN(n657) );
  XOR2_X1 U725 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n654) );
  XNOR2_X1 U726 ( .A(G107), .B(KEYINPUT112), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U728 ( .A(KEYINPUT26), .B(n655), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n657), .B(n656), .ZN(G9) );
  XNOR2_X1 U730 ( .A(G128), .B(n658), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n659), .B(KEYINPUT29), .ZN(G30) );
  XOR2_X1 U732 ( .A(G143), .B(n660), .Z(G45) );
  XOR2_X1 U733 ( .A(G146), .B(n661), .Z(G48) );
  NOR2_X1 U734 ( .A1(n662), .A2(n664), .ZN(n663) );
  XOR2_X1 U735 ( .A(G113), .B(n663), .Z(G15) );
  NOR2_X1 U736 ( .A1(n665), .A2(n664), .ZN(n667) );
  XNOR2_X1 U737 ( .A(G116), .B(KEYINPUT115), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n667), .B(n666), .ZN(G18) );
  XOR2_X1 U739 ( .A(G134), .B(n668), .Z(G36) );
  NAND2_X1 U740 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U741 ( .A(KEYINPUT50), .B(n672), .ZN(n679) );
  NOR2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U743 ( .A(KEYINPUT49), .B(n675), .Z(n676) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U747 ( .A(KEYINPUT51), .B(n682), .Z(n683) );
  NAND2_X1 U748 ( .A1(n701), .A2(n683), .ZN(n696) );
  NOR2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n391), .A2(n690), .ZN(n691) );
  NOR2_X1 U752 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U753 ( .A1(n703), .A2(n693), .ZN(n694) );
  XOR2_X1 U754 ( .A(KEYINPUT116), .B(n694), .Z(n695) );
  NAND2_X1 U755 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U756 ( .A(n697), .B(KEYINPUT117), .ZN(n698) );
  XNOR2_X1 U757 ( .A(n698), .B(KEYINPUT52), .ZN(n699) );
  NOR2_X1 U758 ( .A1(n700), .A2(n699), .ZN(n705) );
  INV_X1 U759 ( .A(n701), .ZN(n702) );
  NOR2_X1 U760 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U761 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U762 ( .A(n706), .B(KEYINPUT118), .ZN(n707) );
  NAND2_X1 U763 ( .A1(n707), .A2(n747), .ZN(n708) );
  NOR2_X1 U764 ( .A1(n669), .A2(n708), .ZN(n709) );
  XNOR2_X1 U765 ( .A(n709), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U766 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n711) );
  XNOR2_X1 U767 ( .A(n711), .B(KEYINPUT55), .ZN(n712) );
  XNOR2_X1 U768 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U769 ( .A1(n719), .A2(G478), .ZN(n716) );
  XNOR2_X1 U770 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U771 ( .A1(n723), .A2(n718), .ZN(G63) );
  NAND2_X1 U772 ( .A1(n719), .A2(G217), .ZN(n721) );
  XNOR2_X1 U773 ( .A(n720), .B(n721), .ZN(n722) );
  NOR2_X1 U774 ( .A1(n723), .A2(n722), .ZN(G66) );
  XNOR2_X1 U775 ( .A(G101), .B(KEYINPUT122), .ZN(n725) );
  XNOR2_X1 U776 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U777 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U778 ( .A1(n730), .A2(n729), .ZN(n739) );
  NOR2_X1 U779 ( .A1(n731), .A2(G953), .ZN(n737) );
  NAND2_X1 U780 ( .A1(G224), .A2(G953), .ZN(n732) );
  XNOR2_X1 U781 ( .A(n732), .B(KEYINPUT61), .ZN(n733) );
  XNOR2_X1 U782 ( .A(KEYINPUT120), .B(n733), .ZN(n734) );
  NAND2_X1 U783 ( .A1(n734), .A2(G898), .ZN(n735) );
  XNOR2_X1 U784 ( .A(n735), .B(KEYINPUT121), .ZN(n736) );
  NOR2_X1 U785 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U786 ( .A(n739), .B(n738), .ZN(G69) );
  XOR2_X1 U787 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n743) );
  XNOR2_X1 U788 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U789 ( .A(n743), .B(n742), .ZN(n744) );
  XOR2_X1 U790 ( .A(n745), .B(n744), .Z(n749) );
  XNOR2_X1 U791 ( .A(n746), .B(n749), .ZN(n748) );
  NAND2_X1 U792 ( .A1(n748), .A2(n747), .ZN(n753) );
  XNOR2_X1 U793 ( .A(G227), .B(n749), .ZN(n750) );
  NAND2_X1 U794 ( .A1(n750), .A2(G900), .ZN(n751) );
  NAND2_X1 U795 ( .A1(n751), .A2(G953), .ZN(n752) );
  NAND2_X1 U796 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U797 ( .A(KEYINPUT125), .B(n754), .Z(G72) );
  XNOR2_X1 U798 ( .A(G125), .B(KEYINPUT37), .ZN(n756) );
  XNOR2_X1 U799 ( .A(n756), .B(n755), .ZN(G27) );
  XNOR2_X1 U800 ( .A(n757), .B(G131), .ZN(G33) );
  XNOR2_X1 U801 ( .A(n758), .B(G137), .ZN(G39) );
  XNOR2_X1 U802 ( .A(G101), .B(n759), .ZN(G3) );
endmodule

