//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  NOR2_X1   g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT93), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n211), .A2(KEYINPUT15), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(KEYINPUT15), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT92), .B(G29gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n214), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  OAI22_X1  g017(.A1(new_n210), .A2(new_n216), .B1(new_n218), .B2(new_n213), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT94), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(KEYINPUT94), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G8gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(G1gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n223), .B1(new_n226), .B2(KEYINPUT95), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(G1gat), .B2(new_n224), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n222), .B(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT96), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT99), .ZN(new_n236));
  INV_X1    g035(.A(new_n222), .ZN(new_n237));
  INV_X1    g036(.A(new_n229), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n219), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n242), .B1(new_n222), .B2(new_n240), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n239), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(KEYINPUT18), .A3(new_n232), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n236), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT97), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n206), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT18), .B1(new_n244), .B2(new_n232), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n250), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G226gat), .A2(G233gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT79), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT27), .B(G183gat), .ZN(new_n257));
  INV_X1    g056(.A(G190gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT28), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  INV_X1    g060(.A(G176gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT26), .ZN(new_n264));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n266), .B(new_n267), .C1(new_n264), .C2(new_n263), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT23), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n265), .B1(new_n263), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n272));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n272), .B1(new_n273), .B2(KEYINPUT23), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n263), .A2(KEYINPUT67), .A3(new_n270), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277));
  AND2_X1   g076(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(G190gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n276), .B(KEYINPUT25), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT24), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n267), .A2(KEYINPUT65), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT65), .B1(new_n267), .B2(new_n283), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n279), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT66), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n279), .B(KEYINPUT66), .C1(new_n284), .C2(new_n285), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n289), .A3(new_n276), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n290), .A2(KEYINPUT68), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT68), .B1(new_n290), .B2(new_n291), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n282), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT69), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n296), .B(new_n282), .C1(new_n292), .C2(new_n293), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n269), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n256), .B1(new_n298), .B2(KEYINPUT29), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT80), .B(new_n256), .C1(new_n298), .C2(KEYINPUT29), .ZN(new_n302));
  INV_X1    g101(.A(new_n269), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(new_n255), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G197gat), .B(G204gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT22), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n311), .A2(KEYINPUT78), .B1(G211gat), .B2(G218gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(KEYINPUT78), .B2(new_n311), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n307), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n255), .B1(new_n304), .B2(KEYINPUT29), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n314), .B(new_n315), .Z(new_n319));
  OAI211_X1 g118(.A(new_n318), .B(new_n319), .C1(new_n298), .C2(new_n256), .ZN(new_n320));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G64gat), .B(G92gat), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n321), .B(new_n322), .Z(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n323), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n305), .B1(new_n299), .B2(new_n300), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n319), .B1(new_n326), .B2(new_n302), .ZN(new_n327));
  INV_X1    g126(.A(new_n320), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n325), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n329), .A3(KEYINPUT30), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT30), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n317), .A2(new_n331), .A3(new_n320), .A4(new_n323), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334));
  INV_X1    g133(.A(G127gat), .ZN(new_n335));
  INV_X1    g134(.A(G134gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(G127gat), .A2(G134gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n334), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G113gat), .B(G120gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n341), .B2(KEYINPUT71), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n341), .A2(KEYINPUT71), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n335), .A2(KEYINPUT70), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n335), .A2(KEYINPUT70), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n338), .B1(new_n347), .B2(G134gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n341), .A2(new_n334), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G141gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G148gat), .ZN(new_n353));
  INV_X1    g152(.A(G148gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G141gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT2), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G155gat), .B(G162gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT82), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n353), .A2(new_n355), .B1(KEYINPUT2), .B2(new_n357), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT82), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n364), .A3(new_n360), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n359), .A2(new_n367), .A3(new_n361), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT81), .B1(new_n363), .B2(new_n360), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT4), .B1(new_n351), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(KEYINPUT83), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n362), .A2(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n342), .A2(new_n343), .B1(new_n348), .B2(new_n349), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n373), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n372), .B1(new_n378), .B2(KEYINPUT4), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT5), .ZN(new_n380));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n377), .B1(new_n371), .B2(KEYINPUT3), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n374), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n382), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n379), .A2(new_n380), .A3(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n373), .A2(new_n376), .A3(KEYINPUT4), .A4(new_n377), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n389), .B1(new_n351), .B2(new_n371), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT84), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n386), .A2(KEYINPUT84), .A3(new_n388), .A4(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n374), .B(new_n377), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n380), .B1(new_n396), .B2(new_n382), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n387), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(G57gat), .B(G85gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  AOI21_X1  g201(.A(KEYINPUT6), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n402), .ZN(new_n404));
  INV_X1    g203(.A(new_n397), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n393), .B2(new_n394), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(new_n406), .B2(new_n387), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT6), .B(new_n404), .C1(new_n406), .C2(new_n387), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n333), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT29), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n319), .B1(new_n413), .B2(new_n385), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n384), .B1(new_n316), .B2(KEYINPUT29), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n373), .A2(new_n376), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n415), .A2(new_n371), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n421), .A2(new_n418), .A3(new_n414), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n412), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT31), .B(G50gat), .ZN(new_n425));
  XOR2_X1   g224(.A(new_n424), .B(new_n425), .Z(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G22gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n420), .A2(new_n422), .ZN(new_n429));
  INV_X1    g228(.A(G22gat), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(new_n430), .A3(new_n426), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n428), .A2(KEYINPUT85), .A3(new_n429), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(KEYINPUT85), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n423), .A2(new_n430), .A3(new_n426), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n423), .B2(new_n426), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n411), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT76), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n295), .A2(new_n297), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT72), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n377), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n303), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n377), .B(KEYINPUT72), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n444), .B(new_n445), .C1(new_n298), .C2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT74), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT34), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(KEYINPUT75), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT75), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n447), .B2(new_n448), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n450), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n439), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT32), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n444), .B1(new_n298), .B2(new_n446), .ZN(new_n459));
  INV_X1    g258(.A(new_n445), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n298), .A2(new_n446), .ZN(new_n463));
  AOI211_X1 g262(.A(new_n269), .B(new_n442), .C1(new_n295), .C2(new_n297), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(G71gat), .B(G99gat), .Z(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G43gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n462), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(KEYINPUT33), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(KEYINPUT32), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT73), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT73), .B1(new_n461), .B2(new_n472), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n455), .A2(new_n450), .B1(new_n452), .B2(new_n447), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n449), .A2(KEYINPUT75), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT34), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT76), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n457), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n473), .A2(new_n474), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n461), .A2(KEYINPUT73), .A3(new_n472), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n485), .A2(new_n471), .A3(new_n480), .A4(new_n478), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(KEYINPUT36), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n478), .A2(new_n480), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n477), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n485), .A2(new_n471), .B1(new_n478), .B2(new_n480), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n407), .A2(KEYINPUT87), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(new_n404), .C1(new_n406), .C2(new_n387), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n403), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n324), .A2(new_n409), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT88), .B(KEYINPUT38), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n323), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n320), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n327), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n316), .B1(new_n326), .B2(new_n302), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n318), .B1(new_n298), .B2(new_n256), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT37), .B1(new_n505), .B2(new_n319), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT89), .B1(new_n498), .B2(new_n508), .ZN(new_n509));
  OAI221_X1 g308(.A(new_n500), .B1(new_n327), .B2(new_n502), .C1(new_n504), .C2(new_n506), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n497), .A2(new_n409), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .A4(new_n324), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n501), .B1(new_n317), .B2(new_n320), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n325), .B1(new_n327), .B2(new_n502), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n499), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n509), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT39), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n396), .A2(new_n382), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(KEYINPUT86), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n383), .A2(new_n385), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n379), .A2(new_n521), .ZN(new_n522));
  OAI221_X1 g321(.A(new_n520), .B1(KEYINPUT86), .B2(new_n519), .C1(new_n522), .C2(new_n381), .ZN(new_n523));
  OR3_X1    g322(.A1(new_n522), .A2(KEYINPUT39), .A3(new_n381), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n402), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT40), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n494), .A2(new_n496), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n525), .A2(new_n526), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n330), .A2(new_n332), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n437), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n438), .B(new_n493), .C1(new_n517), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n482), .A2(new_n532), .A3(new_n486), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT35), .B1(new_n535), .B2(new_n411), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT90), .B1(new_n490), .B2(new_n491), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n437), .B1(new_n332), .B2(new_n330), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n477), .A2(new_n489), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT90), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n486), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT91), .B(KEYINPUT35), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n512), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n537), .A2(new_n538), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n254), .B1(new_n534), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT41), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT101), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(G85gat), .A3(G92gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553));
  INV_X1    g352(.A(G85gat), .ZN(new_n554));
  INV_X1    g353(.A(G92gat), .ZN(new_n555));
  AOI22_X1  g354(.A1(KEYINPUT8), .A2(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n549), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n552), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G99gat), .B(G106gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n548), .B1(new_n237), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n243), .B2(new_n560), .ZN(new_n562));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n547), .A2(KEYINPUT41), .ZN(new_n565));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n568), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G57gat), .B(G64gat), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT100), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G71gat), .B(G78gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(new_n335), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n238), .B1(new_n577), .B2(new_n576), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G155gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n571), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n593));
  OR3_X1    g392(.A1(new_n560), .A2(new_n576), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n560), .B(new_n576), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n594), .B1(new_n595), .B2(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT102), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n595), .A2(G230gat), .A3(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n597), .B(KEYINPUT103), .Z(new_n607));
  AND2_X1   g406(.A1(new_n596), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n604), .B1(new_n608), .B2(new_n600), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n592), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n546), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n410), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G1gat), .ZN(G1324gat));
  INV_X1    g416(.A(new_n333), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n223), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT105), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n225), .A2(new_n223), .ZN(new_n621));
  NAND2_X1  g420(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n614), .A2(new_n618), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT104), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT42), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT42), .B1(new_n623), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n620), .B1(new_n625), .B2(new_n626), .ZN(G1325gat));
  INV_X1    g426(.A(new_n614), .ZN(new_n628));
  OAI21_X1  g427(.A(G15gat), .B1(new_n628), .B2(new_n493), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n537), .A2(new_n541), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n630), .A2(G15gat), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n628), .B2(new_n631), .ZN(G1326gat));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n437), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT43), .B(G22gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(G1327gat));
  NOR2_X1   g434(.A1(new_n590), .A2(new_n610), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n571), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n546), .A2(new_n615), .A3(new_n215), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT45), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n411), .A2(KEYINPUT106), .A3(new_n437), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n615), .B1(new_n330), .B2(new_n332), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(new_n532), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n509), .A2(new_n513), .A3(new_n516), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n531), .A2(new_n532), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n646), .A2(new_n647), .B1(new_n492), .B2(new_n487), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n645), .A2(new_n648), .B1(new_n536), .B2(new_n544), .ZN(new_n649));
  INV_X1    g448(.A(new_n571), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n640), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n534), .A2(new_n545), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n650), .A2(new_n640), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n651), .A2(new_n253), .A3(new_n654), .A4(new_n636), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n410), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n639), .B1(new_n656), .B2(new_n215), .ZN(G1328gat));
  NAND2_X1  g456(.A1(new_n546), .A2(new_n637), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n658), .A2(G36gat), .A3(new_n333), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT46), .ZN(new_n660));
  OAI21_X1  g459(.A(G36gat), .B1(new_n655), .B2(new_n333), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(G1329gat));
  NAND3_X1  g461(.A1(new_n487), .A2(new_n492), .A3(G43gat), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n658), .A2(new_n630), .ZN(new_n664));
  OAI22_X1  g463(.A1(new_n655), .A2(new_n663), .B1(G43gat), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g465(.A1(new_n658), .A2(G50gat), .A3(new_n532), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n655), .A2(new_n532), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n668), .B2(G50gat), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1331gat));
  NAND3_X1  g470(.A1(new_n254), .A2(new_n610), .A3(new_n592), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT108), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n646), .A2(new_n647), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n674), .A2(new_n493), .A3(new_n644), .A4(new_n641), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n545), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n615), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g479(.A1(new_n677), .A2(new_n333), .ZN(new_n681));
  NOR2_X1   g480(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n682));
  AND2_X1   g481(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n681), .B2(new_n682), .ZN(G1333gat));
  OAI21_X1  g484(.A(G71gat), .B1(new_n677), .B2(new_n493), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n630), .A2(G71gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n677), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g488(.A1(new_n678), .A2(new_n437), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g490(.A1(new_n253), .A2(new_n611), .A3(new_n590), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n650), .B1(new_n675), .B2(new_n545), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n654), .B(new_n692), .C1(new_n693), .C2(KEYINPUT44), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT109), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n651), .A2(new_n696), .A3(new_n654), .A4(new_n692), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G85gat), .B1(new_n698), .B2(new_n410), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n649), .B2(new_n650), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n253), .A2(new_n590), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n676), .A2(KEYINPUT110), .A3(new_n571), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT51), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n701), .A2(new_n703), .A3(KEYINPUT51), .A4(new_n702), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n410), .A2(G85gat), .A3(new_n611), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT111), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n699), .B1(new_n708), .B2(new_n710), .ZN(G1336gat));
  AOI21_X1  g510(.A(KEYINPUT51), .B1(new_n704), .B2(KEYINPUT114), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT114), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n701), .A2(new_n703), .A3(new_n713), .A4(new_n702), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n712), .A2(KEYINPUT115), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT115), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n707), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n712), .B2(new_n714), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n333), .A2(G92gat), .A3(new_n611), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT113), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n715), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n695), .A2(new_n618), .A3(new_n697), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G92gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT112), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n722), .A2(new_n725), .A3(G92gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT52), .B1(new_n721), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G92gat), .B1(new_n694), .B2(new_n333), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n706), .A2(new_n707), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(new_n719), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT116), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n728), .A2(new_n735), .ZN(G1337gat));
  OAI21_X1  g535(.A(G99gat), .B1(new_n698), .B2(new_n493), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n630), .A2(G99gat), .A3(new_n611), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n708), .B2(new_n738), .ZN(G1338gat));
  NOR3_X1   g538(.A1(new_n532), .A2(G106gat), .A3(new_n611), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n732), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT53), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT117), .B(G106gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n694), .A2(new_n532), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n698), .A2(new_n532), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n743), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n715), .A2(new_n718), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n740), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n745), .B1(new_n749), .B2(new_n742), .ZN(G1339gat));
  OAI211_X1 g549(.A(new_n599), .B(KEYINPUT54), .C1(new_n596), .C2(new_n607), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n603), .B1(new_n608), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n754), .A2(KEYINPUT55), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(KEYINPUT55), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n606), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n253), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n206), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n244), .A2(new_n232), .B1(new_n230), .B2(new_n234), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n250), .A2(new_n760), .B1(new_n205), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n610), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n571), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n758), .A2(new_n571), .A3(new_n762), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n591), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n254), .A2(new_n611), .A3(new_n592), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n630), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n768), .A2(new_n615), .A3(new_n769), .A4(new_n538), .ZN(new_n770));
  INV_X1    g569(.A(G113gat), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n770), .A2(new_n771), .A3(new_n254), .ZN(new_n772));
  INV_X1    g571(.A(new_n768), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n773), .A2(new_n410), .A3(new_n535), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(new_n333), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n253), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n772), .B1(new_n776), .B2(new_n771), .ZN(G1340gat));
  INV_X1    g576(.A(G120gat), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n770), .A2(new_n778), .A3(new_n611), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n775), .A2(new_n610), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(new_n778), .ZN(G1341gat));
  NAND4_X1  g580(.A1(new_n775), .A2(new_n346), .A3(new_n345), .A4(new_n590), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n347), .B1(new_n770), .B2(new_n591), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1342gat));
  NOR2_X1   g583(.A1(new_n618), .A2(new_n650), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n774), .A2(new_n336), .A3(new_n785), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n786), .A2(KEYINPUT56), .ZN(new_n787));
  OAI21_X1  g586(.A(G134gat), .B1(new_n770), .B2(new_n650), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(KEYINPUT56), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(G1343gat));
  AOI21_X1  g589(.A(new_n532), .B1(new_n766), .B2(new_n767), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n757), .A2(KEYINPUT118), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n757), .A2(KEYINPUT118), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n253), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n571), .B1(new_n796), .B2(new_n763), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n591), .B1(new_n797), .B2(new_n765), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n532), .B1(new_n798), .B2(new_n767), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n793), .B1(new_n799), .B2(new_n792), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n410), .B1(new_n487), .B2(new_n492), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n333), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n800), .A2(new_n254), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n802), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n791), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n253), .A2(new_n352), .ZN(new_n806));
  OAI22_X1  g605(.A1(new_n803), .A2(new_n352), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g607(.A(new_n805), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n354), .A3(new_n610), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n437), .A2(new_n792), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n767), .B(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n798), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n791), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n816), .B2(KEYINPUT57), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n610), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n804), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n811), .B1(new_n819), .B2(G148gat), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n800), .A2(new_n802), .ZN(new_n821));
  AOI211_X1 g620(.A(KEYINPUT59), .B(new_n354), .C1(new_n821), .C2(new_n610), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n810), .B1(new_n820), .B2(new_n822), .ZN(G1345gat));
  INV_X1    g622(.A(G155gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n824), .A3(new_n590), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n800), .A2(new_n591), .A3(new_n802), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n824), .ZN(G1346gat));
  NOR3_X1   g626(.A1(new_n800), .A2(new_n650), .A3(new_n802), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(KEYINPUT120), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(KEYINPUT120), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(G162gat), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(G162gat), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n791), .A2(new_n832), .A3(new_n785), .A4(new_n801), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1347gat));
  NOR4_X1   g633(.A1(new_n773), .A2(new_n615), .A3(new_n333), .A4(new_n535), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n261), .A3(new_n253), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n773), .A2(new_n437), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n333), .A2(new_n615), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n769), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n839), .A2(KEYINPUT121), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(KEYINPUT121), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G169gat), .B1(new_n842), .B2(new_n254), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(KEYINPUT122), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(KEYINPUT122), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n836), .B1(new_n844), .B2(new_n845), .ZN(G1348gat));
  OAI21_X1  g645(.A(G176gat), .B1(new_n842), .B2(new_n611), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n835), .A2(new_n262), .A3(new_n610), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1349gat));
  OAI21_X1  g648(.A(G183gat), .B1(new_n842), .B2(new_n591), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n257), .A3(new_n590), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g651(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n853));
  XNOR2_X1  g652(.A(new_n852), .B(new_n853), .ZN(G1350gat));
  NOR2_X1   g653(.A1(new_n842), .A2(new_n650), .ZN(new_n855));
  NAND2_X1  g654(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G190gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  OR3_X1    g657(.A1(new_n858), .A2(KEYINPUT125), .A3(KEYINPUT61), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n835), .A2(new_n258), .A3(new_n571), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT124), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(G1351gat));
  NAND2_X1  g662(.A1(new_n493), .A2(new_n838), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n816), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(G197gat), .B1(new_n865), .B2(new_n253), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n864), .B(KEYINPUT126), .Z(new_n867));
  AND2_X1   g666(.A1(new_n817), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n253), .A2(G197gat), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(G1352gat));
  INV_X1    g669(.A(new_n865), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(G204gat), .A3(new_n611), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT62), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n818), .A2(new_n867), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G204gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1353gat));
  OR3_X1    g675(.A1(new_n871), .A2(G211gat), .A3(new_n591), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n868), .A2(new_n590), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n878), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT63), .B1(new_n878), .B2(G211gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(G1354gat));
  INV_X1    g680(.A(G218gat), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n882), .B1(new_n868), .B2(new_n571), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT127), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n871), .A2(G218gat), .A3(new_n650), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n884), .B1(new_n883), .B2(new_n885), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1355gat));
endmodule


