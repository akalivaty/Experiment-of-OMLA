//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n203), .A2(G183gat), .A3(G190gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(G183gat), .B(G190gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(new_n203), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NOR3_X1   g013(.A1(new_n210), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n208), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n206), .A2(new_n207), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT25), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n206), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n206), .A2(new_n219), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n215), .A4(new_n222), .ZN(new_n223));
  OR3_X1    g022(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(KEYINPUT69), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n212), .A2(new_n213), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(new_n214), .B2(KEYINPUT26), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(KEYINPUT69), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G183gat), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n230), .A2(KEYINPUT27), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(KEYINPUT27), .ZN(new_n232));
  INV_X1    g031(.A(G190gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n234), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236));
  AOI211_X1 g035(.A(KEYINPUT28), .B(G190gat), .C1(new_n232), .C2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(new_n236), .B2(new_n232), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n231), .B(KEYINPUT68), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n229), .B(new_n235), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n218), .A2(new_n223), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT72), .ZN(new_n242));
  INV_X1    g041(.A(G127gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G134gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT71), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G134gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G127gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT70), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(new_n247), .A3(G127gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n242), .B1(new_n246), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n244), .B(KEYINPUT71), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n254), .A2(KEYINPUT72), .A3(new_n249), .A4(new_n251), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(G113gat), .B(G120gat), .Z(new_n257));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT73), .B(KEYINPUT1), .Z(new_n261));
  NAND4_X1  g060(.A1(new_n257), .A2(new_n261), .A3(new_n244), .A4(new_n248), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT74), .B1(new_n241), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n223), .A2(new_n240), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT74), .ZN(new_n266));
  INV_X1    g065(.A(new_n262), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n256), .B2(new_n259), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n265), .A2(new_n266), .A3(new_n268), .A4(new_n218), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n241), .A2(new_n263), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n264), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n202), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT33), .B1(new_n271), .B2(new_n273), .ZN(new_n275));
  XNOR2_X1  g074(.A(G15gat), .B(G43gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(G71gat), .B(G99gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n274), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n271), .A2(new_n273), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT32), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n278), .A2(KEYINPUT75), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n278), .A2(KEYINPUT75), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT33), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n264), .A2(new_n269), .A3(new_n272), .A4(new_n270), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT34), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n279), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT34), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n287), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n280), .A2(new_n284), .ZN(new_n292));
  INV_X1    g091(.A(new_n278), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n281), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n285), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n274), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n291), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G78gat), .B(G106gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT31), .B(G50gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n301), .A2(KEYINPUT81), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n302), .B(KEYINPUT82), .Z(new_n303));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT76), .B(G218gat), .Z(new_n305));
  INV_X1    g104(.A(G211gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G197gat), .B(G204gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT3), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(G155gat), .B(G162gat), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G155gat), .ZN(new_n319));
  INV_X1    g118(.A(G162gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT2), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G141gat), .B(G148gat), .Z(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n321), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n317), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n323), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n329), .A2(new_n315), .ZN(new_n330));
  OAI22_X1  g129(.A1(new_n316), .A2(new_n327), .B1(new_n314), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G228gat), .A2(G233gat), .ZN(new_n332));
  INV_X1    g131(.A(G22gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n331), .A2(new_n335), .B1(KEYINPUT81), .B2(new_n301), .ZN(new_n336));
  OAI221_X1 g135(.A(new_n334), .B1(new_n314), .B2(new_n330), .C1(new_n316), .C2(new_n327), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n303), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n314), .A2(new_n315), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n327), .B1(new_n339), .B2(new_n328), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n330), .A2(new_n314), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n335), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n301), .A2(KEYINPUT81), .ZN(new_n343));
  AND4_X1   g142(.A1(new_n337), .A2(new_n342), .A3(new_n343), .A4(new_n303), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n289), .A2(new_n297), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT35), .ZN(new_n347));
  XOR2_X1   g146(.A(G1gat), .B(G29gat), .Z(new_n348));
  XNOR2_X1  g147(.A(G57gat), .B(G85gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n326), .A2(KEYINPUT3), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n253), .A2(new_n255), .B1(new_n258), .B2(new_n257), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n329), .B(new_n353), .C1(new_n354), .C2(new_n267), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n260), .A2(new_n262), .A3(new_n327), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT4), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n354), .A2(new_n267), .A3(new_n326), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n327), .B1(new_n260), .B2(new_n262), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(new_n358), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n361), .A2(new_n362), .B1(KEYINPUT5), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n367), .B(new_n363), .C1(new_n357), .C2(new_n360), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n352), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(KEYINPUT5), .ZN(new_n370));
  NOR4_X1   g169(.A1(new_n354), .A2(KEYINPUT4), .A3(new_n267), .A4(new_n326), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n359), .B1(new_n268), .B2(new_n327), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(new_n355), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(new_n363), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n352), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n361), .A2(KEYINPUT5), .A3(new_n362), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n369), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT6), .A4(new_n375), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n241), .A2(new_n315), .ZN(new_n382));
  NAND2_X1  g181(.A1(G226gat), .A2(G233gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT77), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n384), .B(KEYINPUT78), .Z(new_n387));
  NAND2_X1  g186(.A1(new_n241), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n314), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n314), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n385), .B1(new_n265), .B2(new_n218), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n387), .B1(new_n241), .B2(new_n315), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n394), .B(new_n395), .Z(new_n396));
  NAND3_X1  g195(.A1(new_n389), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n389), .A2(new_n393), .A3(KEYINPUT30), .A4(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n389), .A2(new_n393), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n396), .B(KEYINPUT79), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n399), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n346), .A2(new_n347), .A3(new_n381), .A4(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n288), .B1(new_n279), .B2(new_n286), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n294), .A2(new_n296), .A3(new_n291), .ZN(new_n407));
  INV_X1    g206(.A(new_n345), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n406), .A2(new_n404), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n381), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT35), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n338), .B2(new_n344), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n342), .A2(new_n337), .A3(new_n343), .ZN(new_n415));
  INV_X1    g214(.A(new_n303), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n336), .A2(new_n337), .A3(new_n303), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT83), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n381), .B2(new_n404), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT36), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n289), .B2(new_n297), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n406), .A2(KEYINPUT36), .A3(new_n407), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT39), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n357), .A2(new_n426), .A3(new_n360), .A4(new_n363), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n352), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(KEYINPUT84), .A3(new_n352), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n373), .A2(new_n363), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n364), .A2(new_n358), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n426), .B1(new_n433), .B2(new_n362), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n430), .A2(new_n431), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT85), .B1(new_n435), .B2(KEYINPUT40), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n434), .ZN(new_n437));
  INV_X1    g236(.A(new_n431), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT84), .B1(new_n427), .B2(new_n352), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT40), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n366), .A2(new_n368), .A3(new_n352), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n397), .A2(new_n398), .B1(new_n401), .B2(new_n402), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n400), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n435), .A2(KEYINPUT40), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n436), .A2(new_n443), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n386), .A2(new_n390), .A3(new_n388), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n314), .B1(new_n391), .B2(new_n392), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT37), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT38), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n402), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n451), .B(new_n453), .C1(new_n401), .C2(KEYINPUT37), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n454), .A2(new_n397), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n401), .A2(KEYINPUT37), .ZN(new_n456));
  INV_X1    g255(.A(new_n396), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n401), .B2(KEYINPUT37), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT38), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n455), .A2(new_n459), .A3(new_n380), .A4(new_n379), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n448), .A2(new_n408), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n425), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n412), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G57gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G64gat), .ZN(new_n465));
  INV_X1    g264(.A(G64gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(G57gat), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT9), .ZN(new_n468));
  NAND2_X1  g267(.A1(G71gat), .A2(G78gat), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n465), .A2(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n469), .ZN(new_n471));
  NOR2_X1   g270(.A1(G71gat), .A2(G78gat), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G71gat), .ZN(new_n474));
  INV_X1    g273(.A(G78gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT94), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT94), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(G71gat), .B2(G78gat), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n471), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n469), .A2(new_n468), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n466), .A2(G57gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n464), .A2(G64gat), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n479), .A2(new_n483), .A3(KEYINPUT95), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT95), .B1(new_n479), .B2(new_n483), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n473), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT21), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G127gat), .B(G155gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(new_n489), .Z(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT16), .ZN(new_n492));
  AOI21_X1  g291(.A(G1gat), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n333), .A2(G15gat), .ZN(new_n494));
  INV_X1    g293(.A(G15gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G22gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT90), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G8gat), .ZN(new_n498));
  INV_X1    g297(.A(G8gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n491), .A2(KEYINPUT90), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n493), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n493), .B1(new_n498), .B2(new_n500), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n486), .A2(KEYINPUT97), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT95), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n477), .A2(G71gat), .A3(G78gat), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT94), .B1(new_n474), .B2(new_n475), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n469), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n506), .B1(new_n509), .B2(new_n470), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n479), .A2(new_n483), .A3(KEYINPUT95), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT97), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n473), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n504), .B1(new_n515), .B2(new_n487), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n490), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n488), .A2(new_n489), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n488), .A2(new_n489), .ZN(new_n519));
  OAI221_X1 g318(.A(new_n504), .B1(new_n515), .B2(new_n487), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G231gat), .A2(G233gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT96), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G183gat), .B(G211gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n517), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n526), .B1(new_n517), .B2(new_n520), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT88), .ZN(new_n530));
  NOR2_X1   g329(.A1(G29gat), .A2(G36gat), .ZN(new_n531));
  OR2_X1    g330(.A1(KEYINPUT86), .A2(KEYINPUT14), .ZN(new_n532));
  NAND2_X1  g331(.A1(KEYINPUT86), .A2(KEYINPUT14), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n533), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n530), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n538));
  INV_X1    g337(.A(G43gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n540));
  INV_X1    g339(.A(G50gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G43gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(G50gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n538), .B(new_n540), .C1(new_n544), .C2(KEYINPUT87), .ZN(new_n545));
  AND2_X1   g344(.A1(KEYINPUT86), .A2(KEYINPUT14), .ZN(new_n546));
  NOR2_X1   g345(.A1(KEYINPUT86), .A2(KEYINPUT14), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(KEYINPUT88), .B(new_n535), .C1(new_n548), .C2(new_n531), .ZN(new_n549));
  AND2_X1   g348(.A1(G29gat), .A2(G36gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(G43gat), .B(G50gat), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(KEYINPUT15), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n537), .A2(new_n545), .A3(new_n549), .A4(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n544), .A2(new_n538), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n534), .A2(new_n536), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n555), .B2(new_n550), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT89), .B(KEYINPUT17), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n553), .A2(KEYINPUT17), .A3(new_n556), .ZN(new_n560));
  XOR2_X1   g359(.A(G99gat), .B(G106gat), .Z(new_n561));
  INV_X1    g360(.A(KEYINPUT100), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(G85gat), .A3(G92gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT7), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT7), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n562), .A2(new_n565), .A3(G85gat), .A4(G92gat), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT101), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT101), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(G85gat), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G99gat), .ZN(new_n574));
  INV_X1    g373(.A(G106gat), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT8), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n561), .B1(new_n567), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n561), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n566), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n573), .A4(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n559), .A2(new_n560), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT98), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT41), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n582), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n590), .B2(new_n557), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n583), .A2(new_n585), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT102), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT99), .B(G134gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G162gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n587), .A2(new_n588), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n591), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n584), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n592), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n601), .A2(KEYINPUT102), .A3(new_n592), .A4(new_n598), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT103), .B1(new_n529), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n517), .A2(new_n520), .ZN(new_n608));
  INV_X1    g407(.A(new_n526), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n517), .A2(new_n520), .A3(new_n526), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT103), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n607), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n486), .A2(new_n582), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n512), .A2(new_n581), .A3(new_n578), .A4(new_n473), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n578), .A2(KEYINPUT10), .A3(new_n581), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n505), .A2(new_n514), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n615), .A2(new_n616), .ZN(new_n624));
  INV_X1    g423(.A(new_n622), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT104), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n623), .A2(new_n626), .A3(new_n631), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n606), .A2(new_n614), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n559), .A2(new_n504), .A3(new_n560), .ZN(new_n640));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT91), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n503), .A2(new_n557), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n503), .B2(new_n557), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n640), .B(new_n641), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT92), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT18), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n503), .A2(new_n557), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT91), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n503), .A2(new_n557), .A3(new_n642), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT92), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n651), .A2(new_n652), .A3(new_n641), .A4(new_n640), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n646), .A2(new_n647), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n651), .A2(KEYINPUT18), .A3(new_n641), .A4(new_n640), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n503), .A2(new_n557), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n643), .B2(new_n644), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n641), .B(KEYINPUT13), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n655), .A2(new_n659), .A3(KEYINPUT93), .ZN(new_n662));
  XNOR2_X1  g461(.A(G113gat), .B(G141gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G197gat), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT11), .B(G169gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT12), .Z(new_n667));
  NAND3_X1  g466(.A1(new_n661), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n667), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n654), .B(new_n660), .C1(KEYINPUT93), .C2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n606), .A2(new_n614), .A3(KEYINPUT105), .A4(new_n636), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n639), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n463), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n410), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g476(.A1(new_n674), .A2(new_n404), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n499), .B2(new_n678), .ZN(new_n681));
  MUX2_X1   g480(.A(new_n680), .B(new_n681), .S(KEYINPUT42), .Z(G1325gat));
  AND2_X1   g481(.A1(new_n423), .A2(new_n424), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n675), .A2(G15gat), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n289), .A2(new_n297), .ZN(new_n685));
  AOI21_X1  g484(.A(G15gat), .B1(new_n675), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n420), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n411), .A2(new_n405), .B1(new_n425), .B2(new_n461), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n607), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n463), .A2(KEYINPUT44), .A3(new_n605), .ZN(new_n697));
  INV_X1    g496(.A(new_n671), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(new_n612), .A3(new_n635), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n381), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n695), .A2(new_n607), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n699), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(G29gat), .A3(new_n381), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n705), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n707), .B1(new_n706), .B2(new_n708), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n701), .B1(new_n709), .B2(new_n710), .ZN(G1328gat));
  NOR3_X1   g510(.A1(new_n703), .A2(G36gat), .A3(new_n404), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT46), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n700), .B2(new_n404), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1329gat));
  INV_X1    g514(.A(new_n685), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n539), .B1(new_n703), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n683), .A2(G43gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n700), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g519(.A1(new_n696), .A2(new_n697), .A3(new_n345), .A4(new_n699), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n541), .B1(new_n721), .B2(KEYINPUT108), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(KEYINPUT108), .B2(new_n721), .ZN(new_n723));
  INV_X1    g522(.A(new_n420), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n702), .A2(new_n541), .A3(new_n724), .A4(new_n699), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n723), .A2(KEYINPUT48), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G50gat), .B1(new_n700), .B2(new_n420), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n727), .A2(new_n725), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n728), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g528(.A1(new_n606), .A2(new_n614), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n671), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n635), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT109), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n463), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n381), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n464), .ZN(G1332gat));
  AOI211_X1 g535(.A(new_n404), .B(new_n734), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1333gat));
  OAI21_X1  g538(.A(new_n474), .B1(new_n734), .B2(new_n716), .ZN(new_n740));
  INV_X1    g539(.A(new_n734), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n683), .A2(G71gat), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n741), .A2(KEYINPUT110), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT110), .B1(new_n741), .B2(new_n743), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n740), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g546(.A1(new_n734), .A2(new_n420), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n475), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n698), .A2(new_n529), .ZN(new_n750));
  AOI211_X1 g549(.A(new_n607), .B(new_n750), .C1(new_n412), .C2(new_n462), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT51), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(new_n635), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n569), .A2(new_n571), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n410), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n750), .A2(new_n636), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n696), .A2(new_n697), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT111), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n696), .A2(new_n697), .A3(new_n759), .A4(new_n756), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n758), .A2(new_n410), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n755), .B1(new_n754), .B2(new_n761), .ZN(G1336gat));
  INV_X1    g561(.A(new_n404), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n758), .A2(new_n763), .A3(new_n760), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(G92gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n751), .B2(KEYINPUT112), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n463), .A2(new_n605), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n768), .B(KEYINPUT51), .C1(new_n769), .C2(new_n750), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n404), .A2(G92gat), .A3(new_n636), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n767), .A2(new_n770), .A3(KEYINPUT113), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT52), .B1(new_n765), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(new_n752), .B2(new_n771), .ZN(new_n778));
  OAI21_X1  g577(.A(G92gat), .B1(new_n757), .B2(new_n404), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(G1337gat));
  NAND3_X1  g580(.A1(new_n753), .A2(new_n574), .A3(new_n685), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n758), .A2(new_n683), .A3(new_n760), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n574), .B2(new_n783), .ZN(G1338gat));
  NAND4_X1  g583(.A1(new_n696), .A2(new_n697), .A3(new_n345), .A4(new_n756), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n575), .B1(new_n785), .B2(KEYINPUT115), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(KEYINPUT115), .B2(new_n785), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n345), .A2(new_n575), .A3(new_n635), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT114), .Z(new_n789));
  AOI21_X1  g588(.A(KEYINPUT53), .B1(new_n752), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n758), .A2(new_n724), .A3(new_n760), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n767), .A2(new_n770), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n792), .A2(G106gat), .B1(new_n793), .B2(new_n789), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(G1339gat));
  NOR3_X1   g595(.A1(new_n730), .A2(new_n671), .A3(new_n635), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n618), .A2(new_n620), .A3(new_n625), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n623), .A2(KEYINPUT54), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n625), .B1(new_n618), .B2(new_n620), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n631), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n804), .A2(new_n634), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n800), .A2(new_n803), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g608(.A(KEYINPUT116), .B(KEYINPUT55), .C1(new_n800), .C2(new_n803), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n805), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n654), .A2(new_n660), .A3(new_n669), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n657), .A2(new_n658), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n641), .B1(new_n651), .B2(new_n640), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n666), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n812), .A2(new_n605), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n798), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n812), .A2(new_n605), .A3(new_n816), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n618), .A2(new_n620), .A3(new_n625), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n820), .A2(new_n801), .A3(new_n802), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n621), .A2(new_n802), .A3(new_n622), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n632), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n808), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT116), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT55), .B1(new_n800), .B2(new_n803), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n806), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n819), .A2(new_n828), .A3(KEYINPUT117), .A4(new_n805), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n812), .A2(new_n816), .A3(new_n635), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n804), .A2(new_n634), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n825), .B2(new_n827), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n830), .B1(new_n832), .B2(new_n671), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n818), .B(new_n829), .C1(new_n833), .C2(new_n605), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n797), .B1(new_n834), .B2(new_n529), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(new_n381), .A3(new_n409), .ZN(new_n836));
  AOI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n671), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n671), .ZN(new_n838));
  INV_X1    g637(.A(new_n830), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n605), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n818), .A2(new_n829), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n529), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n797), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n420), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n410), .A2(new_n404), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n845), .A2(new_n716), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n671), .A2(G113gat), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n837), .B1(new_n847), .B2(new_n848), .ZN(G1340gat));
  AOI21_X1  g648(.A(G120gat), .B1(new_n836), .B2(new_n635), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n635), .A2(G120gat), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n847), .B2(new_n851), .ZN(G1341gat));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n612), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n855));
  AOI21_X1  g654(.A(G127gat), .B1(new_n854), .B2(KEYINPUT118), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n529), .A2(new_n243), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n855), .A2(new_n856), .B1(new_n847), .B2(new_n857), .ZN(G1342gat));
  AND2_X1   g657(.A1(new_n847), .A2(new_n605), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(new_n247), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n836), .A2(new_n247), .A3(new_n605), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(KEYINPUT56), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(KEYINPUT56), .B2(new_n861), .ZN(G1343gat));
  AOI211_X1 g662(.A(new_n831), .B(new_n826), .C1(new_n668), .C2(new_n670), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n607), .B1(new_n864), .B2(new_n830), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n818), .A3(new_n829), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n797), .B1(new_n866), .B2(new_n529), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT57), .B1(new_n867), .B2(new_n420), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n408), .B1(new_n842), .B2(new_n843), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n683), .A2(new_n846), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n868), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n873), .B2(new_n698), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n844), .A2(new_n410), .ZN(new_n875));
  NOR4_X1   g674(.A1(new_n875), .A2(new_n763), .A3(new_n408), .A4(new_n683), .ZN(new_n876));
  INV_X1    g675(.A(G141gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n671), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g678(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n880));
  XNOR2_X1  g679(.A(new_n879), .B(new_n880), .ZN(G1344gat));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n882), .B(G148gat), .C1(new_n876), .C2(new_n635), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n873), .B2(new_n636), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n420), .A2(KEYINPUT57), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n832), .A2(new_n819), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n612), .B1(new_n865), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n639), .A2(new_n698), .A3(new_n672), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n869), .B2(new_n870), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n872), .A2(KEYINPUT59), .A3(new_n635), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n884), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n883), .B1(new_n892), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g692(.A(G155gat), .B1(new_n873), .B2(new_n529), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n876), .A2(new_n319), .A3(new_n612), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT120), .ZN(G1346gat));
  NOR3_X1   g696(.A1(new_n873), .A2(new_n320), .A3(new_n607), .ZN(new_n898));
  AOI21_X1  g697(.A(G162gat), .B1(new_n876), .B2(new_n605), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n835), .A2(new_n410), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n346), .A2(new_n763), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT121), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n671), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n763), .A2(new_n381), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n845), .A2(new_n716), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n698), .A2(new_n212), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(G1348gat));
  NAND3_X1  g708(.A1(new_n904), .A2(new_n213), .A3(new_n635), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n907), .A2(new_n635), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n213), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT122), .Z(G1349gat));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n904), .A2(new_n231), .A3(new_n232), .A4(new_n612), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n907), .A2(new_n612), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n914), .B(new_n915), .C1(new_n916), .C2(new_n230), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g717(.A(new_n233), .B1(new_n907), .B2(new_n605), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT61), .Z(new_n920));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n233), .A3(new_n605), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1351gat));
  OAI21_X1  g721(.A(KEYINPUT57), .B1(new_n835), .B2(new_n408), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n923), .A2(KEYINPUT124), .A3(new_n889), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT124), .B1(new_n923), .B2(new_n889), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n683), .A2(new_n906), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n671), .A2(G197gat), .ZN(new_n927));
  NOR4_X1   g726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n683), .A2(new_n404), .A3(new_n408), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n901), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n671), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n928), .A2(new_n931), .ZN(G1352gat));
  XOR2_X1   g731(.A(KEYINPUT125), .B(G204gat), .Z(new_n933));
  NOR2_X1   g732(.A1(new_n636), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n901), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT62), .Z(new_n936));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n924), .A2(new_n925), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n926), .A2(new_n636), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n890), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n923), .A2(KEYINPUT124), .A3(new_n889), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n942), .A2(new_n937), .A3(new_n943), .A4(new_n939), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n933), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n936), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g747(.A(KEYINPUT127), .B(new_n936), .C1(new_n940), .C2(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1353gat));
  NOR3_X1   g749(.A1(new_n890), .A2(new_n529), .A3(new_n926), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(new_n306), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT63), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n930), .A2(new_n306), .A3(new_n612), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1354gat));
  AOI21_X1  g754(.A(G218gat), .B1(new_n930), .B2(new_n605), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n926), .A2(new_n305), .A3(new_n607), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n938), .B2(new_n957), .ZN(G1355gat));
endmodule


