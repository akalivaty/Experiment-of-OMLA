//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT27), .B(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT28), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT28), .B1(new_n208), .B2(new_n209), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NOR3_X1   g015(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n212), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n210), .A2(new_n211), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n221), .A2(new_n213), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n212), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n213), .A3(new_n223), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n227), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n212), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n228), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n231), .B1(new_n228), .B2(new_n236), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n220), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G113gat), .ZN(new_n240));
  INV_X1    g039(.A(G120gat), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT1), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT66), .B(G113gat), .Z(new_n244));
  OAI211_X1 g043(.A(new_n242), .B(new_n243), .C1(new_n244), .C2(new_n241), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n242), .B1(new_n240), .B2(new_n241), .ZN(new_n246));
  INV_X1    g045(.A(new_n243), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n239), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n233), .A2(new_n235), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n233), .A2(new_n235), .ZN(new_n252));
  OAI22_X1  g051(.A1(new_n251), .A2(new_n252), .B1(new_n229), .B2(new_n230), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n231), .A3(new_n236), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n219), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(new_n248), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G227gat), .ZN(new_n258));
  INV_X1    g057(.A(G233gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n250), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n205), .B1(new_n261), .B2(KEYINPUT32), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT33), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n261), .B2(new_n264), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n205), .A2(new_n264), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n261), .A2(KEYINPUT32), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n261), .A2(KEYINPUT68), .A3(KEYINPUT32), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n267), .A2(new_n273), .A3(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n250), .A2(new_n257), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n258), .B2(new_n259), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n276), .A2(new_n277), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G197gat), .B(G204gat), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT72), .B(G218gat), .Z(new_n284));
  INV_X1    g083(.A(G211gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(KEYINPUT71), .B(KEYINPUT22), .Z(new_n287));
  OAI21_X1  g086(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G211gat), .B(G218gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n290), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT2), .ZN(new_n294));
  INV_X1    g093(.A(G141gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(G148gat), .ZN(new_n296));
  INV_X1    g095(.A(G148gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(G141gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n294), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300));
  INV_X1    g099(.A(G155gat), .ZN(new_n301));
  INV_X1    g100(.A(G162gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT74), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(G155gat), .B2(G162gat), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n299), .A2(new_n300), .A3(new_n303), .A4(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n294), .A2(new_n301), .A3(new_n302), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n300), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT75), .B1(new_n295), .B2(G148gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(G141gat), .B2(new_n297), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n295), .A2(KEYINPUT75), .A3(G148gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT29), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n293), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n291), .B2(new_n292), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n306), .A2(new_n312), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n321));
  INV_X1    g120(.A(G228gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(new_n259), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n317), .A2(new_n320), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G78gat), .B(G106gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT31), .B(G50gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G22gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(new_n327), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n316), .B(KEYINPUT82), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n318), .A2(KEYINPUT81), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n314), .B1(new_n318), .B2(KEYINPUT81), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n319), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n324), .B(new_n332), .C1(new_n337), .C2(new_n323), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n323), .B1(new_n333), .B2(new_n336), .ZN(new_n339));
  INV_X1    g138(.A(new_n324), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n331), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n261), .A2(new_n264), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT67), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n346), .A2(new_n262), .B1(new_n271), .B2(new_n272), .ZN(new_n347));
  INV_X1    g146(.A(new_n281), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n342), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n282), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n350), .B1(new_n282), .B2(new_n349), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n319), .A2(new_n256), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n306), .A2(new_n312), .A3(new_n245), .A4(new_n248), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n356), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n361), .ZN(new_n363));
  OAI211_X1 g162(.A(KEYINPUT78), .B(new_n363), .C1(new_n357), .C2(new_n359), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n355), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(new_n358), .B2(KEYINPUT4), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n313), .A2(new_n249), .A3(KEYINPUT76), .A4(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n367), .B(new_n369), .C1(new_n368), .C2(new_n359), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n249), .B1(KEYINPUT3), .B2(new_n319), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n313), .A2(new_n314), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n363), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n370), .A2(new_n373), .A3(KEYINPUT77), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT77), .B1(new_n370), .B2(new_n373), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n365), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT79), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT79), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n365), .B(new_n378), .C1(new_n374), .C2(new_n375), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n358), .B(KEYINPUT4), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n373), .A2(new_n355), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT0), .ZN(new_n386));
  XNOR2_X1  g185(.A(G57gat), .B(G85gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n386), .B(new_n387), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT6), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n354), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n382), .B1(new_n377), .B2(new_n379), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n388), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT80), .A3(KEYINPUT6), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(KEYINPUT6), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n388), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n392), .A2(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n255), .B2(KEYINPUT29), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n239), .A2(G226gat), .A3(G233gat), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n400), .A2(new_n401), .A3(new_n293), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n293), .B1(new_n400), .B2(new_n401), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G8gat), .B(G36gat), .Z(new_n405));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n404), .A2(new_n407), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n407), .B(KEYINPUT73), .Z(new_n412));
  NOR2_X1   g211(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n410), .B1(new_n414), .B2(new_n409), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n202), .B1(new_n353), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n347), .A2(new_n348), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n274), .A2(new_n281), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n342), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR4_X1   g221(.A1(new_n398), .A2(new_n422), .A3(KEYINPUT35), .A4(new_n415), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n390), .A2(new_n391), .A3(new_n397), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT80), .B1(new_n394), .B2(KEYINPUT6), .ZN(new_n425));
  NOR4_X1   g224(.A1(new_n393), .A2(new_n354), .A3(new_n391), .A4(new_n388), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n415), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n421), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(KEYINPUT84), .B(KEYINPUT38), .Z(new_n430));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n407), .B1(new_n404), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT37), .B1(new_n402), .B2(new_n403), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n400), .A2(new_n401), .ZN(new_n435));
  INV_X1    g234(.A(new_n293), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n400), .A2(new_n401), .A3(new_n293), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n431), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n430), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n412), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n408), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(new_n424), .C1(new_n425), .C2(new_n426), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n371), .A2(new_n372), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n381), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n363), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n360), .B2(new_n361), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(new_n449), .A3(new_n363), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n388), .A3(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n453), .B(KEYINPUT40), .Z(new_n454));
  NOR2_X1   g253(.A1(new_n394), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n342), .B1(new_n415), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n445), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT36), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n347), .B2(new_n348), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n282), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n418), .A2(new_n419), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n458), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  OAI22_X1  g263(.A1(new_n417), .A2(new_n423), .B1(new_n429), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G113gat), .B(G141gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(G197gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT11), .B(G169gat), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n467), .B(new_n468), .Z(new_n469));
  XOR2_X1   g268(.A(new_n469), .B(KEYINPUT12), .Z(new_n470));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n471));
  INV_X1    g270(.A(G29gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT14), .ZN(new_n473));
  AND2_X1   g272(.A1(G43gat), .A2(G50gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(G43gat), .A2(G50gat), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT15), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT14), .ZN(new_n477));
  AOI21_X1  g276(.A(G36gat), .B1(new_n477), .B2(G29gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G43gat), .B(G50gat), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n478), .B1(new_n481), .B2(KEYINPUT15), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n473), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n476), .A2(new_n479), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(KEYINPUT15), .A3(new_n478), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT14), .A4(new_n472), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  OR2_X1    g286(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n489));
  AOI21_X1  g288(.A(G50gat), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G43gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(G50gat), .ZN(new_n493));
  INV_X1    g292(.A(G50gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(KEYINPUT87), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n490), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(KEYINPUT87), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n492), .A2(G50gat), .ZN(new_n500));
  AOI21_X1  g299(.A(G43gat), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT88), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT15), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n471), .B1(new_n487), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT15), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n488), .A2(new_n489), .ZN(new_n506));
  OAI22_X1  g305(.A1(new_n506), .A2(G50gat), .B1(new_n501), .B2(KEYINPUT88), .ZN(new_n507));
  INV_X1    g306(.A(new_n502), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n509), .A2(KEYINPUT89), .A3(new_n486), .A4(new_n483), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(G1gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(G1gat), .B2(new_n511), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(G8gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n504), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT90), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n504), .A2(new_n510), .A3(new_n518), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n509), .A2(new_n486), .A3(new_n483), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n515), .B1(new_n522), .B2(KEYINPUT17), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n510), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n520), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(KEYINPUT18), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT18), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n517), .A2(new_n519), .B1(new_n525), .B2(new_n523), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(new_n521), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n521), .B(KEYINPUT13), .Z(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n517), .A2(KEYINPUT91), .A3(new_n519), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n504), .A2(new_n510), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(new_n515), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n534), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n470), .B1(new_n532), .B2(new_n541), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n517), .A2(KEYINPUT91), .A3(new_n519), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT91), .B1(new_n517), .B2(new_n519), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n533), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n527), .A2(KEYINPUT18), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n529), .A3(new_n521), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n470), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n542), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G134gat), .B(G162gat), .Z(new_n553));
  AOI21_X1  g352(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g358(.A1(G85gat), .A2(G92gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n559), .A2(new_n562), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G99gat), .B(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n558), .B1(new_n563), .B2(new_n564), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n571), .A2(new_n568), .A3(new_n562), .A4(new_n566), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n574), .B1(new_n522), .B2(KEYINPUT17), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n525), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n504), .A2(new_n510), .A3(new_n574), .ZN(new_n577));
  NAND3_X1  g376(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT95), .ZN(new_n580));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n555), .A2(new_n556), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n582), .B(new_n583), .C1(new_n579), .C2(new_n581), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n580), .B1(new_n579), .B2(new_n581), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n557), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n579), .A2(new_n581), .ZN(new_n587));
  INV_X1    g386(.A(new_n583), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n585), .ZN(new_n590));
  INV_X1    g389(.A(new_n557), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n589), .A2(new_n590), .A3(new_n591), .A4(new_n582), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n595));
  INV_X1    g394(.A(G57gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(G64gat), .ZN(new_n597));
  INV_X1    g396(.A(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(G57gat), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n595), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT92), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT92), .ZN(new_n605));
  NAND2_X1  g404(.A1(G71gat), .A2(G78gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n600), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n606), .ZN(new_n609));
  XNOR2_X1  g408(.A(G57gat), .B(G64gat), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n609), .B(KEYINPUT92), .C1(new_n610), .C2(new_n595), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT93), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n615), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT94), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n612), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n608), .A2(new_n611), .A3(KEYINPUT94), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n515), .B1(KEYINPUT21), .B2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n620), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n620), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n594), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT97), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n573), .A2(new_n612), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n570), .A2(new_n608), .A3(new_n611), .A4(new_n572), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT10), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n570), .A2(KEYINPUT10), .A3(new_n572), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n622), .B2(new_n623), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n634), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G120gat), .B(G148gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT98), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n635), .A2(new_n633), .A3(new_n636), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n640), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g449(.A(KEYINPUT99), .B(new_n634), .C1(new_n637), .C2(new_n639), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n645), .B1(new_n652), .B2(new_n646), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n653), .A2(KEYINPUT100), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(KEYINPUT100), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n648), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n631), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n465), .A2(new_n552), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n465), .A2(KEYINPUT101), .A3(new_n552), .A4(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n398), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n428), .B1(new_n660), .B2(new_n661), .ZN(new_n666));
  INV_X1    g465(.A(G8gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n662), .ZN(new_n669));
  OAI211_X1 g468(.A(KEYINPUT104), .B(G8gat), .C1(new_n669), .C2(new_n428), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n672), .B2(KEYINPUT42), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n666), .B(new_n673), .C1(new_n672), .C2(new_n671), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n675), .B2(KEYINPUT42), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n666), .B2(new_n671), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n668), .B(new_n670), .C1(new_n676), .C2(new_n678), .ZN(G1325gat));
  OR3_X1    g478(.A1(new_n669), .A2(G15gat), .A3(new_n461), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n669), .B2(new_n463), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(G1326gat));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n683), .B1(new_n662), .B2(new_n342), .ZN(new_n684));
  AOI211_X1 g483(.A(KEYINPUT105), .B(new_n421), .C1(new_n660), .C2(new_n661), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n687), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n684), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(G1327gat));
  AND2_X1   g490(.A1(new_n465), .A2(new_n552), .ZN(new_n692));
  INV_X1    g491(.A(new_n630), .ZN(new_n693));
  INV_X1    g492(.A(new_n656), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n594), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n472), .A3(new_n398), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n464), .B2(new_n429), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n445), .A2(new_n456), .B1(new_n460), .B2(new_n462), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n342), .B1(new_n398), .B2(new_n415), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n705), .A3(KEYINPUT106), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n282), .A2(new_n349), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT85), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n282), .A2(new_n350), .A3(new_n349), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n708), .A2(new_n427), .A3(new_n709), .A4(new_n428), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT35), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n416), .A2(new_n202), .A3(new_n421), .A4(new_n420), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n703), .A2(new_n706), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n701), .B1(new_n713), .B2(new_n594), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n465), .A2(KEYINPUT44), .A3(new_n593), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n552), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n695), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n427), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n700), .A2(new_n720), .ZN(G1328gat));
  NOR3_X1   g520(.A1(new_n697), .A2(G36gat), .A3(new_n428), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  OAI21_X1  g522(.A(G36gat), .B1(new_n719), .B2(new_n428), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1329gat));
  NOR2_X1   g524(.A1(new_n463), .A2(new_n506), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n716), .A2(new_n718), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n692), .A2(new_n420), .A3(new_n696), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n728), .A2(new_n506), .B1(new_n729), .B2(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n729), .A2(KEYINPUT47), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1330gat));
  NAND4_X1  g532(.A1(new_n714), .A2(new_n342), .A3(new_n715), .A4(new_n718), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n499), .A2(new_n500), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n421), .A2(new_n735), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n698), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT108), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1331gat));
  AND3_X1   g540(.A1(new_n704), .A2(new_n705), .A3(KEYINPUT106), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT106), .B1(new_n704), .B2(new_n705), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n742), .A2(new_n743), .B1(new_n417), .B2(new_n423), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n631), .A2(new_n552), .A3(new_n694), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n427), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(new_n596), .ZN(G1332gat));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n428), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  AND2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n749), .B2(new_n750), .ZN(G1333gat));
  INV_X1    g552(.A(G71gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n746), .B2(new_n461), .ZN(new_n755));
  INV_X1    g554(.A(new_n746), .ZN(new_n756));
  INV_X1    g555(.A(new_n463), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(G71gat), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n755), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT50), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n764), .B(new_n755), .C1(new_n760), .C2(new_n761), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1334gat));
  NAND2_X1  g565(.A1(new_n756), .A2(new_n342), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g567(.A1(new_n552), .A2(new_n630), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n694), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n716), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n427), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n703), .A2(new_n706), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n711), .A2(new_n712), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n594), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n770), .B1(new_n776), .B2(KEYINPUT111), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n713), .B2(new_n594), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT51), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n744), .A2(KEYINPUT111), .A3(new_n593), .ZN(new_n781));
  AND4_X1   g580(.A1(KEYINPUT51), .A2(new_n779), .A3(new_n769), .A4(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n398), .A2(new_n563), .A3(new_n656), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n773), .B1(new_n783), .B2(new_n784), .ZN(G1336gat));
  NOR3_X1   g584(.A1(new_n428), .A2(G92gat), .A3(new_n694), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n780), .B2(new_n782), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n714), .A2(new_n415), .A3(new_n715), .A4(new_n771), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G92gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n787), .B(new_n789), .C1(KEYINPUT112), .C2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n789), .B2(KEYINPUT112), .ZN(new_n792));
  INV_X1    g591(.A(new_n786), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n781), .A2(new_n769), .ZN(new_n795));
  INV_X1    g594(.A(new_n779), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n777), .A2(KEYINPUT51), .A3(new_n779), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n789), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n792), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n791), .A2(new_n801), .ZN(G1337gat));
  OAI21_X1  g601(.A(G99gat), .B1(new_n772), .B2(new_n463), .ZN(new_n803));
  OR3_X1    g602(.A1(new_n461), .A2(G99gat), .A3(new_n694), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n783), .B2(new_n804), .ZN(G1338gat));
  NOR3_X1   g604(.A1(new_n421), .A2(new_n694), .A3(G106gat), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT114), .Z(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n797), .B2(new_n798), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n714), .A2(new_n342), .A3(new_n715), .A4(new_n771), .ZN(new_n809));
  XOR2_X1   g608(.A(KEYINPUT113), .B(G106gat), .Z(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT53), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(KEYINPUT53), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n806), .B1(new_n780), .B2(new_n782), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(G1339gat));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n650), .A2(new_n818), .A3(new_n651), .ZN(new_n819));
  INV_X1    g618(.A(new_n638), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n624), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT10), .ZN(new_n822));
  INV_X1    g621(.A(new_n636), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n572), .A2(new_n570), .B1(new_n608), .B2(new_n611), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n821), .A2(new_n825), .A3(new_n633), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n640), .A3(KEYINPUT54), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n819), .A2(new_n644), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n644), .A4(new_n827), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT115), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n827), .A2(KEYINPUT55), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n644), .A4(new_n819), .ZN(new_n833));
  AOI221_X4 g632(.A(new_n647), .B1(new_n817), .B2(new_n828), .C1(new_n830), .C2(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n550), .B1(new_n546), .B2(new_n549), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n469), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n534), .B(new_n540), .C1(new_n543), .C2(new_n544), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n530), .A2(new_n521), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n656), .A3(new_n551), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n593), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n533), .A2(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n841), .B1(new_n845), .B2(new_n550), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n593), .A2(new_n834), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT116), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n593), .A2(new_n834), .A3(new_n846), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n552), .A2(new_n834), .B1(new_n846), .B2(new_n656), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n593), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n848), .A2(new_n693), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n657), .A2(new_n717), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n427), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(new_n428), .A3(new_n421), .A4(new_n420), .ZN(new_n856));
  OAI21_X1  g655(.A(G113gat), .B1(new_n856), .B2(new_n717), .ZN(new_n857));
  INV_X1    g656(.A(new_n353), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n415), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n552), .A2(new_n244), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(G1340gat));
  NOR3_X1   g661(.A1(new_n856), .A2(new_n241), .A3(new_n694), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n855), .A2(new_n656), .A3(new_n859), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n241), .B2(new_n864), .ZN(G1341gat));
  OAI21_X1  g664(.A(G127gat), .B1(new_n856), .B2(new_n693), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n693), .A2(G127gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n860), .B2(new_n867), .ZN(G1342gat));
  OR3_X1    g667(.A1(new_n860), .A2(G134gat), .A3(new_n594), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n870));
  OAI21_X1  g669(.A(G134gat), .B1(new_n856), .B2(new_n594), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G1343gat));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n421), .B1(new_n853), .B2(new_n854), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n463), .A2(new_n398), .A3(new_n428), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(G141gat), .A3(new_n717), .ZN(new_n879));
  XOR2_X1   g678(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n853), .A2(new_n854), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n342), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n647), .B1(new_n830), .B2(new_n833), .ZN(new_n885));
  INV_X1    g684(.A(new_n828), .ZN(new_n886));
  XNOR2_X1  g685(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n552), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n593), .B1(new_n888), .B2(new_n843), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n693), .B1(new_n889), .B2(new_n847), .ZN(new_n890));
  AOI211_X1 g689(.A(new_n884), .B(new_n421), .C1(new_n890), .C2(new_n854), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n552), .B(new_n877), .C1(new_n883), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G141gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n879), .B1(new_n893), .B2(KEYINPUT119), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n895), .A3(G141gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n874), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n879), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n893), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT121), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n892), .A2(new_n895), .A3(G141gat), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n895), .B1(new_n892), .B2(G141gat), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n904), .A2(new_n905), .A3(new_n879), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n903), .B(new_n900), .C1(new_n906), .C2(new_n874), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n902), .A2(new_n907), .ZN(G1344gat));
  INV_X1    g707(.A(new_n878), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n297), .A3(new_n656), .ZN(new_n910));
  XOR2_X1   g709(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n911));
  NAND2_X1  g710(.A1(new_n890), .A2(new_n854), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT57), .B1(new_n912), .B2(new_n342), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT123), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n875), .A2(new_n881), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n656), .B(new_n877), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n911), .B1(new_n916), .B2(G148gat), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n883), .A2(new_n891), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n876), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n297), .C1(new_n919), .C2(new_n656), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n910), .B1(new_n917), .B2(new_n920), .ZN(G1345gat));
  NAND3_X1  g720(.A1(new_n909), .A2(new_n301), .A3(new_n630), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n918), .A2(new_n693), .A3(new_n876), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n301), .ZN(G1346gat));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n302), .A3(new_n593), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n918), .A2(new_n594), .A3(new_n876), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n302), .ZN(G1347gat));
  AOI21_X1  g726(.A(new_n398), .B1(new_n853), .B2(new_n854), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n422), .A2(new_n428), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(G169gat), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n930), .A2(new_n931), .A3(new_n717), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n858), .A2(new_n428), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n552), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n932), .B1(new_n931), .B2(new_n936), .ZN(G1348gat));
  OAI21_X1  g736(.A(G176gat), .B1(new_n930), .B2(new_n694), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n694), .A2(G176gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n934), .B2(new_n939), .ZN(G1349gat));
  NAND3_X1  g739(.A1(new_n935), .A2(new_n206), .A3(new_n630), .ZN(new_n941));
  OAI21_X1  g740(.A(G183gat), .B1(new_n930), .B2(new_n693), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(KEYINPUT124), .A3(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n935), .A2(new_n207), .A3(new_n593), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n593), .A3(new_n929), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(KEYINPUT61), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n207), .B1(new_n947), .B2(KEYINPUT61), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n946), .B2(new_n949), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  NAND3_X1  g751(.A1(new_n463), .A2(new_n415), .A3(new_n342), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT126), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(new_n928), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n552), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n914), .A2(new_n915), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n757), .A2(new_n398), .A3(new_n428), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n552), .A2(G197gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(G1352gat));
  XNOR2_X1  g761(.A(KEYINPUT127), .B(G204gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n959), .B2(new_n694), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n694), .A2(new_n963), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n955), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT62), .Z(new_n967));
  NAND2_X1  g766(.A1(new_n964), .A2(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n955), .A2(new_n285), .A3(new_n630), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n630), .B(new_n958), .C1(new_n914), .C2(new_n915), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  AOI21_X1  g772(.A(G218gat), .B1(new_n955), .B2(new_n593), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n594), .A2(new_n284), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n974), .B1(new_n960), .B2(new_n975), .ZN(G1355gat));
endmodule


