

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798;

  INV_X2 U380 ( .A(G125), .ZN(n429) );
  OR2_X1 U381 ( .A1(n397), .A2(n658), .ZN(n564) );
  INV_X2 U382 ( .A(G953), .ZN(n554) );
  XOR2_X1 U383 ( .A(n568), .B(KEYINPUT39), .Z(n360) );
  NOR2_X1 U384 ( .A1(n452), .A2(KEYINPUT64), .ZN(n447) );
  NAND2_X1 U385 ( .A1(n364), .A2(n654), .ZN(n791) );
  NAND2_X1 U386 ( .A1(n647), .A2(n759), .ZN(n707) );
  NOR2_X1 U387 ( .A1(G953), .A2(G237), .ZN(n539) );
  NOR2_X1 U388 ( .A1(n791), .A2(n689), .ZN(n690) );
  INV_X1 U389 ( .A(n791), .ZN(n693) );
  XNOR2_X1 U390 ( .A(n366), .B(n365), .ZN(n364) );
  AND2_X1 U391 ( .A1(n646), .A2(n772), .ZN(n367) );
  XNOR2_X1 U392 ( .A(n370), .B(n360), .ZN(n423) );
  XNOR2_X1 U393 ( .A(n591), .B(KEYINPUT42), .ZN(n650) );
  INV_X1 U394 ( .A(n718), .ZN(n621) );
  XNOR2_X1 U395 ( .A(n361), .B(KEYINPUT38), .ZN(n702) );
  NAND2_X1 U396 ( .A1(n361), .A2(n406), .ZN(n405) );
  INV_X1 U397 ( .A(KEYINPUT48), .ZN(n365) );
  XNOR2_X1 U398 ( .A(G110), .B(G107), .ZN(n402) );
  NOR2_X1 U399 ( .A1(n666), .A2(n755), .ZN(n668) );
  NOR2_X1 U400 ( .A1(n686), .A2(n755), .ZN(n426) );
  NOR2_X1 U401 ( .A1(n680), .A2(n755), .ZN(n681) );
  NOR2_X1 U402 ( .A1(n673), .A2(n755), .ZN(n674) );
  NOR2_X1 U403 ( .A1(n738), .A2(n737), .ZN(n739) );
  BUF_X1 U404 ( .A(n749), .Z(n752) );
  XNOR2_X1 U405 ( .A(n657), .B(n454), .ZN(n452) );
  NOR2_X1 U406 ( .A1(n691), .A2(n661), .ZN(n411) );
  XNOR2_X1 U407 ( .A(n660), .B(KEYINPUT82), .ZN(n661) );
  NAND2_X1 U408 ( .A1(n368), .A2(n367), .ZN(n366) );
  NOR2_X1 U409 ( .A1(n616), .A2(n617), .ZN(n417) );
  XNOR2_X1 U410 ( .A(n651), .B(n369), .ZN(n368) );
  AND2_X1 U411 ( .A1(n363), .A2(n418), .ZN(n387) );
  AND2_X1 U412 ( .A1(n413), .A2(n607), .ZN(n617) );
  NAND2_X1 U413 ( .A1(n470), .A2(n471), .ZN(n469) );
  NAND2_X1 U414 ( .A1(n604), .A2(n472), .ZN(n606) );
  NAND2_X1 U415 ( .A1(n371), .A2(n567), .ZN(n370) );
  OR2_X1 U416 ( .A1(n732), .A2(n590), .ZN(n591) );
  BUF_X1 U417 ( .A(n602), .Z(n624) );
  INV_X1 U418 ( .A(n566), .ZN(n371) );
  XNOR2_X1 U419 ( .A(n410), .B(KEYINPUT0), .ZN(n602) );
  NOR2_X1 U420 ( .A1(n506), .A2(n505), .ZN(n524) );
  NAND2_X1 U421 ( .A1(n407), .A2(n405), .ZN(n636) );
  AND2_X1 U422 ( .A1(n409), .A2(n408), .ZN(n407) );
  INV_X2 U423 ( .A(n593), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n428), .B(n486), .ZN(n570) );
  XNOR2_X1 U425 ( .A(n397), .B(n677), .ZN(n678) );
  XNOR2_X1 U426 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U427 ( .A(n402), .B(G104), .ZN(n558) );
  XNOR2_X1 U428 ( .A(n473), .B(G140), .ZN(n396) );
  XNOR2_X1 U429 ( .A(G902), .B(KEYINPUT15), .ZN(n655) );
  INV_X1 U430 ( .A(KEYINPUT46), .ZN(n369) );
  XOR2_X1 U431 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n473) );
  INV_X1 U432 ( .A(n362), .ZN(n691) );
  NAND2_X1 U433 ( .A1(n656), .A2(n362), .ZN(n657) );
  XNOR2_X2 U434 ( .A(n398), .B(n384), .ZN(n362) );
  NOR2_X1 U435 ( .A1(n372), .A2(n694), .ZN(n695) );
  NAND2_X1 U436 ( .A1(n690), .A2(n362), .ZN(n425) );
  AND2_X1 U437 ( .A1(n363), .A2(n415), .ZN(n388) );
  NAND2_X1 U438 ( .A1(n700), .A2(KEYINPUT34), .ZN(n363) );
  INV_X1 U439 ( .A(n423), .ZN(n648) );
  INV_X1 U440 ( .A(n691), .ZN(n372) );
  NOR2_X2 U441 ( .A1(n682), .A2(G902), .ZN(n390) );
  XNOR2_X2 U442 ( .A(n786), .B(n504), .ZN(n682) );
  AND2_X1 U443 ( .A1(n465), .A2(n610), .ZN(n389) );
  NOR2_X2 U444 ( .A1(n373), .A2(n374), .ZN(n446) );
  NOR2_X1 U445 ( .A1(n592), .A2(n463), .ZN(n373) );
  AND2_X1 U446 ( .A1(n718), .A2(KEYINPUT73), .ZN(n374) );
  NAND2_X1 U447 ( .A1(n445), .A2(n444), .ZN(n375) );
  NAND2_X1 U448 ( .A1(n445), .A2(n444), .ZN(n613) );
  XNOR2_X2 U449 ( .A(n515), .B(n499), .ZN(n786) );
  NAND2_X1 U450 ( .A1(n644), .A2(n434), .ZN(n431) );
  NOR2_X1 U451 ( .A1(KEYINPUT77), .A2(n435), .ZN(n434) );
  NAND2_X1 U452 ( .A1(n433), .A2(KEYINPUT47), .ZN(n432) );
  INV_X1 U453 ( .A(n707), .ZN(n433) );
  AND2_X1 U454 ( .A1(n607), .A2(n438), .ZN(n587) );
  AND2_X1 U455 ( .A1(n714), .A2(n571), .ZN(n438) );
  XNOR2_X1 U456 ( .A(n480), .B(G137), .ZN(n498) );
  INV_X1 U457 ( .A(KEYINPUT70), .ZN(n480) );
  NAND2_X1 U458 ( .A1(n467), .A2(n614), .ZN(n466) );
  NAND2_X1 U459 ( .A1(n624), .A2(KEYINPUT34), .ZN(n467) );
  OR2_X1 U460 ( .A1(n662), .A2(G902), .ZN(n517) );
  XNOR2_X1 U461 ( .A(n460), .B(n459), .ZN(n559) );
  XNOR2_X1 U462 ( .A(G128), .B(KEYINPUT23), .ZN(n476) );
  XNOR2_X1 U463 ( .A(n498), .B(n394), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n395), .B(G119), .ZN(n394) );
  INV_X1 U465 ( .A(G110), .ZN(n395) );
  XOR2_X1 U466 ( .A(G122), .B(KEYINPUT97), .Z(n541) );
  XNOR2_X1 U467 ( .A(n548), .B(n421), .ZN(n420) );
  INV_X1 U468 ( .A(G113), .ZN(n421) );
  XNOR2_X1 U469 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U470 ( .A(G143), .B(G104), .ZN(n546) );
  XNOR2_X1 U471 ( .A(G101), .B(G146), .ZN(n501) );
  AND2_X1 U472 ( .A1(n577), .A2(n441), .ZN(n427) );
  INV_X1 U473 ( .A(G237), .ZN(n518) );
  NOR2_X1 U474 ( .A1(n465), .A2(n610), .ZN(n442) );
  INV_X1 U475 ( .A(KEYINPUT73), .ZN(n464) );
  NOR2_X1 U476 ( .A1(n701), .A2(KEYINPUT19), .ZN(n406) );
  XNOR2_X1 U477 ( .A(G146), .B(G137), .ZN(n510) );
  NOR2_X1 U478 ( .A1(n645), .A2(n430), .ZN(n646) );
  NAND2_X1 U479 ( .A1(n431), .A2(n432), .ZN(n430) );
  INV_X1 U480 ( .A(n383), .ZN(n451) );
  NAND2_X1 U481 ( .A1(G234), .A2(G237), .ZN(n490) );
  NOR2_X2 U482 ( .A1(n702), .A2(n701), .ZN(n706) );
  INV_X1 U483 ( .A(n624), .ZN(n470) );
  INV_X1 U484 ( .A(G902), .ZN(n551) );
  AND2_X1 U485 ( .A1(n584), .A2(n583), .ZN(n703) );
  XOR2_X1 U486 ( .A(KEYINPUT101), .B(G107), .Z(n527) );
  XNOR2_X1 U487 ( .A(G116), .B(G122), .ZN(n526) );
  INV_X1 U488 ( .A(G128), .ZN(n495) );
  NAND2_X1 U489 ( .A1(n425), .A2(n382), .ZN(n696) );
  AND2_X1 U490 ( .A1(n589), .A2(n588), .ZN(n637) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n588) );
  INV_X1 U492 ( .A(KEYINPUT28), .ZN(n436) );
  NOR2_X1 U493 ( .A1(n466), .A2(n615), .ZN(n415) );
  INV_X1 U494 ( .A(n466), .ZN(n418) );
  XNOR2_X1 U495 ( .A(n662), .B(KEYINPUT62), .ZN(n663) );
  XNOR2_X1 U496 ( .A(n559), .B(n458), .ZN(n776) );
  XNOR2_X1 U497 ( .A(n479), .B(n478), .ZN(n481) );
  XNOR2_X1 U498 ( .A(n788), .B(n393), .ZN(n422) );
  XNOR2_X1 U499 ( .A(n788), .B(n420), .ZN(n549) );
  XNOR2_X1 U500 ( .A(n682), .B(n683), .ZN(n684) );
  XOR2_X1 U501 ( .A(KEYINPUT87), .B(n665), .Z(n755) );
  XNOR2_X1 U502 ( .A(n404), .B(n403), .ZN(n616) );
  INV_X1 U503 ( .A(KEYINPUT32), .ZN(n403) );
  XNOR2_X1 U504 ( .A(n462), .B(KEYINPUT65), .ZN(n413) );
  XNOR2_X1 U505 ( .A(n620), .B(KEYINPUT104), .ZN(n688) );
  XNOR2_X1 U506 ( .A(n392), .B(KEYINPUT85), .ZN(n619) );
  AND2_X1 U507 ( .A1(n451), .A2(n453), .ZN(n376) );
  AND2_X1 U508 ( .A1(n688), .A2(n627), .ZN(n377) );
  INV_X1 U509 ( .A(n716), .ZN(n461) );
  XOR2_X1 U510 ( .A(KEYINPUT16), .B(G122), .Z(n378) );
  XOR2_X1 U511 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n379) );
  AND2_X1 U512 ( .A1(n577), .A2(n461), .ZN(n380) );
  AND2_X1 U513 ( .A1(n632), .A2(n608), .ZN(n381) );
  INV_X1 U514 ( .A(n769), .ZN(n647) );
  XNOR2_X1 U515 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n615) );
  NAND2_X1 U516 ( .A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(n382) );
  XOR2_X1 U517 ( .A(n659), .B(KEYINPUT67), .Z(n383) );
  XOR2_X1 U518 ( .A(KEYINPUT81), .B(KEYINPUT45), .Z(n384) );
  XNOR2_X1 U519 ( .A(n422), .B(n481), .ZN(n748) );
  INV_X1 U520 ( .A(KEYINPUT47), .ZN(n435) );
  INV_X1 U521 ( .A(KEYINPUT64), .ZN(n453) );
  AND2_X1 U522 ( .A1(n383), .A2(KEYINPUT64), .ZN(n385) );
  XNOR2_X1 U523 ( .A(n613), .B(n612), .ZN(n386) );
  XNOR2_X1 U524 ( .A(n375), .B(n612), .ZN(n700) );
  NAND2_X1 U525 ( .A1(n388), .A2(n412), .ZN(n414) );
  NAND2_X1 U526 ( .A1(n416), .A2(n414), .ZN(n745) );
  INV_X1 U527 ( .A(n446), .ZN(n424) );
  XNOR2_X2 U528 ( .A(n390), .B(G469), .ZN(n576) );
  NAND2_X1 U529 ( .A1(n391), .A2(n615), .ZN(n416) );
  NAND2_X1 U530 ( .A1(n387), .A2(n412), .ZN(n391) );
  XNOR2_X1 U531 ( .A(n557), .B(n456), .ZN(n455) );
  XNOR2_X1 U532 ( .A(n401), .B(n379), .ZN(n457) );
  NAND2_X1 U533 ( .A1(n609), .A2(n427), .ZN(n392) );
  XNOR2_X1 U534 ( .A(n400), .B(n439), .ZN(n399) );
  XNOR2_X2 U535 ( .A(n396), .B(n401), .ZN(n788) );
  XNOR2_X2 U536 ( .A(n429), .B(G146), .ZN(n401) );
  XNOR2_X1 U537 ( .A(n455), .B(n776), .ZN(n397) );
  NAND2_X1 U538 ( .A1(n399), .A2(n377), .ZN(n398) );
  NAND2_X1 U539 ( .A1(n745), .A2(n417), .ZN(n400) );
  NAND2_X1 U540 ( .A1(n609), .A2(n381), .ZN(n404) );
  XNOR2_X2 U541 ( .A(n606), .B(n605), .ZN(n609) );
  NAND2_X1 U542 ( .A1(n361), .A2(n582), .ZN(n629) );
  NAND2_X1 U543 ( .A1(n701), .A2(KEYINPUT19), .ZN(n408) );
  NAND2_X1 U544 ( .A1(n593), .A2(KEYINPUT19), .ZN(n409) );
  NAND2_X1 U545 ( .A1(n636), .A2(n597), .ZN(n410) );
  NOR2_X1 U546 ( .A1(n411), .A2(n376), .ZN(n450) );
  NOR2_X1 U547 ( .A1(n697), .A2(n411), .ZN(n698) );
  INV_X1 U548 ( .A(n468), .ZN(n412) );
  NAND2_X1 U549 ( .A1(n424), .A2(KEYINPUT105), .ZN(n444) );
  NAND2_X1 U550 ( .A1(n419), .A2(n639), .ZN(n641) );
  NAND2_X1 U551 ( .A1(n635), .A2(n643), .ZN(n419) );
  AND2_X2 U552 ( .A1(n573), .A2(n584), .ZN(n769) );
  NAND2_X1 U553 ( .A1(n423), .A2(n769), .ZN(n649) );
  NAND2_X1 U554 ( .A1(n531), .A2(G221), .ZN(n479) );
  XNOR2_X1 U555 ( .A(n474), .B(n475), .ZN(n531) );
  NOR2_X1 U556 ( .A1(n442), .A2(n441), .ZN(n440) );
  NAND2_X1 U557 ( .A1(n446), .A2(n389), .ZN(n443) );
  NOR2_X1 U558 ( .A1(n386), .A2(n469), .ZN(n468) );
  XNOR2_X1 U559 ( .A(n426), .B(n687), .ZN(G54) );
  XNOR2_X1 U560 ( .A(n558), .B(n378), .ZN(n458) );
  AND2_X2 U561 ( .A1(n443), .A2(n440), .ZN(n445) );
  XNOR2_X1 U562 ( .A(n507), .B(KEYINPUT3), .ZN(n459) );
  NAND2_X1 U563 ( .A1(n748), .A2(n551), .ZN(n428) );
  NAND2_X1 U564 ( .A1(n587), .A2(n716), .ZN(n437) );
  INV_X1 U565 ( .A(KEYINPUT44), .ZN(n439) );
  INV_X1 U566 ( .A(n618), .ZN(n441) );
  NAND2_X1 U567 ( .A1(n446), .A2(n465), .ZN(n611) );
  NOR2_X4 U568 ( .A1(n448), .A2(n447), .ZN(n749) );
  NAND2_X1 U569 ( .A1(n449), .A2(n450), .ZN(n448) );
  NAND2_X1 U570 ( .A1(n452), .A2(n385), .ZN(n449) );
  XNOR2_X2 U571 ( .A(n564), .B(n563), .ZN(n593) );
  INV_X1 U572 ( .A(KEYINPUT79), .ZN(n454) );
  XNOR2_X1 U573 ( .A(n457), .B(n556), .ZN(n456) );
  XNOR2_X2 U574 ( .A(n525), .B(KEYINPUT4), .ZN(n557) );
  XNOR2_X1 U575 ( .A(n508), .B(n509), .ZN(n460) );
  NAND2_X1 U576 ( .A1(n609), .A2(n380), .ZN(n462) );
  NAND2_X1 U577 ( .A1(n621), .A2(n464), .ZN(n463) );
  NAND2_X1 U578 ( .A1(n592), .A2(KEYINPUT73), .ZN(n465) );
  XNOR2_X2 U579 ( .A(n576), .B(n575), .ZN(n592) );
  INV_X1 U580 ( .A(KEYINPUT34), .ZN(n471) );
  AND2_X1 U581 ( .A1(n703), .A2(n603), .ZN(n472) );
  INV_X1 U582 ( .A(KEYINPUT105), .ZN(n610) );
  INV_X1 U583 ( .A(n498), .ZN(n499) );
  INV_X1 U584 ( .A(KEYINPUT33), .ZN(n612) );
  BUF_X1 U585 ( .A(n386), .Z(n733) );
  XNOR2_X1 U586 ( .A(n649), .B(KEYINPUT40), .ZN(n743) );
  NAND2_X1 U587 ( .A1(G234), .A2(n554), .ZN(n475) );
  XOR2_X1 U588 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n474) );
  XOR2_X1 U589 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n477) );
  XNOR2_X1 U590 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U591 ( .A1(n655), .A2(G234), .ZN(n482) );
  XNOR2_X1 U592 ( .A(n482), .B(KEYINPUT20), .ZN(n483) );
  XNOR2_X1 U593 ( .A(KEYINPUT92), .B(n483), .ZN(n487) );
  NAND2_X1 U594 ( .A1(G217), .A2(n487), .ZN(n485) );
  XNOR2_X1 U595 ( .A(KEYINPUT25), .B(KEYINPUT93), .ZN(n484) );
  XNOR2_X1 U596 ( .A(n485), .B(n484), .ZN(n486) );
  NAND2_X1 U597 ( .A1(n487), .A2(G221), .ZN(n489) );
  INV_X1 U598 ( .A(KEYINPUT21), .ZN(n488) );
  XNOR2_X1 U599 ( .A(n489), .B(n488), .ZN(n714) );
  XNOR2_X1 U600 ( .A(n714), .B(KEYINPUT94), .ZN(n603) );
  NAND2_X1 U601 ( .A1(n570), .A2(n603), .ZN(n718) );
  XNOR2_X1 U602 ( .A(n490), .B(KEYINPUT14), .ZN(n699) );
  NAND2_X1 U603 ( .A1(G953), .A2(G900), .ZN(n493) );
  NOR2_X1 U604 ( .A1(G953), .A2(G952), .ZN(n492) );
  NOR2_X1 U605 ( .A1(G902), .A2(n554), .ZN(n491) );
  NOR2_X1 U606 ( .A1(n492), .A2(n491), .ZN(n594) );
  AND2_X1 U607 ( .A1(n493), .A2(n594), .ZN(n494) );
  AND2_X1 U608 ( .A1(n699), .A2(n494), .ZN(n571) );
  NAND2_X1 U609 ( .A1(n621), .A2(n571), .ZN(n506) );
  XNOR2_X2 U610 ( .A(G143), .B(KEYINPUT76), .ZN(n496) );
  XNOR2_X2 U611 ( .A(n496), .B(n495), .ZN(n525) );
  XNOR2_X1 U612 ( .A(G134), .B(G131), .ZN(n497) );
  XNOR2_X2 U613 ( .A(n557), .B(n497), .ZN(n515) );
  NAND2_X1 U614 ( .A1(n554), .A2(G227), .ZN(n500) );
  XNOR2_X1 U615 ( .A(n500), .B(G140), .ZN(n502) );
  XNOR2_X1 U616 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U617 ( .A(n503), .B(n558), .ZN(n504) );
  BUF_X1 U618 ( .A(n576), .Z(n505) );
  XNOR2_X1 U619 ( .A(G119), .B(G116), .ZN(n508) );
  XNOR2_X1 U620 ( .A(KEYINPUT71), .B(KEYINPUT88), .ZN(n507) );
  XNOR2_X1 U621 ( .A(G113), .B(G101), .ZN(n509) );
  NAND2_X1 U622 ( .A1(n539), .A2(G210), .ZN(n511) );
  XNOR2_X1 U623 ( .A(n511), .B(n510), .ZN(n513) );
  XNOR2_X1 U624 ( .A(KEYINPUT74), .B(KEYINPUT5), .ZN(n512) );
  XNOR2_X1 U625 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U626 ( .A(n559), .B(n514), .ZN(n516) );
  XNOR2_X1 U627 ( .A(n515), .B(n516), .ZN(n662) );
  XNOR2_X2 U628 ( .A(n517), .B(G472), .ZN(n716) );
  NAND2_X1 U629 ( .A1(n551), .A2(n518), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n560), .A2(G214), .ZN(n520) );
  INV_X1 U631 ( .A(KEYINPUT90), .ZN(n519) );
  XNOR2_X1 U632 ( .A(n520), .B(n519), .ZN(n701) );
  INV_X1 U633 ( .A(n701), .ZN(n582) );
  NAND2_X1 U634 ( .A1(n716), .A2(n582), .ZN(n522) );
  XNOR2_X1 U635 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n521) );
  XNOR2_X1 U636 ( .A(n522), .B(n521), .ZN(n523) );
  NAND2_X1 U637 ( .A1(n524), .A2(n523), .ZN(n566) );
  XNOR2_X1 U638 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U639 ( .A(n525), .B(n528), .ZN(n535) );
  XOR2_X1 U640 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n530) );
  XNOR2_X1 U641 ( .A(G134), .B(KEYINPUT100), .ZN(n529) );
  XNOR2_X1 U642 ( .A(n530), .B(n529), .ZN(n533) );
  NAND2_X1 U643 ( .A1(G217), .A2(n531), .ZN(n532) );
  XNOR2_X1 U644 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U645 ( .A(n535), .B(n534), .ZN(n753) );
  NOR2_X1 U646 ( .A1(G902), .A2(n753), .ZN(n536) );
  XOR2_X1 U647 ( .A(G478), .B(n536), .Z(n538) );
  INV_X1 U648 ( .A(KEYINPUT102), .ZN(n537) );
  XNOR2_X1 U649 ( .A(n538), .B(n537), .ZN(n584) );
  NAND2_X1 U650 ( .A1(G214), .A2(n539), .ZN(n540) );
  XNOR2_X1 U651 ( .A(n541), .B(n540), .ZN(n545) );
  XOR2_X1 U652 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n543) );
  XNOR2_X1 U653 ( .A(G131), .B(KEYINPUT11), .ZN(n542) );
  XNOR2_X1 U654 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U655 ( .A(n545), .B(n544), .Z(n550) );
  XOR2_X1 U656 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n547) );
  XNOR2_X1 U657 ( .A(n550), .B(n549), .ZN(n670) );
  NAND2_X1 U658 ( .A1(n670), .A2(n551), .ZN(n553) );
  XOR2_X1 U659 ( .A(KEYINPUT13), .B(G475), .Z(n552) );
  XNOR2_X1 U660 ( .A(n553), .B(n552), .ZN(n573) );
  INV_X1 U661 ( .A(n573), .ZN(n583) );
  NOR2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n614) );
  NAND2_X1 U663 ( .A1(n554), .A2(G224), .ZN(n555) );
  XNOR2_X1 U664 ( .A(n555), .B(KEYINPUT75), .ZN(n556) );
  INV_X1 U665 ( .A(n655), .ZN(n658) );
  NAND2_X1 U666 ( .A1(n560), .A2(G210), .ZN(n562) );
  INV_X1 U667 ( .A(KEYINPUT89), .ZN(n561) );
  XNOR2_X1 U668 ( .A(n562), .B(n561), .ZN(n563) );
  NAND2_X1 U669 ( .A1(n614), .A2(n361), .ZN(n565) );
  OR2_X1 U670 ( .A1(n566), .A2(n565), .ZN(n640) );
  XNOR2_X1 U671 ( .A(n640), .B(G143), .ZN(G45) );
  INV_X1 U672 ( .A(n702), .ZN(n567) );
  INV_X1 U673 ( .A(KEYINPUT84), .ZN(n568) );
  INV_X1 U674 ( .A(n584), .ZN(n569) );
  NAND2_X1 U675 ( .A1(n569), .A2(n583), .ZN(n759) );
  OR2_X1 U676 ( .A1(n648), .A2(n759), .ZN(n652) );
  XNOR2_X1 U677 ( .A(n652), .B(G134), .ZN(G36) );
  INV_X1 U678 ( .A(n570), .ZN(n607) );
  XNOR2_X1 U679 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n572) );
  XNOR2_X1 U680 ( .A(n716), .B(n572), .ZN(n618) );
  AND2_X1 U681 ( .A1(n618), .A2(n769), .ZN(n574) );
  AND2_X1 U682 ( .A1(n587), .A2(n574), .ZN(n628) );
  AND2_X1 U683 ( .A1(n628), .A2(n582), .ZN(n578) );
  XNOR2_X1 U684 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n575) );
  BUF_X1 U685 ( .A(n592), .Z(n577) );
  NAND2_X1 U686 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U687 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n579) );
  XNOR2_X1 U688 ( .A(n580), .B(n579), .ZN(n581) );
  NAND2_X1 U689 ( .A1(n581), .A2(n593), .ZN(n653) );
  XNOR2_X1 U690 ( .A(n653), .B(G140), .ZN(G42) );
  NAND2_X1 U691 ( .A1(n706), .A2(n703), .ZN(n586) );
  INV_X1 U692 ( .A(KEYINPUT41), .ZN(n585) );
  XNOR2_X1 U693 ( .A(n586), .B(n585), .ZN(n732) );
  INV_X1 U694 ( .A(n505), .ZN(n589) );
  INV_X1 U695 ( .A(n637), .ZN(n590) );
  XNOR2_X1 U696 ( .A(n650), .B(G137), .ZN(G39) );
  NAND2_X1 U697 ( .A1(n611), .A2(n716), .ZN(n723) );
  NAND2_X1 U698 ( .A1(G953), .A2(G898), .ZN(n595) );
  AND2_X1 U699 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U700 ( .A1(n699), .A2(n596), .ZN(n597) );
  NOR2_X1 U701 ( .A1(n723), .A2(n624), .ZN(n599) );
  XOR2_X1 U702 ( .A(KEYINPUT95), .B(KEYINPUT31), .Z(n598) );
  XNOR2_X1 U703 ( .A(n599), .B(n598), .ZN(n625) );
  NOR2_X1 U704 ( .A1(n625), .A2(n759), .ZN(n600) );
  XOR2_X1 U705 ( .A(G116), .B(n600), .Z(G18) );
  NOR2_X1 U706 ( .A1(n625), .A2(n647), .ZN(n601) );
  XOR2_X1 U707 ( .A(G113), .B(n601), .Z(G15) );
  INV_X1 U708 ( .A(n602), .ZN(n604) );
  INV_X1 U709 ( .A(KEYINPUT22), .ZN(n605) );
  INV_X1 U710 ( .A(n577), .ZN(n632) );
  INV_X1 U711 ( .A(n607), .ZN(n713) );
  NOR2_X1 U712 ( .A1(n618), .A2(n713), .ZN(n608) );
  XOR2_X1 U713 ( .A(G119), .B(n616), .Z(G21) );
  XOR2_X1 U714 ( .A(n617), .B(G110), .Z(G12) );
  NAND2_X1 U715 ( .A1(n619), .A2(n713), .ZN(n620) );
  NAND2_X1 U716 ( .A1(n621), .A2(n461), .ZN(n622) );
  OR2_X1 U717 ( .A1(n622), .A2(n505), .ZN(n623) );
  OR2_X1 U718 ( .A1(n624), .A2(n623), .ZN(n757) );
  NAND2_X1 U719 ( .A1(n625), .A2(n757), .ZN(n626) );
  NAND2_X1 U720 ( .A1(n626), .A2(n707), .ZN(n627) );
  XOR2_X1 U721 ( .A(KEYINPUT108), .B(n628), .Z(n630) );
  NOR2_X1 U722 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U723 ( .A(n631), .B(KEYINPUT36), .ZN(n633) );
  NAND2_X1 U724 ( .A1(n633), .A2(n632), .ZN(n772) );
  INV_X1 U725 ( .A(KEYINPUT77), .ZN(n643) );
  XNOR2_X1 U726 ( .A(KEYINPUT72), .B(n707), .ZN(n634) );
  NAND2_X1 U727 ( .A1(n634), .A2(n435), .ZN(n635) );
  NAND2_X1 U728 ( .A1(n637), .A2(n636), .ZN(n764) );
  OR2_X1 U729 ( .A1(KEYINPUT47), .A2(n643), .ZN(n638) );
  NAND2_X1 U730 ( .A1(n764), .A2(n638), .ZN(n639) );
  NAND2_X1 U731 ( .A1(n641), .A2(n640), .ZN(n645) );
  INV_X1 U732 ( .A(KEYINPUT72), .ZN(n642) );
  OR2_X1 U733 ( .A1(n764), .A2(n642), .ZN(n644) );
  NAND2_X1 U734 ( .A1(n743), .A2(n650), .ZN(n651) );
  AND2_X1 U735 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U736 ( .A1(n791), .A2(n655), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n658), .A2(KEYINPUT2), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n693), .A2(KEYINPUT2), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n749), .A2(G472), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n664), .B(n663), .ZN(n666) );
  NOR2_X1 U741 ( .A1(n554), .A2(G952), .ZN(n665) );
  INV_X1 U742 ( .A(KEYINPUT63), .ZN(n667) );
  XNOR2_X1 U743 ( .A(n668), .B(n667), .ZN(G57) );
  NAND2_X1 U744 ( .A1(n749), .A2(G475), .ZN(n672) );
  XNOR2_X1 U745 ( .A(KEYINPUT118), .B(KEYINPUT59), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U747 ( .A(n674), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U748 ( .A1(n749), .A2(G210), .ZN(n679) );
  XOR2_X1 U749 ( .A(KEYINPUT116), .B(KEYINPUT54), .Z(n676) );
  XNOR2_X1 U750 ( .A(KEYINPUT55), .B(KEYINPUT86), .ZN(n675) );
  XNOR2_X1 U751 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U752 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U753 ( .A(n681), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U754 ( .A(KEYINPUT117), .ZN(n687) );
  NAND2_X1 U755 ( .A1(n749), .A2(G469), .ZN(n685) );
  XOR2_X1 U756 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n683) );
  XNOR2_X1 U757 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n688), .B(G101), .ZN(G3) );
  INV_X1 U759 ( .A(KEYINPUT78), .ZN(n689) );
  NOR2_X1 U760 ( .A1(KEYINPUT2), .A2(KEYINPUT78), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U763 ( .A(n698), .B(KEYINPUT80), .ZN(n738) );
  NAND2_X1 U764 ( .A1(G952), .A2(n699), .ZN(n731) );
  INV_X1 U765 ( .A(n733), .ZN(n712) );
  NAND2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U767 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U768 ( .A(KEYINPUT111), .B(n705), .Z(n710) );
  NAND2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U770 ( .A(n708), .B(KEYINPUT112), .ZN(n709) );
  NAND2_X1 U771 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U772 ( .A1(n712), .A2(n711), .ZN(n728) );
  NOR2_X1 U773 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U774 ( .A(KEYINPUT49), .B(n715), .Z(n717) );
  NOR2_X1 U775 ( .A1(n717), .A2(n716), .ZN(n721) );
  NAND2_X1 U776 ( .A1(n577), .A2(n718), .ZN(n719) );
  XNOR2_X1 U777 ( .A(n719), .B(KEYINPUT50), .ZN(n720) );
  NAND2_X1 U778 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U779 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U780 ( .A(KEYINPUT51), .B(n724), .Z(n726) );
  INV_X1 U781 ( .A(n732), .ZN(n725) );
  NAND2_X1 U782 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U783 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U784 ( .A(KEYINPUT52), .B(n729), .Z(n730) );
  NOR2_X1 U785 ( .A1(n731), .A2(n730), .ZN(n735) );
  NOR2_X1 U786 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U787 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U788 ( .A(n736), .B(KEYINPUT113), .ZN(n737) );
  XNOR2_X1 U789 ( .A(n739), .B(KEYINPUT114), .ZN(n740) );
  NAND2_X1 U790 ( .A1(n740), .A2(n554), .ZN(n742) );
  XNOR2_X1 U791 ( .A(KEYINPUT115), .B(KEYINPUT53), .ZN(n741) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(G75) );
  XNOR2_X1 U793 ( .A(G131), .B(KEYINPUT127), .ZN(n744) );
  XOR2_X1 U794 ( .A(n744), .B(n743), .Z(G33) );
  BUF_X1 U795 ( .A(n745), .Z(n746) );
  XNOR2_X1 U796 ( .A(G122), .B(KEYINPUT126), .ZN(n747) );
  XNOR2_X1 U797 ( .A(n746), .B(n747), .ZN(G24) );
  NAND2_X1 U798 ( .A1(n752), .A2(G217), .ZN(n750) );
  XOR2_X1 U799 ( .A(n748), .B(n750), .Z(n751) );
  NOR2_X1 U800 ( .A1(n751), .A2(n755), .ZN(G66) );
  NAND2_X1 U801 ( .A1(n752), .A2(G478), .ZN(n754) );
  XNOR2_X1 U802 ( .A(n754), .B(n753), .ZN(n756) );
  NOR2_X1 U803 ( .A1(n756), .A2(n755), .ZN(G63) );
  INV_X1 U804 ( .A(n757), .ZN(n760) );
  NAND2_X1 U805 ( .A1(n760), .A2(n769), .ZN(n758) );
  XNOR2_X1 U806 ( .A(n758), .B(G104), .ZN(G6) );
  XOR2_X1 U807 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n762) );
  INV_X1 U808 ( .A(n759), .ZN(n765) );
  NAND2_X1 U809 ( .A1(n760), .A2(n765), .ZN(n761) );
  XNOR2_X1 U810 ( .A(n762), .B(n761), .ZN(n763) );
  XNOR2_X1 U811 ( .A(G107), .B(n763), .ZN(G9) );
  XOR2_X1 U812 ( .A(KEYINPUT109), .B(KEYINPUT29), .Z(n767) );
  INV_X1 U813 ( .A(n764), .ZN(n770) );
  NAND2_X1 U814 ( .A1(n770), .A2(n765), .ZN(n766) );
  XNOR2_X1 U815 ( .A(n767), .B(n766), .ZN(n768) );
  XOR2_X1 U816 ( .A(G128), .B(n768), .Z(G30) );
  NAND2_X1 U817 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U818 ( .A(n771), .B(G146), .ZN(G48) );
  XOR2_X1 U819 ( .A(KEYINPUT110), .B(n772), .Z(n773) );
  XNOR2_X1 U820 ( .A(n773), .B(KEYINPUT37), .ZN(n774) );
  XNOR2_X1 U821 ( .A(G125), .B(n774), .ZN(G27) );
  NOR2_X1 U822 ( .A1(G898), .A2(n554), .ZN(n775) );
  NOR2_X1 U823 ( .A1(n776), .A2(n775), .ZN(n784) );
  NAND2_X1 U824 ( .A1(n372), .A2(n554), .ZN(n777) );
  XOR2_X1 U825 ( .A(KEYINPUT120), .B(n777), .Z(n782) );
  NAND2_X1 U826 ( .A1(G953), .A2(G224), .ZN(n778) );
  XNOR2_X1 U827 ( .A(KEYINPUT61), .B(n778), .ZN(n779) );
  NAND2_X1 U828 ( .A1(n779), .A2(G898), .ZN(n780) );
  XNOR2_X1 U829 ( .A(KEYINPUT119), .B(n780), .ZN(n781) );
  NOR2_X1 U830 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U831 ( .A(n784), .B(n783), .Z(n785) );
  XOR2_X1 U832 ( .A(KEYINPUT121), .B(n785), .Z(G69) );
  XOR2_X1 U833 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n787) );
  XNOR2_X1 U834 ( .A(n788), .B(n787), .ZN(n789) );
  XNOR2_X1 U835 ( .A(n786), .B(n789), .ZN(n793) );
  XOR2_X1 U836 ( .A(KEYINPUT124), .B(n793), .Z(n790) );
  XNOR2_X1 U837 ( .A(n791), .B(n790), .ZN(n792) );
  NAND2_X1 U838 ( .A1(n792), .A2(n554), .ZN(n798) );
  XNOR2_X1 U839 ( .A(n793), .B(G227), .ZN(n794) );
  XNOR2_X1 U840 ( .A(n794), .B(KEYINPUT125), .ZN(n795) );
  NAND2_X1 U841 ( .A1(n795), .A2(G900), .ZN(n796) );
  NAND2_X1 U842 ( .A1(n796), .A2(G953), .ZN(n797) );
  NAND2_X1 U843 ( .A1(n798), .A2(n797), .ZN(G72) );
endmodule

