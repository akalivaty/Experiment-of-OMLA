//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NOR3_X1   g008(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n189), .B2(new_n191), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G137), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n202), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(G137), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G134), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(G131), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n212), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n204), .A2(new_n202), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n209), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n214), .A2(KEYINPUT66), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n222), .B(G131), .C1(new_n208), .C2(new_n213), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n221), .B1(new_n220), .B2(new_n223), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n201), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G116), .B(G119), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT2), .B(G113), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n192), .A2(G128), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n189), .B(new_n191), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n211), .A2(new_n209), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n219), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n226), .A2(new_n229), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT26), .B(G101), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n241), .B(KEYINPUT69), .ZN(new_n242));
  INV_X1    g056(.A(G237), .ZN(new_n243));
  INV_X1    g057(.A(G953), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(G210), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n242), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT29), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n237), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n220), .A2(new_n223), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT67), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n252), .B1(new_n256), .B2(new_n201), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(new_n229), .ZN(new_n258));
  INV_X1    g072(.A(new_n238), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n240), .B(new_n251), .C1(new_n260), .C2(new_n239), .ZN(new_n261));
  INV_X1    g075(.A(G902), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n229), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n226), .B2(new_n237), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n220), .A2(new_n201), .A3(new_n223), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n237), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(KEYINPUT30), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n264), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n238), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT76), .B1(new_n271), .B2(new_n249), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT76), .ZN(new_n273));
  AOI211_X1 g087(.A(new_n273), .B(new_n248), .C1(new_n270), .C2(new_n238), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n272), .A2(new_n274), .A3(KEYINPUT29), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n268), .B2(new_n264), .ZN(new_n277));
  AOI211_X1 g091(.A(KEYINPUT72), .B(new_n229), .C1(new_n267), .C2(new_n237), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n279), .A2(new_n238), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n248), .B(new_n240), .C1(new_n280), .C2(new_n239), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT75), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n239), .B1(new_n279), .B2(new_n238), .ZN(new_n283));
  INV_X1    g097(.A(new_n240), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n248), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n263), .B1(new_n275), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G472), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n187), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n286), .B1(new_n285), .B2(new_n248), .ZN(new_n292));
  NOR4_X1   g106(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT75), .A4(new_n249), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n269), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(new_n257), .B2(new_n265), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n259), .B1(new_n296), .B2(new_n264), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n273), .B1(new_n297), .B2(new_n248), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n271), .A2(KEYINPUT76), .A3(new_n249), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n250), .A3(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT77), .B(G472), .C1(new_n301), .C2(new_n263), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n291), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT70), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n238), .A2(new_n304), .A3(new_n248), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n270), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n304), .B1(new_n238), .B2(new_n248), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT71), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n238), .A2(new_n248), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT70), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n310), .A2(new_n270), .A3(new_n311), .A4(new_n305), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n308), .A2(KEYINPUT31), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n249), .B1(new_n283), .B2(new_n284), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT31), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n310), .A2(new_n270), .A3(new_n315), .A4(new_n305), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(KEYINPUT32), .A3(new_n290), .A4(new_n262), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT74), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n290), .A3(new_n262), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(KEYINPUT74), .A3(new_n323), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n303), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n328), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n328), .B2(KEYINPUT81), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT81), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(G125), .A3(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n329), .B1(new_n334), .B2(KEYINPUT16), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n335), .A2(G146), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(G146), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XOR2_X1   g152(.A(G119), .B(G128), .Z(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT24), .B(G110), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n342));
  INV_X1    g156(.A(G119), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n342), .B1(new_n343), .B2(G128), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n344), .A2(KEYINPUT23), .B1(new_n343), .B2(G128), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(KEYINPUT23), .B2(new_n344), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT80), .ZN(new_n347));
  INV_X1    g161(.A(G110), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n338), .B(new_n341), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n339), .A2(new_n340), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n346), .B2(G110), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n354), .A2(KEYINPUT83), .A3(G146), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT83), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n352), .B(KEYINPUT82), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(new_n188), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n337), .B(new_n351), .C1(new_n355), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n349), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT22), .B(G137), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n244), .A2(G221), .A3(G234), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n349), .A2(KEYINPUT84), .A3(new_n359), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n362), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n349), .A2(new_n359), .A3(new_n365), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n262), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT25), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n368), .A2(new_n372), .A3(new_n262), .A4(new_n369), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT78), .B(G217), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(G234), .B2(new_n262), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n368), .A2(new_n369), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n375), .A2(G902), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n234), .A2(new_n328), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n244), .A2(G224), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT7), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n199), .B1(new_n196), .B2(new_n197), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n383), .B(new_n385), .C1(new_n328), .C2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n328), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n231), .A2(new_n233), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G125), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT7), .B(new_n384), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n343), .A2(G116), .ZN(new_n392));
  INV_X1    g206(.A(G116), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G119), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT5), .ZN(new_n395));
  OR3_X1    g209(.A1(new_n393), .A2(KEYINPUT5), .A3(G119), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n396), .A3(G113), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT2), .B(G113), .Z(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n227), .ZN(new_n399));
  INV_X1    g213(.A(G104), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT3), .B1(new_n400), .B2(G107), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n402));
  INV_X1    g216(.A(G107), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G104), .ZN(new_n404));
  INV_X1    g218(.A(G101), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(G107), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n401), .A2(new_n404), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n400), .A2(G107), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n403), .A2(G104), .ZN(new_n409));
  OAI21_X1  g223(.A(G101), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n397), .A2(new_n399), .A3(new_n407), .A4(new_n410), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n397), .A2(new_n399), .B1(new_n407), .B2(new_n410), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT91), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n397), .A2(new_n399), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n407), .A2(new_n410), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n415), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(KEYINPUT90), .B(KEYINPUT8), .Z(new_n419));
  XNOR2_X1  g233(.A(G110), .B(G122), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n387), .B(new_n391), .C1(new_n418), .C2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n401), .A2(new_n404), .A3(new_n406), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n423), .A2(new_n424), .A3(G101), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n229), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(G101), .ZN(new_n427));
  AND4_X1   g241(.A1(KEYINPUT86), .A2(new_n427), .A3(KEYINPUT4), .A4(new_n407), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n424), .B1(new_n423), .B2(G101), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT86), .B1(new_n429), .B2(new_n407), .ZN(new_n430));
  OAI211_X1 g244(.A(KEYINPUT89), .B(new_n426), .C1(new_n428), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n411), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n427), .A2(KEYINPUT4), .A3(new_n407), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n429), .A2(KEYINPUT86), .A3(new_n407), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT89), .B1(new_n437), .B2(new_n426), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n422), .B1(new_n439), .B2(new_n420), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n382), .B1(new_n440), .B2(G902), .ZN(new_n441));
  INV_X1    g255(.A(new_n420), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n432), .B2(new_n438), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n426), .B1(new_n428), .B2(new_n430), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n446), .A2(new_n431), .A3(new_n411), .A4(new_n420), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n443), .A2(KEYINPUT6), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n388), .A2(new_n390), .ZN(new_n449));
  INV_X1    g263(.A(new_n384), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n452), .B(new_n442), .C1(new_n432), .C2(new_n438), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n448), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G210), .B1(G237), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(new_n447), .ZN(new_n456));
  OAI211_X1 g270(.A(KEYINPUT92), .B(new_n262), .C1(new_n456), .C2(new_n422), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n441), .A2(new_n454), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n441), .A2(new_n457), .A3(new_n454), .ZN(new_n460));
  INV_X1    g274(.A(new_n455), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(KEYINPUT93), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT93), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n460), .A2(new_n464), .A3(new_n461), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G214), .B1(G237), .B2(G902), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT88), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G469), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n389), .A2(new_n416), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n231), .A2(new_n233), .A3(new_n407), .A4(new_n410), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND4_X1   g288(.A1(KEYINPUT12), .A2(new_n474), .A3(new_n223), .A4(new_n220), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n474), .B1(new_n224), .B2(new_n225), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n386), .A2(new_n425), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n428), .B2(new_n430), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n407), .A2(new_n410), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n234), .A2(KEYINPUT87), .A3(new_n481), .A4(KEYINPUT10), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT10), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(new_n473), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n473), .A2(new_n484), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n480), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(new_n256), .ZN(new_n489));
  XNOR2_X1  g303(.A(G110), .B(G140), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n244), .A2(G227), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n490), .B(new_n491), .Z(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n478), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n224), .A2(new_n225), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(new_n486), .A3(new_n480), .A4(new_n487), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n488), .A2(new_n256), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n471), .B(new_n262), .C1(new_n494), .C2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n493), .B1(new_n478), .B2(new_n489), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n496), .A2(new_n497), .A3(new_n492), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(G469), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n471), .A2(new_n262), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT9), .B(G234), .ZN(new_n506));
  OAI21_X1  g320(.A(G221), .B1(new_n506), .B2(G902), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(KEYINPUT85), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n393), .A3(G122), .ZN(new_n512));
  INV_X1    g326(.A(G122), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT14), .B1(new_n513), .B2(G116), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(G116), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G107), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT99), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(KEYINPUT99), .A3(G107), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(G116), .B(G122), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n522), .A2(KEYINPUT95), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(KEYINPUT95), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n403), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT98), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n232), .A2(G143), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT96), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n190), .A2(G128), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n528), .A3(new_n531), .ZN(new_n534));
  AOI21_X1  g348(.A(G134), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n534), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n536), .A2(new_n532), .A3(new_n203), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n527), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n203), .B1(new_n536), .B2(new_n532), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n531), .B(KEYINPUT13), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n530), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n540), .B1(new_n543), .B2(new_n203), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(KEYINPUT97), .A3(G134), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n523), .A2(G107), .A3(new_n524), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n526), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n539), .A2(new_n544), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n374), .A2(new_n506), .A3(G953), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n538), .A2(new_n548), .A3(new_n550), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G478), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n554), .A2(KEYINPUT100), .A3(new_n262), .A4(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n538), .A2(new_n548), .A3(new_n550), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n550), .B1(new_n538), .B2(new_n548), .ZN(new_n559));
  OAI211_X1 g373(.A(KEYINPUT100), .B(new_n262), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n556), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT100), .B1(new_n554), .B2(new_n262), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n557), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(G234), .A2(G237), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(G952), .A3(new_n244), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT21), .B(G898), .Z(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(G902), .A3(G953), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n569), .B(KEYINPUT101), .Z(new_n570));
  NAND3_X1  g384(.A1(new_n243), .A2(new_n244), .A3(G214), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(new_n190), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G131), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n571), .B(G143), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n218), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n574), .A2(new_n218), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT17), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n577), .A2(new_n579), .A3(new_n336), .A4(new_n337), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT83), .B1(new_n354), .B2(G146), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n357), .A2(new_n356), .A3(new_n188), .ZN(new_n582));
  INV_X1    g396(.A(new_n334), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n581), .A2(new_n582), .B1(G146), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n578), .A2(KEYINPUT18), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT18), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n574), .B1(new_n586), .B2(new_n218), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n580), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(G113), .B(G122), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(new_n400), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n580), .B(new_n591), .C1(new_n584), .C2(new_n588), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT94), .B(G475), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OAI22_X1  g412(.A1(new_n355), .A2(new_n358), .B1(new_n188), .B2(new_n334), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n585), .A3(new_n587), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n573), .A2(new_n575), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT19), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n583), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n354), .B2(new_n602), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n337), .B(new_n601), .C1(new_n604), .C2(G146), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n591), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n594), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(G475), .A2(G902), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT20), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT20), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n612), .B(new_n609), .C1(new_n606), .C2(new_n607), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n598), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n564), .A2(new_n570), .A3(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n470), .A2(new_n510), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n327), .A2(new_n381), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  AOI21_X1  g432(.A(new_n468), .B1(new_n462), .B2(new_n458), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n554), .A2(KEYINPUT33), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n552), .B2(new_n553), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n262), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(G478), .ZN(new_n625));
  INV_X1    g439(.A(new_n614), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n554), .A2(new_n555), .A3(new_n262), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n570), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n620), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT102), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n318), .A2(new_n262), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G472), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n380), .A2(new_n510), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n633), .A2(new_n321), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  INV_X1    g452(.A(new_n564), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n614), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n620), .A2(new_n629), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NAND2_X1  g458(.A1(new_n633), .A2(new_n321), .ZN(new_n645));
  INV_X1    g459(.A(new_n367), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT84), .B1(new_n349), .B2(new_n359), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT103), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n362), .A2(new_n649), .A3(new_n367), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n366), .A2(KEYINPUT36), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n648), .B(new_n650), .C1(KEYINPUT36), .C2(new_n366), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(new_n378), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n376), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n645), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n616), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  NOR2_X1   g475(.A1(new_n620), .A2(new_n657), .ZN(new_n662));
  INV_X1    g476(.A(new_n640), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n568), .A2(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n566), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n510), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n327), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  AND2_X1   g483(.A1(new_n308), .A2(new_n312), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n260), .A2(new_n248), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n262), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n325), .A2(new_n326), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n564), .A2(new_n614), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n657), .A2(new_n469), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n665), .B(KEYINPUT39), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n505), .A2(new_n509), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n466), .B(KEYINPUT38), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n675), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  INV_X1    g499(.A(new_n665), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n628), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n510), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n327), .A2(new_n662), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  INV_X1    g505(.A(new_n327), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n494), .A2(new_n498), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n262), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n695), .A2(new_n499), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n509), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n692), .A2(new_n380), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n631), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NAND2_X1  g515(.A1(new_n698), .A2(new_n641), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  NAND4_X1  g517(.A1(new_n695), .A2(new_n509), .A3(new_n499), .A4(new_n570), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n704), .A2(new_n626), .A3(new_n639), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n327), .A2(new_n662), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  NOR2_X1   g521(.A1(G472), .A2(G902), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n240), .B1(new_n260), .B2(new_n239), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n249), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n313), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n316), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n709), .B1(new_n313), .B2(new_n711), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n708), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n380), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n619), .A2(new_n676), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n704), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n715), .A2(new_n717), .A3(new_n719), .A4(new_n633), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n290), .B1(new_n318), .B2(new_n262), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n313), .A2(new_n711), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n316), .A3(new_n712), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n723), .B1(new_n726), .B2(new_n708), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(KEYINPUT106), .A3(new_n717), .A4(new_n719), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n722), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  INV_X1    g544(.A(new_n697), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n619), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n688), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n715), .A2(new_n633), .A3(new_n656), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT107), .B(G125), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G27));
  NAND2_X1  g551(.A1(new_n462), .A2(KEYINPUT93), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n469), .A3(new_n465), .A4(new_n458), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT110), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n463), .A2(new_n741), .A3(new_n469), .A4(new_n465), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n502), .A2(KEYINPUT108), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n500), .A2(new_n501), .A3(new_n744), .A4(G469), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n743), .A2(new_n499), .A3(new_n504), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n509), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT109), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n746), .A2(new_n749), .A3(new_n509), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n740), .A2(new_n742), .A3(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n327), .A2(new_n381), .A3(new_n687), .A4(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n717), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n321), .B(KEYINPUT32), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n756), .B1(new_n757), .B2(new_n303), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n687), .A2(new_n740), .A3(new_n742), .A4(new_n751), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(KEYINPUT42), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  INV_X1    g576(.A(new_n666), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n327), .A2(new_n381), .A3(new_n763), .A4(new_n752), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NOR2_X1   g579(.A1(new_n558), .A2(new_n559), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n622), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n554), .A2(KEYINPUT33), .ZN(new_n768));
  AOI21_X1  g582(.A(G902), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n627), .B1(new_n769), .B2(new_n555), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT43), .B1(new_n770), .B2(new_n626), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n625), .A2(new_n772), .A3(new_n614), .A4(new_n627), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n771), .A2(new_n656), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n645), .A2(new_n774), .A3(KEYINPUT44), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n740), .A2(new_n742), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT46), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n500), .A2(new_n501), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT45), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(KEYINPUT45), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n471), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n779), .B1(new_n783), .B2(new_n503), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT111), .ZN(new_n785));
  OR3_X1    g599(.A1(new_n783), .A2(new_n779), .A3(new_n503), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n787), .B(new_n779), .C1(new_n783), .C2(new_n503), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n785), .A2(new_n499), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n509), .A3(new_n678), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT112), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n789), .A2(new_n792), .A3(new_n509), .A4(new_n678), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n778), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n645), .A2(new_n774), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(KEYINPUT113), .A3(new_n796), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  NAND2_X1  g617(.A1(new_n789), .A2(new_n509), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT47), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n789), .A2(KEYINPUT47), .A3(new_n509), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n777), .A2(new_n380), .A3(new_n687), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n692), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  XNOR2_X1  g626(.A(new_n696), .B(KEYINPUT49), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n770), .A2(new_n626), .A3(new_n468), .A4(new_n508), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n717), .A3(new_n814), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n675), .A2(new_n815), .A3(new_n683), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n727), .A2(new_n717), .ZN(new_n818));
  INV_X1    g632(.A(new_n566), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n771), .A2(new_n819), .A3(new_n773), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n731), .A2(new_n468), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n822), .A2(new_n683), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT50), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n777), .A2(new_n381), .A3(new_n819), .A4(new_n731), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n675), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n626), .B1(new_n625), .B2(new_n627), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n776), .A2(new_n697), .A3(new_n820), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n827), .A2(new_n828), .B1(new_n734), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT117), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n696), .A2(new_n508), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n777), .B(new_n821), .C1(new_n808), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT116), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n817), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n758), .A2(new_n829), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n836), .A2(KEYINPUT118), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(KEYINPUT118), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(KEYINPUT48), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(KEYINPUT48), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n826), .A2(new_n628), .A3(new_n675), .ZN(new_n842));
  OAI211_X1 g656(.A(G952), .B(new_n244), .C1(new_n822), .C2(new_n732), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n833), .A2(KEYINPUT51), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n817), .A2(KEYINPUT117), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n825), .B(new_n830), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n835), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n657), .A2(new_n665), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n852), .B2(new_n747), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n656), .A2(new_n686), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(KEYINPUT114), .A3(new_n509), .A4(new_n746), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n718), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n675), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n668), .A2(new_n690), .A3(new_n735), .A4(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT52), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n629), .B1(new_n628), .B2(new_n640), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n860), .A2(new_n469), .A3(new_n466), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n616), .A2(new_n658), .B1(new_n861), .B2(new_n635), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n617), .A2(new_n729), .A3(new_n706), .A4(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n321), .A2(KEYINPUT74), .A3(new_n323), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n324), .B2(new_n320), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n380), .B1(new_n865), .B2(new_n303), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n866), .B(new_n731), .C1(new_n631), .C2(new_n641), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n639), .A2(new_n626), .A3(new_n686), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n509), .A3(new_n505), .A4(new_n656), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n776), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n327), .A2(new_n870), .B1(new_n734), .B2(new_n759), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n871), .A2(new_n764), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n863), .A2(new_n761), .A3(new_n867), .A4(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n850), .B1(new_n859), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n668), .A2(new_n735), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(KEYINPUT52), .A3(new_n690), .A4(new_n857), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n858), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n729), .A2(new_n706), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n617), .A2(new_n862), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n867), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n871), .A2(new_n764), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n755), .B2(new_n760), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n879), .A2(KEYINPUT53), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n874), .A2(KEYINPUT54), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT54), .B1(new_n874), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n849), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  INV_X1    g703(.A(new_n873), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT53), .B1(new_n890), .B2(new_n879), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n859), .A2(new_n873), .A3(new_n850), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n874), .A2(new_n885), .A3(KEYINPUT54), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(KEYINPUT115), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n848), .B1(new_n888), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(G952), .A2(G953), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n816), .B1(new_n896), .B2(new_n897), .ZN(G75));
  OR2_X1    g712(.A1(new_n244), .A2(G952), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT120), .Z(new_n900));
  AOI21_X1  g714(.A(new_n262), .B1(new_n874), .B2(new_n885), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT56), .B1(new_n901), .B2(new_n461), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n448), .A2(new_n453), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n451), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n900), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n901), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n461), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n906), .B1(new_n909), .B2(new_n911), .ZN(G51));
  INV_X1    g726(.A(new_n900), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n908), .A2(new_n783), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n893), .A2(new_n894), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n503), .B(KEYINPUT57), .Z(new_n916));
  OAI21_X1  g730(.A(new_n693), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n913), .B1(new_n914), .B2(new_n917), .ZN(G54));
  OAI21_X1  g732(.A(G902), .B1(new_n891), .B2(new_n892), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n907), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n901), .A2(KEYINPUT119), .ZN(new_n921));
  AND2_X1   g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n608), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n920), .A2(new_n608), .A3(new_n921), .A4(new_n922), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n913), .B1(new_n925), .B2(new_n926), .ZN(G60));
  INV_X1    g741(.A(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n767), .A2(new_n768), .ZN(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n555), .A2(new_n262), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n886), .A2(new_n887), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n928), .B1(new_n934), .B2(new_n913), .ZN(new_n935));
  OAI211_X1 g749(.A(KEYINPUT122), .B(new_n900), .C1(new_n915), .C2(new_n933), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n888), .A2(new_n895), .A3(new_n932), .ZN(new_n937));
  INV_X1    g751(.A(new_n929), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n935), .A2(new_n936), .B1(new_n937), .B2(new_n938), .ZN(G63));
  XNOR2_X1  g753(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT124), .ZN(new_n941));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n941), .B(new_n942), .Z(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n874), .B2(new_n885), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n944), .A2(new_n377), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n653), .A3(new_n654), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n945), .A2(new_n900), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n945), .A2(KEYINPUT61), .A3(new_n900), .A4(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(G66));
  NAND3_X1  g765(.A1(new_n567), .A2(G224), .A3(G953), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n867), .A2(new_n880), .A3(new_n881), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n903), .B1(G898), .B2(new_n244), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n954), .B(new_n955), .Z(G69));
  AOI21_X1  g770(.A(new_n244), .B1(G227), .B2(G900), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n296), .B(new_n604), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n679), .B1(new_n628), .B2(new_n640), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n866), .A2(new_n777), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n799), .A2(new_n800), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n778), .A2(new_n791), .A3(new_n793), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n811), .B(new_n962), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n668), .A2(new_n690), .A3(new_n684), .A4(new_n735), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n967), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n960), .B1(new_n970), .B2(G953), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n960), .B1(G900), .B2(G953), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n809), .B1(new_n806), .B2(new_n807), .ZN(new_n973));
  AOI22_X1  g787(.A1(new_n794), .A2(new_n801), .B1(new_n692), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n875), .A2(new_n690), .ZN(new_n975));
  INV_X1    g789(.A(new_n718), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n791), .A2(new_n758), .A3(new_n976), .A4(new_n793), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n977), .A2(new_n764), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n974), .A2(new_n975), .A3(new_n761), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n972), .B1(new_n979), .B2(G953), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n971), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT126), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n971), .B2(new_n980), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT126), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n959), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n985), .A2(new_n986), .ZN(new_n989));
  AOI211_X1 g803(.A(KEYINPUT126), .B(new_n983), .C1(new_n971), .C2(new_n980), .ZN(new_n990));
  INV_X1    g804(.A(new_n959), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n988), .A2(new_n992), .ZN(G72));
  XNOR2_X1  g807(.A(new_n271), .B(KEYINPUT127), .ZN(new_n994));
  OR3_X1    g808(.A1(new_n979), .A2(new_n248), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n248), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n970), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n953), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  NAND2_X1  g815(.A1(new_n298), .A2(new_n299), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1001), .B1(new_n671), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(new_n874), .B2(new_n885), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n994), .B(new_n249), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n900), .B1(new_n1005), .B2(new_n1001), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n999), .A2(new_n1004), .A3(new_n1006), .ZN(G57));
endmodule


