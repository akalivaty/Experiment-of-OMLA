

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716;

  NAND2_X1 U374 ( .A1(n591), .A2(n592), .ZN(n588) );
  INV_X1 U375 ( .A(G953), .ZN(n707) );
  NOR2_X2 U376 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X2 U377 ( .A(n393), .B(G134), .ZN(n433) );
  XNOR2_X2 U378 ( .A(n372), .B(n371), .ZN(n393) );
  XNOR2_X2 U379 ( .A(n572), .B(n571), .ZN(n685) );
  NOR2_X1 U380 ( .A1(n591), .A2(n544), .ZN(n646) );
  NOR2_X1 U381 ( .A1(n712), .A2(n716), .ZN(n520) );
  XNOR2_X1 U382 ( .A(n519), .B(KEYINPUT39), .ZN(n529) );
  XNOR2_X1 U383 ( .A(G475), .B(n419), .ZN(n513) );
  OR2_X1 U384 ( .A1(n667), .A2(G902), .ZN(n374) );
  XNOR2_X1 U385 ( .A(n413), .B(KEYINPUT70), .ZN(n431) );
  XNOR2_X1 U386 ( .A(G131), .B(KEYINPUT71), .ZN(n413) );
  INV_X1 U387 ( .A(n558), .ZN(n351) );
  XNOR2_X1 U388 ( .A(n500), .B(n373), .ZN(n589) );
  XNOR2_X2 U389 ( .A(n422), .B(n421), .ZN(n467) );
  XOR2_X2 U390 ( .A(G119), .B(KEYINPUT3), .Z(n422) );
  XNOR2_X1 U391 ( .A(n474), .B(n473), .ZN(n630) );
  XNOR2_X1 U392 ( .A(n428), .B(n355), .ZN(n491) );
  NAND2_X1 U393 ( .A1(n630), .A2(n477), .ZN(n360) );
  NAND2_X1 U394 ( .A1(n574), .A2(n575), .ZN(n623) );
  XNOR2_X1 U395 ( .A(G137), .B(G140), .ZN(n449) );
  XOR2_X1 U396 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n410) );
  XNOR2_X1 U397 ( .A(n431), .B(n416), .ZN(n367) );
  XNOR2_X1 U398 ( .A(G113), .B(G143), .ZN(n406) );
  XOR2_X1 U399 ( .A(G104), .B(G140), .Z(n408) );
  INV_X1 U400 ( .A(KEYINPUT64), .ZN(n371) );
  XOR2_X1 U401 ( .A(KEYINPUT4), .B(KEYINPUT69), .Z(n430) );
  XOR2_X1 U402 ( .A(KEYINPUT68), .B(G101), .Z(n429) );
  XNOR2_X1 U403 ( .A(G146), .B(G125), .ZN(n414) );
  XNOR2_X1 U404 ( .A(G104), .B(G107), .ZN(n420) );
  XNOR2_X1 U405 ( .A(G128), .B(G119), .ZN(n440) );
  XNOR2_X1 U406 ( .A(KEYINPUT10), .B(n414), .ZN(n695) );
  XNOR2_X1 U407 ( .A(n429), .B(n414), .ZN(n392) );
  XNOR2_X1 U408 ( .A(n427), .B(n388), .ZN(n387) );
  XNOR2_X1 U409 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n388) );
  XNOR2_X1 U410 ( .A(n540), .B(n539), .ZN(n610) );
  INV_X1 U411 ( .A(KEYINPUT33), .ZN(n539) );
  AND2_X1 U412 ( .A1(n653), .A2(n354), .ZN(n365) );
  XNOR2_X1 U413 ( .A(n503), .B(n492), .ZN(n535) );
  INV_X1 U414 ( .A(n493), .ZN(n482) );
  INV_X1 U415 ( .A(KEYINPUT1), .ZN(n373) );
  INV_X1 U416 ( .A(n595), .ZN(n381) );
  NOR2_X1 U417 ( .A1(n624), .A2(G902), .ZN(n418) );
  XNOR2_X1 U418 ( .A(n459), .B(n456), .ZN(n370) );
  INV_X1 U419 ( .A(KEYINPUT22), .ZN(n383) );
  XNOR2_X1 U420 ( .A(n632), .B(n631), .ZN(n633) );
  NOR2_X1 U421 ( .A1(G952), .A2(n707), .ZN(n680) );
  NOR2_X1 U422 ( .A1(G953), .A2(G237), .ZN(n464) );
  XNOR2_X1 U423 ( .A(KEYINPUT23), .B(KEYINPUT83), .ZN(n442) );
  XNOR2_X1 U424 ( .A(G113), .B(G116), .ZN(n421) );
  XNOR2_X1 U425 ( .A(n522), .B(KEYINPUT48), .ZN(n528) );
  XNOR2_X1 U426 ( .A(n520), .B(KEYINPUT46), .ZN(n521) );
  XNOR2_X1 U427 ( .A(G122), .B(G107), .ZN(n397) );
  XNOR2_X1 U428 ( .A(n415), .B(n366), .ZN(n624) );
  XNOR2_X1 U429 ( .A(n695), .B(n367), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n474), .B(n439), .ZN(n667) );
  INV_X1 U431 ( .A(n504), .ZN(n523) );
  XNOR2_X1 U432 ( .A(n541), .B(KEYINPUT34), .ZN(n364) );
  NOR2_X1 U433 ( .A1(n546), .A2(n554), .ZN(n378) );
  NOR2_X2 U434 ( .A1(n462), .A2(n588), .ZN(n563) );
  OR2_X2 U435 ( .A1(n535), .A2(n352), .ZN(n538) );
  XNOR2_X1 U436 ( .A(n695), .B(n451), .ZN(n452) );
  XNOR2_X1 U437 ( .A(n450), .B(KEYINPUT90), .ZN(n451) );
  AND2_X2 U438 ( .A1(n623), .A2(n622), .ZN(n676) );
  AND2_X1 U439 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U440 ( .A(n392), .B(n387), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n369), .B(n356), .ZN(n712) );
  NOR2_X1 U442 ( .A1(n504), .A2(n503), .ZN(n506) );
  XNOR2_X1 U443 ( .A(n363), .B(n361), .ZN(n713) );
  XNOR2_X1 U444 ( .A(n362), .B(KEYINPUT79), .ZN(n361) );
  NAND2_X1 U445 ( .A1(n364), .A2(n532), .ZN(n363) );
  INV_X1 U446 ( .A(KEYINPUT35), .ZN(n362) );
  XNOR2_X1 U447 ( .A(n375), .B(KEYINPUT32), .ZN(n715) );
  NOR2_X1 U448 ( .A1(n553), .A2(n376), .ZN(n375) );
  XNOR2_X1 U449 ( .A(n378), .B(n377), .ZN(n376) );
  INV_X1 U450 ( .A(KEYINPUT80), .ZN(n377) );
  NAND2_X1 U451 ( .A1(n382), .A2(n380), .ZN(n544) );
  AND2_X1 U452 ( .A1(n351), .A2(n381), .ZN(n380) );
  NOR2_X1 U453 ( .A1(n513), .A2(n487), .ZN(n653) );
  NOR2_X1 U454 ( .A1(n680), .A2(n635), .ZN(n638) );
  NOR2_X1 U455 ( .A1(G953), .A2(n616), .ZN(n618) );
  XNOR2_X1 U456 ( .A(n649), .B(n368), .ZN(G30) );
  INV_X1 U457 ( .A(G128), .ZN(n368) );
  OR2_X1 U458 ( .A1(n534), .A2(n357), .ZN(n352) );
  XOR2_X1 U459 ( .A(G472), .B(KEYINPUT73), .Z(n353) );
  AND2_X1 U460 ( .A1(n494), .A2(n592), .ZN(n354) );
  AND2_X1 U461 ( .A1(G210), .A2(n463), .ZN(n355) );
  XNOR2_X1 U462 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n356) );
  AND2_X1 U463 ( .A1(G898), .A2(G953), .ZN(n357) );
  XOR2_X1 U464 ( .A(n624), .B(KEYINPUT59), .Z(n358) );
  XNOR2_X1 U465 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n359) );
  XNOR2_X2 U466 ( .A(n360), .B(n353), .ZN(n502) );
  XNOR2_X2 U467 ( .A(n700), .B(n434), .ZN(n474) );
  NAND2_X1 U468 ( .A1(n554), .A2(n365), .ZN(n504) );
  AND2_X2 U469 ( .A1(n543), .A2(n562), .ZN(n379) );
  NAND2_X1 U470 ( .A1(n529), .A2(n653), .ZN(n369) );
  XNOR2_X2 U471 ( .A(n457), .B(n370), .ZN(n591) );
  INV_X1 U472 ( .A(n393), .ZN(n426) );
  XNOR2_X2 U473 ( .A(G143), .B(G128), .ZN(n372) );
  XNOR2_X2 U474 ( .A(n374), .B(G469), .ZN(n500) );
  XNOR2_X2 U475 ( .A(n379), .B(n383), .ZN(n553) );
  NAND2_X1 U476 ( .A1(n491), .A2(n579), .ZN(n503) );
  INV_X1 U477 ( .A(n553), .ZN(n382) );
  XNOR2_X1 U478 ( .A(n688), .B(n384), .ZN(n662) );
  XNOR2_X1 U479 ( .A(n386), .B(n385), .ZN(n384) );
  XNOR2_X1 U480 ( .A(n425), .B(n426), .ZN(n385) );
  NOR2_X1 U481 ( .A1(n626), .A2(n680), .ZN(n629) );
  XNOR2_X1 U482 ( .A(n625), .B(n358), .ZN(n626) );
  NAND2_X1 U483 ( .A1(n676), .A2(G475), .ZN(n625) );
  XNOR2_X1 U484 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n662), .B(n359), .ZN(n663) );
  AND2_X1 U487 ( .A1(n576), .A2(KEYINPUT2), .ZN(n389) );
  XNOR2_X1 U488 ( .A(KEYINPUT72), .B(n511), .ZN(n390) );
  AND2_X1 U489 ( .A1(n485), .A2(n484), .ZN(n391) );
  XNOR2_X1 U490 ( .A(n468), .B(n467), .ZN(n472) );
  NAND2_X1 U491 ( .A1(n559), .A2(n554), .ZN(n540) );
  XNOR2_X1 U492 ( .A(n472), .B(n471), .ZN(n473) );
  AND2_X1 U493 ( .A1(n483), .A2(n482), .ZN(n484) );
  INV_X1 U494 ( .A(KEYINPUT77), .ZN(n454) );
  INV_X1 U495 ( .A(KEYINPUT45), .ZN(n571) );
  XNOR2_X1 U496 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U497 ( .A(n636), .B(KEYINPUT63), .ZN(n637) );
  XNOR2_X1 U498 ( .A(n627), .B(KEYINPUT60), .ZN(n628) );
  XNOR2_X1 U499 ( .A(n618), .B(n617), .ZN(G75) );
  XOR2_X1 U500 ( .A(KEYINPUT7), .B(KEYINPUT99), .Z(n395) );
  XNOR2_X1 U501 ( .A(KEYINPUT9), .B(KEYINPUT100), .ZN(n394) );
  XNOR2_X1 U502 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U503 ( .A(n433), .B(n396), .ZN(n404) );
  XOR2_X1 U504 ( .A(KEYINPUT101), .B(KEYINPUT98), .Z(n398) );
  XNOR2_X1 U505 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U506 ( .A(G116), .B(n399), .Z(n402) );
  NAND2_X1 U507 ( .A1(G234), .A2(n707), .ZN(n400) );
  XOR2_X1 U508 ( .A(KEYINPUT8), .B(n400), .Z(n446) );
  NAND2_X1 U509 ( .A1(G217), .A2(n446), .ZN(n401) );
  XNOR2_X1 U510 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U511 ( .A(n404), .B(n403), .ZN(n674) );
  NOR2_X1 U512 ( .A1(G902), .A2(n674), .ZN(n405) );
  XOR2_X1 U513 ( .A(G478), .B(n405), .Z(n487) );
  XNOR2_X1 U514 ( .A(n406), .B(KEYINPUT12), .ZN(n416) );
  NAND2_X1 U515 ( .A1(G214), .A2(n464), .ZN(n407) );
  XNOR2_X1 U516 ( .A(n408), .B(n407), .ZN(n412) );
  XNOR2_X1 U517 ( .A(G122), .B(KEYINPUT95), .ZN(n409) );
  XNOR2_X1 U518 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U519 ( .A(n412), .B(n411), .Z(n415) );
  XNOR2_X1 U520 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n417) );
  XNOR2_X1 U521 ( .A(n418), .B(n417), .ZN(n419) );
  AND2_X1 U522 ( .A1(n513), .A2(n487), .ZN(n655) );
  NOR2_X1 U523 ( .A1(n653), .A2(n655), .ZN(n584) );
  NAND2_X1 U524 ( .A1(n584), .A2(KEYINPUT47), .ZN(n489) );
  XNOR2_X1 U525 ( .A(n420), .B(G110), .ZN(n435) );
  XOR2_X1 U526 ( .A(n435), .B(KEYINPUT16), .Z(n424) );
  XNOR2_X1 U527 ( .A(n467), .B(G122), .ZN(n423) );
  XNOR2_X1 U528 ( .A(n424), .B(n423), .ZN(n688) );
  XNOR2_X1 U529 ( .A(n430), .B(KEYINPUT86), .ZN(n425) );
  NAND2_X1 U530 ( .A1(G224), .A2(n707), .ZN(n427) );
  XNOR2_X1 U531 ( .A(G902), .B(KEYINPUT15), .ZN(n619) );
  NAND2_X1 U532 ( .A1(n662), .A2(n619), .ZN(n428) );
  OR2_X1 U533 ( .A1(G237), .A2(G902), .ZN(n463) );
  BUF_X1 U534 ( .A(n491), .Z(n527) );
  XNOR2_X1 U535 ( .A(G146), .B(n429), .ZN(n434) );
  XNOR2_X2 U536 ( .A(n433), .B(n432), .ZN(n700) );
  INV_X1 U537 ( .A(n435), .ZN(n436) );
  XNOR2_X1 U538 ( .A(KEYINPUT89), .B(n449), .ZN(n696) );
  XNOR2_X1 U539 ( .A(n436), .B(n696), .ZN(n438) );
  NAND2_X1 U540 ( .A1(n707), .A2(G227), .ZN(n437) );
  XNOR2_X1 U541 ( .A(n438), .B(n437), .ZN(n439) );
  INV_X1 U542 ( .A(n500), .ZN(n462) );
  XOR2_X1 U543 ( .A(KEYINPUT78), .B(G110), .Z(n441) );
  XNOR2_X1 U544 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U545 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n443) );
  XNOR2_X1 U546 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U547 ( .A(n445), .B(n444), .Z(n448) );
  NAND2_X1 U548 ( .A1(G221), .A2(n446), .ZN(n447) );
  XNOR2_X1 U549 ( .A(n448), .B(n447), .ZN(n453) );
  INV_X1 U550 ( .A(n449), .ZN(n450) );
  XNOR2_X1 U551 ( .A(n453), .B(n452), .ZN(n678) );
  NOR2_X1 U552 ( .A1(G902), .A2(n678), .ZN(n457) );
  XNOR2_X1 U553 ( .A(KEYINPUT25), .B(KEYINPUT92), .ZN(n455) );
  NAND2_X1 U554 ( .A1(G234), .A2(n619), .ZN(n458) );
  XNOR2_X1 U555 ( .A(KEYINPUT20), .B(n458), .ZN(n460) );
  NAND2_X1 U556 ( .A1(n460), .A2(G217), .ZN(n459) );
  NAND2_X1 U557 ( .A1(n460), .A2(G221), .ZN(n461) );
  XOR2_X1 U558 ( .A(KEYINPUT21), .B(n461), .Z(n592) );
  XNOR2_X1 U559 ( .A(n563), .B(KEYINPUT104), .ZN(n485) );
  NAND2_X1 U560 ( .A1(G214), .A2(n463), .ZN(n579) );
  INV_X1 U561 ( .A(G902), .ZN(n477) );
  XOR2_X1 U562 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n466) );
  NAND2_X1 U563 ( .A1(n464), .A2(G210), .ZN(n465) );
  XOR2_X1 U564 ( .A(n466), .B(n465), .Z(n468) );
  XOR2_X1 U565 ( .A(KEYINPUT74), .B(KEYINPUT94), .Z(n470) );
  XNOR2_X1 U566 ( .A(G137), .B(KEYINPUT75), .ZN(n469) );
  XNOR2_X1 U567 ( .A(n470), .B(n469), .ZN(n471) );
  NAND2_X1 U568 ( .A1(n579), .A2(n502), .ZN(n475) );
  XOR2_X1 U569 ( .A(n475), .B(KEYINPUT30), .Z(n483) );
  NAND2_X1 U570 ( .A1(G234), .A2(G237), .ZN(n476) );
  XNOR2_X1 U571 ( .A(n476), .B(KEYINPUT14), .ZN(n578) );
  NAND2_X1 U572 ( .A1(G953), .A2(n477), .ZN(n478) );
  NAND2_X1 U573 ( .A1(n578), .A2(n478), .ZN(n480) );
  NOR2_X1 U574 ( .A1(G953), .A2(G952), .ZN(n479) );
  NOR2_X1 U575 ( .A1(n480), .A2(n479), .ZN(n533) );
  NAND2_X1 U576 ( .A1(G953), .A2(G900), .ZN(n481) );
  NAND2_X1 U577 ( .A1(n533), .A2(n481), .ZN(n493) );
  NAND2_X1 U578 ( .A1(n527), .A2(n391), .ZN(n486) );
  XNOR2_X1 U579 ( .A(KEYINPUT105), .B(n486), .ZN(n488) );
  INV_X1 U580 ( .A(n487), .ZN(n512) );
  NOR2_X1 U581 ( .A1(n513), .A2(n512), .ZN(n532) );
  NAND2_X1 U582 ( .A1(n488), .A2(n532), .ZN(n650) );
  NAND2_X1 U583 ( .A1(n489), .A2(n650), .ZN(n490) );
  XNOR2_X1 U584 ( .A(n490), .B(KEYINPUT82), .ZN(n510) );
  XOR2_X1 U585 ( .A(KEYINPUT76), .B(KEYINPUT19), .Z(n492) );
  NOR2_X1 U586 ( .A1(n591), .A2(n493), .ZN(n494) );
  BUF_X1 U587 ( .A(n502), .Z(n595) );
  NAND2_X1 U588 ( .A1(n354), .A2(n595), .ZN(n496) );
  XOR2_X1 U589 ( .A(KEYINPUT106), .B(KEYINPUT28), .Z(n495) );
  XNOR2_X1 U590 ( .A(n496), .B(n495), .ZN(n497) );
  NAND2_X1 U591 ( .A1(n497), .A2(n500), .ZN(n517) );
  NOR2_X2 U592 ( .A1(n535), .A2(n517), .ZN(n651) );
  XOR2_X1 U593 ( .A(n651), .B(KEYINPUT47), .Z(n499) );
  NAND2_X1 U594 ( .A1(n651), .A2(n584), .ZN(n498) );
  NAND2_X1 U595 ( .A1(n499), .A2(n498), .ZN(n508) );
  INV_X1 U596 ( .A(n589), .ZN(n558) );
  INV_X1 U597 ( .A(KEYINPUT6), .ZN(n501) );
  XNOR2_X1 U598 ( .A(n502), .B(n501), .ZN(n554) );
  XOR2_X1 U599 ( .A(KEYINPUT109), .B(KEYINPUT36), .Z(n505) );
  XNOR2_X1 U600 ( .A(n506), .B(n505), .ZN(n507) );
  NAND2_X1 U601 ( .A1(n558), .A2(n507), .ZN(n659) );
  NAND2_X1 U602 ( .A1(n508), .A2(n659), .ZN(n509) );
  NAND2_X1 U603 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U604 ( .A(KEYINPUT102), .B(n514), .ZN(n582) );
  XOR2_X1 U605 ( .A(KEYINPUT38), .B(n527), .Z(n580) );
  NAND2_X1 U606 ( .A1(n580), .A2(n579), .ZN(n583) );
  NOR2_X1 U607 ( .A1(n582), .A2(n583), .ZN(n516) );
  XNOR2_X1 U608 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n515) );
  XNOR2_X1 U609 ( .A(n516), .B(n515), .ZN(n611) );
  NOR2_X1 U610 ( .A1(n517), .A2(n611), .ZN(n518) );
  XNOR2_X1 U611 ( .A(n518), .B(KEYINPUT42), .ZN(n716) );
  NAND2_X1 U612 ( .A1(n391), .A2(n580), .ZN(n519) );
  NAND2_X1 U613 ( .A1(n390), .A2(n521), .ZN(n522) );
  NAND2_X1 U614 ( .A1(n523), .A2(n579), .ZN(n524) );
  NOR2_X1 U615 ( .A1(n558), .A2(n524), .ZN(n525) );
  XNOR2_X1 U616 ( .A(n525), .B(KEYINPUT43), .ZN(n526) );
  NOR2_X1 U617 ( .A1(n527), .A2(n526), .ZN(n661) );
  NOR2_X2 U618 ( .A1(n528), .A2(n661), .ZN(n704) );
  NAND2_X1 U619 ( .A1(n655), .A2(n529), .ZN(n703) );
  INV_X1 U620 ( .A(KEYINPUT81), .ZN(n530) );
  AND2_X1 U621 ( .A1(n703), .A2(n530), .ZN(n531) );
  AND2_X1 U622 ( .A1(n704), .A2(n531), .ZN(n573) );
  INV_X1 U623 ( .A(n533), .ZN(n534) );
  XOR2_X1 U624 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n536) );
  XNOR2_X1 U625 ( .A(KEYINPUT67), .B(n536), .ZN(n537) );
  XNOR2_X2 U626 ( .A(n538), .B(n537), .ZN(n562) );
  INV_X1 U627 ( .A(n562), .ZN(n560) );
  NOR2_X1 U628 ( .A1(n589), .A2(n588), .ZN(n559) );
  NOR2_X1 U629 ( .A1(n560), .A2(n610), .ZN(n541) );
  INV_X1 U630 ( .A(n592), .ZN(n542) );
  NOR2_X1 U631 ( .A1(n542), .A2(n582), .ZN(n543) );
  NOR2_X1 U632 ( .A1(n589), .A2(n591), .ZN(n545) );
  XNOR2_X1 U633 ( .A(n545), .B(KEYINPUT103), .ZN(n546) );
  NOR2_X1 U634 ( .A1(n646), .A2(n715), .ZN(n549) );
  INV_X1 U635 ( .A(KEYINPUT44), .ZN(n547) );
  NAND2_X1 U636 ( .A1(n549), .A2(n547), .ZN(n548) );
  OR2_X1 U637 ( .A1(n713), .A2(n548), .ZN(n552) );
  NOR2_X1 U638 ( .A1(n549), .A2(n547), .ZN(n550) );
  XNOR2_X1 U639 ( .A(n550), .B(KEYINPUT65), .ZN(n551) );
  NAND2_X1 U640 ( .A1(n552), .A2(n551), .ZN(n570) );
  NOR2_X1 U641 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U642 ( .A(KEYINPUT84), .B(n555), .ZN(n556) );
  NAND2_X1 U643 ( .A1(n556), .A2(n591), .ZN(n557) );
  NOR2_X1 U644 ( .A1(n558), .A2(n557), .ZN(n639) );
  NAND2_X1 U645 ( .A1(n595), .A2(n559), .ZN(n598) );
  NOR2_X1 U646 ( .A1(n560), .A2(n598), .ZN(n561) );
  XOR2_X1 U647 ( .A(KEYINPUT31), .B(n561), .Z(n656) );
  NAND2_X1 U648 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U649 ( .A1(n595), .A2(n564), .ZN(n641) );
  NOR2_X1 U650 ( .A1(n656), .A2(n641), .ZN(n565) );
  NOR2_X1 U651 ( .A1(n584), .A2(n565), .ZN(n566) );
  NOR2_X1 U652 ( .A1(n639), .A2(n566), .ZN(n568) );
  NAND2_X1 U653 ( .A1(n713), .A2(KEYINPUT44), .ZN(n567) );
  NAND2_X1 U654 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X2 U655 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U656 ( .A1(n573), .A2(n685), .ZN(n574) );
  INV_X1 U657 ( .A(KEYINPUT2), .ZN(n575) );
  XOR2_X1 U658 ( .A(n703), .B(KEYINPUT81), .Z(n576) );
  AND2_X1 U659 ( .A1(n704), .A2(n389), .ZN(n577) );
  NAND2_X1 U660 ( .A1(n577), .A2(n685), .ZN(n620) );
  NAND2_X1 U661 ( .A1(n623), .A2(n620), .ZN(n609) );
  NAND2_X1 U662 ( .A1(G952), .A2(n578), .ZN(n606) );
  NOR2_X1 U663 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U664 ( .A1(n582), .A2(n581), .ZN(n586) );
  NOR2_X1 U665 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U666 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U667 ( .A1(n587), .A2(n610), .ZN(n603) );
  NAND2_X1 U668 ( .A1(n351), .A2(n588), .ZN(n590) );
  XNOR2_X1 U669 ( .A(n590), .B(KEYINPUT50), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U671 ( .A(KEYINPUT49), .B(n593), .Z(n594) );
  NOR2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U675 ( .A(KEYINPUT51), .B(n600), .ZN(n601) );
  NOR2_X1 U676 ( .A1(n611), .A2(n601), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U678 ( .A(n604), .B(KEYINPUT52), .ZN(n605) );
  NOR2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT113), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n614) );
  NOR2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n612), .B(KEYINPUT114), .ZN(n613) );
  NOR2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n615), .B(KEYINPUT115), .ZN(n616) );
  XNOR2_X1 U686 ( .A(KEYINPUT116), .B(KEYINPUT53), .ZN(n617) );
  INV_X1 U687 ( .A(n619), .ZN(n621) );
  XNOR2_X1 U688 ( .A(KEYINPUT66), .B(KEYINPUT118), .ZN(n627) );
  XNOR2_X1 U689 ( .A(n629), .B(n628), .ZN(G60) );
  NAND2_X1 U690 ( .A1(n676), .A2(G472), .ZN(n634) );
  XOR2_X1 U691 ( .A(n630), .B(KEYINPUT87), .Z(n632) );
  INV_X1 U692 ( .A(KEYINPUT62), .ZN(n631) );
  XNOR2_X1 U693 ( .A(n634), .B(n633), .ZN(n635) );
  INV_X1 U694 ( .A(KEYINPUT88), .ZN(n636) );
  XNOR2_X1 U695 ( .A(n638), .B(n637), .ZN(G57) );
  XOR2_X1 U696 ( .A(G101), .B(n639), .Z(G3) );
  NAND2_X1 U697 ( .A1(n641), .A2(n653), .ZN(n640) );
  XNOR2_X1 U698 ( .A(n640), .B(G104), .ZN(G6) );
  XNOR2_X1 U699 ( .A(G107), .B(KEYINPUT110), .ZN(n645) );
  XOR2_X1 U700 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n643) );
  NAND2_X1 U701 ( .A1(n641), .A2(n655), .ZN(n642) );
  XNOR2_X1 U702 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U703 ( .A(n645), .B(n644), .ZN(G9) );
  XOR2_X1 U704 ( .A(G110), .B(n646), .Z(G12) );
  XOR2_X1 U705 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n648) );
  NAND2_X1 U706 ( .A1(n651), .A2(n655), .ZN(n647) );
  XNOR2_X1 U707 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U708 ( .A(G143), .B(n650), .ZN(G45) );
  NAND2_X1 U709 ( .A1(n651), .A2(n653), .ZN(n652) );
  XNOR2_X1 U710 ( .A(n652), .B(G146), .ZN(G48) );
  NAND2_X1 U711 ( .A1(n656), .A2(n653), .ZN(n654) );
  XNOR2_X1 U712 ( .A(n654), .B(G113), .ZN(G15) );
  NAND2_X1 U713 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U714 ( .A(n657), .B(G116), .ZN(G18) );
  XOR2_X1 U715 ( .A(KEYINPUT37), .B(KEYINPUT112), .Z(n658) );
  XNOR2_X1 U716 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U717 ( .A(G125), .B(n660), .ZN(G27) );
  XNOR2_X1 U718 ( .A(G134), .B(n703), .ZN(G36) );
  XOR2_X1 U719 ( .A(G140), .B(n661), .Z(G42) );
  NAND2_X1 U720 ( .A1(n676), .A2(G210), .ZN(n664) );
  NOR2_X2 U721 ( .A1(n680), .A2(n665), .ZN(n666) );
  XNOR2_X1 U722 ( .A(KEYINPUT56), .B(n666), .ZN(G51) );
  XNOR2_X1 U723 ( .A(KEYINPUT58), .B(KEYINPUT117), .ZN(n669) );
  XNOR2_X1 U724 ( .A(n667), .B(KEYINPUT57), .ZN(n668) );
  XNOR2_X1 U725 ( .A(n669), .B(n668), .ZN(n671) );
  NAND2_X1 U726 ( .A1(n676), .A2(G469), .ZN(n670) );
  XNOR2_X1 U727 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U728 ( .A1(n680), .A2(n672), .ZN(G54) );
  NAND2_X1 U729 ( .A1(G478), .A2(n676), .ZN(n673) );
  XNOR2_X1 U730 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U731 ( .A1(n680), .A2(n675), .ZN(G63) );
  NAND2_X1 U732 ( .A1(G217), .A2(n676), .ZN(n677) );
  XNOR2_X1 U733 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X1 U734 ( .A1(n680), .A2(n679), .ZN(G66) );
  XOR2_X1 U735 ( .A(KEYINPUT119), .B(KEYINPUT61), .Z(n682) );
  NAND2_X1 U736 ( .A1(G224), .A2(G953), .ZN(n681) );
  XNOR2_X1 U737 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U738 ( .A1(G898), .A2(n683), .ZN(n684) );
  XNOR2_X1 U739 ( .A(n684), .B(KEYINPUT120), .ZN(n687) );
  NAND2_X1 U740 ( .A1(n685), .A2(n707), .ZN(n686) );
  NAND2_X1 U741 ( .A1(n687), .A2(n686), .ZN(n694) );
  XNOR2_X1 U742 ( .A(n688), .B(G101), .ZN(n690) );
  NOR2_X1 U743 ( .A1(n707), .A2(G898), .ZN(n689) );
  NOR2_X1 U744 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U745 ( .A(n691), .B(KEYINPUT121), .Z(n692) );
  XNOR2_X1 U746 ( .A(KEYINPUT122), .B(n692), .ZN(n693) );
  XNOR2_X1 U747 ( .A(n694), .B(n693), .ZN(G69) );
  XOR2_X1 U748 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n698) );
  XNOR2_X1 U749 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U750 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U751 ( .A(n700), .B(n699), .ZN(n706) );
  XNOR2_X1 U752 ( .A(G227), .B(n706), .ZN(n701) );
  NAND2_X1 U753 ( .A1(G900), .A2(n701), .ZN(n702) );
  NAND2_X1 U754 ( .A1(n702), .A2(G953), .ZN(n710) );
  NAND2_X1 U755 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U756 ( .A(n706), .B(n705), .ZN(n708) );
  NAND2_X1 U757 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U758 ( .A1(n710), .A2(n709), .ZN(G72) );
  XOR2_X1 U759 ( .A(G131), .B(KEYINPUT126), .Z(n711) );
  XNOR2_X1 U760 ( .A(n712), .B(n711), .ZN(G33) );
  XNOR2_X1 U761 ( .A(G122), .B(n713), .ZN(n714) );
  XNOR2_X1 U762 ( .A(n714), .B(KEYINPUT125), .ZN(G24) );
  XOR2_X1 U763 ( .A(n715), .B(G119), .Z(G21) );
  XOR2_X1 U764 ( .A(G137), .B(n716), .Z(G39) );
endmodule

