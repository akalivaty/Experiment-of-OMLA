//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149, new_n1150;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n464), .B2(G101), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n459), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n459), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n488), .A3(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n460), .B2(new_n461), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n492), .B(new_n495), .C1(new_n461), .C2(new_n460), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n490), .B1(new_n494), .B2(new_n496), .ZN(G164));
  NAND2_X1  g072(.A1(KEYINPUT67), .A2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(KEYINPUT67), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n505), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  INV_X1    g090(.A(G51), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n502), .A2(new_n506), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n517), .B1(G89), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT68), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  AOI22_X1  g098(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n504), .ZN(new_n525));
  INV_X1    g100(.A(G90), .ZN(new_n526));
  INV_X1    g101(.A(G52), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n507), .A2(new_n526), .B1(new_n509), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G171));
  AOI22_X1  g104(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n504), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT69), .B(G81), .ZN(new_n532));
  INV_X1    g107(.A(G43), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n507), .A2(new_n532), .B1(new_n509), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n535));
  OR3_X1    g110(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n531), .B2(new_n534), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  NAND4_X1  g115(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND4_X1  g118(.A1(G319), .A2(G483), .A3(G661), .A4(new_n543), .ZN(G188));
  NAND3_X1  g119(.A1(new_n506), .A2(G53), .A3(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT9), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT9), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n506), .A2(new_n547), .A3(G53), .A4(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G65), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n500), .B2(new_n501), .ZN(new_n551));
  AND2_X1   g126(.A1(G78), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n502), .A2(G91), .A3(new_n506), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(G299));
  INV_X1    g130(.A(G171), .ZN(G301));
  NAND2_X1  g131(.A1(new_n518), .A2(G87), .ZN(new_n557));
  INV_X1    g132(.A(new_n509), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G49), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(G288));
  NAND2_X1  g136(.A1(new_n518), .A2(G86), .ZN(new_n562));
  AND2_X1   g137(.A1(KEYINPUT6), .A2(G651), .ZN(new_n563));
  NOR2_X1   g138(.A1(KEYINPUT6), .A2(G651), .ZN(new_n564));
  OAI211_X1 g139(.A(G48), .B(G543), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT71), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n506), .A2(KEYINPUT71), .A3(G48), .A4(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G61), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n500), .B2(new_n501), .ZN(new_n571));
  AND2_X1   g146(.A1(G73), .A2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n562), .A2(new_n569), .A3(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n504), .ZN(new_n576));
  INV_X1    g151(.A(G85), .ZN(new_n577));
  INV_X1    g152(.A(G47), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n507), .A2(new_n577), .B1(new_n509), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n504), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(new_n584), .B2(new_n583), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n518), .A2(KEYINPUT10), .A3(G92), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n507), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n587), .A2(new_n590), .B1(G54), .B2(new_n558), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G321));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G299), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(G168), .B2(new_n595), .ZN(G297));
  XOR2_X1   g172(.A(G297), .B(KEYINPUT73), .Z(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n538), .A2(new_n595), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n586), .A2(new_n591), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n603), .B2(new_n595), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n474), .A2(new_n464), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(G2100), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT74), .Z(new_n611));
  NAND2_X1  g186(.A1(new_n476), .A2(G135), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n479), .A2(G123), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n459), .A2(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2096), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n609), .B2(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n611), .A2(new_n618), .ZN(G156));
  INV_X1    g194(.A(KEYINPUT14), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(new_n622), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n625), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G14), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n630), .A2(new_n631), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(G401));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2072), .B(G2078), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT75), .Z(new_n638));
  INV_X1    g213(.A(KEYINPUT76), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2084), .B(G2090), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n638), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n636), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n641), .B(new_n642), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n642), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n638), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT18), .Z(new_n649));
  NOR2_X1   g224(.A1(new_n636), .A2(new_n642), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n646), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2096), .B(G2100), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  XOR2_X1   g231(.A(G1956), .B(G2474), .Z(new_n657));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  AND2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT78), .B(KEYINPUT20), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n658), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  MUX2_X1   g239(.A(new_n664), .B(new_n663), .S(new_n656), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G1981), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G1986), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT79), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  NOR2_X1   g248(.A1(G29), .A2(G33), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT25), .Z(new_n676));
  INV_X1    g251(.A(G139), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(new_n677), .B2(new_n475), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n474), .A2(G127), .ZN(new_n679));
  INV_X1    g254(.A(G115), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n463), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n678), .B1(G2105), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n674), .B1(new_n682), .B2(G29), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT88), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(G2072), .Z(new_n685));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G35), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G162), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT29), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(G2090), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G19), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n539), .B2(new_n692), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT84), .B(G1341), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n690), .A2(new_n691), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n685), .B(new_n696), .C1(new_n694), .C2(new_n695), .ZN(new_n697));
  NOR2_X1   g272(.A1(G168), .A2(new_n692), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n692), .B2(G21), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT89), .B(G1966), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT90), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n692), .A2(G20), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT23), .ZN(new_n704));
  INV_X1    g279(.A(G299), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n692), .ZN(new_n706));
  INV_X1    g281(.A(G1956), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n690), .B2(new_n691), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n697), .A2(new_n702), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G4), .A2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT83), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n602), .B2(new_n692), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1348), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT31), .B(G11), .Z(new_n715));
  NOR2_X1   g290(.A1(new_n616), .A2(new_n686), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT30), .B(G28), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n715), .B(new_n716), .C1(new_n686), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n686), .A2(G27), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT91), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(KEYINPUT91), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n720), .B(new_n721), .C1(G164), .C2(new_n686), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n718), .B1(G2078), .B2(new_n722), .C1(new_n699), .C2(new_n700), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n692), .A2(G5), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G171), .B2(new_n692), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1961), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n689), .A2(G2090), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n722), .A2(G2078), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n686), .B1(new_n730), .B2(G34), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(G34), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G160), .B2(G29), .ZN(new_n733));
  INV_X1    g308(.A(G2084), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n686), .A2(G32), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n476), .A2(G141), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT26), .Z(new_n741));
  INV_X1    g316(.A(G129), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n478), .B2(new_n742), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n464), .A2(G105), .ZN(new_n744));
  OR3_X1    g319(.A1(new_n739), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n737), .B1(new_n746), .B2(new_n686), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT27), .ZN(new_n748));
  INV_X1    g323(.A(G1996), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n686), .A2(G26), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  OR2_X1    g328(.A1(G104), .A2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT85), .Z(new_n756));
  INV_X1    g331(.A(G128), .ZN(new_n757));
  INV_X1    g332(.A(G140), .ZN(new_n758));
  OAI22_X1  g333(.A1(new_n757), .A2(new_n478), .B1(new_n475), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(KEYINPUT86), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(KEYINPUT86), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n753), .B1(new_n763), .B2(G29), .ZN(new_n764));
  INV_X1    g339(.A(G2067), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n736), .A2(new_n750), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n710), .A2(new_n714), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n692), .A2(G22), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G166), .B2(new_n692), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1971), .ZN(new_n771));
  OR2_X1    g346(.A1(G6), .A2(G16), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G305), .B2(new_n692), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT32), .B(G1981), .Z(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G16), .A2(G23), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT80), .ZN(new_n778));
  NAND2_X1  g353(.A1(G288), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n557), .A2(new_n559), .A3(KEYINPUT80), .A4(new_n560), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n777), .B1(new_n781), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT33), .B(G1976), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n773), .A2(new_n774), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n776), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT34), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n776), .A2(new_n784), .A3(new_n788), .A4(new_n785), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT81), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n686), .A2(G25), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n476), .A2(G131), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n479), .A2(G119), .ZN(new_n793));
  OR2_X1    g368(.A1(G95), .A2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n791), .B1(new_n797), .B2(new_n686), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT35), .B(G1991), .Z(new_n799));
  XOR2_X1   g374(.A(new_n798), .B(new_n799), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n692), .A2(G24), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n580), .B2(new_n692), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1986), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  AND3_X1   g379(.A1(new_n789), .A2(new_n790), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n790), .B1(new_n789), .B2(new_n804), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n787), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(KEYINPUT82), .A2(KEYINPUT36), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n807), .A2(KEYINPUT82), .A3(KEYINPUT36), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n768), .B1(new_n809), .B2(new_n810), .ZN(G311));
  XNOR2_X1  g386(.A(G311), .B(KEYINPUT93), .ZN(G150));
  AOI22_X1  g387(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n504), .ZN(new_n814));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n507), .A2(new_n815), .B1(new_n509), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G860), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT37), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n602), .A2(new_n599), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n818), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n538), .A2(new_n825), .ZN(new_n826));
  OR3_X1    g401(.A1(new_n825), .A2(new_n531), .A3(new_n534), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n824), .B(new_n828), .Z(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n819), .B1(new_n830), .B2(KEYINPUT39), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n821), .B1(new_n831), .B2(new_n832), .ZN(G145));
  XNOR2_X1  g408(.A(new_n763), .B(G164), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n796), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n745), .B(new_n682), .ZN(new_n836));
  AOI22_X1  g411(.A1(G130), .A2(new_n479), .B1(new_n476), .B2(G142), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  OR3_X1    g416(.A1(new_n459), .A2(KEYINPUT95), .A3(G118), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT95), .B1(new_n459), .B2(G118), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n837), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(new_n607), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n836), .B(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n835), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n835), .A2(new_n847), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n616), .B(new_n483), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(G160), .Z(new_n852));
  AOI21_X1  g427(.A(G37), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n848), .A2(new_n849), .ZN(new_n855));
  INV_X1    g430(.A(new_n852), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI211_X1 g432(.A(KEYINPUT97), .B(new_n852), .C1(new_n848), .C2(new_n849), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g435(.A1(new_n825), .A2(new_n595), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n580), .B(KEYINPUT98), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n781), .ZN(new_n863));
  XNOR2_X1  g438(.A(G303), .B(G305), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT99), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n863), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n862), .A2(new_n781), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n862), .A2(new_n781), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n870), .A2(KEYINPUT99), .A3(new_n865), .A4(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT42), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n828), .B(new_n603), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n592), .A2(new_n705), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n602), .A2(G299), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(KEYINPUT41), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(new_n876), .B2(new_n877), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n876), .A2(new_n877), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(new_n875), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n874), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n861), .B1(new_n885), .B2(new_n595), .ZN(G295));
  OAI21_X1  g461(.A(new_n861), .B1(new_n885), .B2(new_n595), .ZN(G331));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n888));
  NAND3_X1  g463(.A1(G168), .A2(KEYINPUT100), .A3(G171), .ZN(new_n889));
  NAND2_X1  g464(.A1(G171), .A2(KEYINPUT100), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n525), .B2(new_n528), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(G286), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n828), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n826), .A2(new_n889), .A3(new_n827), .A4(new_n893), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT102), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n883), .B1(new_n894), .B2(new_n828), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n828), .A2(new_n894), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n898), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n881), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n881), .B2(new_n903), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n873), .B(new_n901), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n873), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n897), .A2(new_n902), .A3(new_n899), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n911), .A2(new_n881), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n900), .A2(new_n898), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n902), .A2(new_n898), .ZN(new_n915));
  INV_X1    g490(.A(new_n880), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n878), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT101), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n881), .A2(new_n903), .A3(new_n904), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n920), .A2(KEYINPUT103), .A3(new_n873), .A4(new_n901), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n909), .A2(new_n914), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT104), .ZN(new_n924));
  AOI21_X1  g499(.A(G37), .B1(new_n907), .B2(new_n908), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n925), .A2(new_n926), .A3(new_n914), .A4(new_n921), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n888), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n920), .A2(new_n901), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n925), .B(new_n921), .C1(new_n873), .C2(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n930), .A2(new_n888), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(KEYINPUT43), .B2(new_n923), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n936), .ZN(G397));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G164), .B2(G1384), .ZN(new_n939));
  INV_X1    g514(.A(new_n472), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n465), .A2(new_n468), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n940), .A2(new_n941), .A3(G40), .A4(new_n462), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n763), .A2(G2067), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n761), .A2(new_n765), .A3(new_n762), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n943), .B1(new_n946), .B2(new_n745), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n749), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT46), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT125), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT47), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n946), .A2(new_n943), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT106), .ZN(new_n954));
  NOR4_X1   g529(.A1(G290), .A2(new_n939), .A3(G1986), .A4(new_n942), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT126), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT48), .Z(new_n957));
  NOR2_X1   g532(.A1(new_n948), .A2(new_n745), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n958), .B(KEYINPUT105), .Z(new_n959));
  NOR2_X1   g534(.A1(new_n746), .A2(new_n749), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n943), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n796), .B(new_n799), .Z(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n943), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n954), .A2(new_n957), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n952), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n954), .A2(new_n961), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n797), .A2(new_n799), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n945), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n965), .B1(new_n943), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n970));
  INV_X1    g545(.A(G40), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n469), .A2(new_n472), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n494), .A2(new_n496), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n485), .A2(new_n489), .ZN(new_n974));
  AOI21_X1  g549(.A(G1384), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR3_X1   g552(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n707), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT57), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n553), .A2(KEYINPUT112), .A3(new_n554), .ZN(new_n981));
  NAND3_X1  g556(.A1(G299), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n553), .A2(new_n554), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n983), .B(new_n549), .C1(KEYINPUT112), .C2(KEYINPUT57), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  INV_X1    g561(.A(new_n496), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n495), .B1(new_n474), .B2(new_n492), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(KEYINPUT45), .B(new_n986), .C1(new_n989), .C2(new_n490), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT56), .B(G2072), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n939), .A2(new_n990), .A3(new_n972), .A4(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n979), .A2(new_n985), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT113), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n979), .A2(new_n985), .A3(new_n995), .A4(new_n992), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n979), .A2(new_n992), .ZN(new_n998));
  INV_X1    g573(.A(new_n985), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT61), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT114), .B(G1996), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n939), .A2(new_n990), .A3(new_n972), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n975), .A2(new_n972), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT58), .B(G1341), .Z(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n539), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT59), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT59), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n539), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1000), .A2(KEYINPUT61), .A3(new_n993), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n970), .B1(new_n1001), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT61), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n998), .B2(new_n999), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n993), .A2(new_n1017), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n994), .A2(new_n996), .B1(new_n999), .B2(new_n998), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1018), .B(KEYINPUT115), .C1(KEYINPUT61), .C2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1004), .A2(G2067), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n986), .B1(new_n989), .B2(new_n490), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n942), .B1(new_n1022), .B2(KEYINPUT50), .ZN(new_n1023));
  NOR4_X1   g598(.A1(G164), .A2(KEYINPUT107), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT107), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n975), .B2(new_n976), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1023), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1348), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1021), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT60), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(new_n592), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n602), .B1(new_n1029), .B2(KEYINPUT60), .ZN(new_n1032));
  OAI22_X1  g607(.A1(new_n1031), .A2(new_n1032), .B1(KEYINPUT60), .B2(new_n1029), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1015), .A2(new_n1020), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1000), .B1(new_n1029), .B2(new_n602), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n997), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1034), .A2(KEYINPUT116), .A3(new_n1036), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1023), .B(new_n734), .C1(new_n1026), .C2(new_n1024), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n939), .A2(new_n972), .A3(new_n990), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n700), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1042), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G286), .A2(G8), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT119), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1041), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(KEYINPUT120), .B(new_n1041), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1047), .A2(new_n1054), .ZN(new_n1055));
  OR3_X1    g630(.A1(new_n1046), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1053), .B1(new_n1046), .B2(new_n1055), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1051), .A2(new_n1052), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1047), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1059));
  XOR2_X1   g634(.A(new_n1059), .B(KEYINPUT117), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1961), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n1063));
  INV_X1    g638(.A(G2078), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n939), .A2(new_n990), .A3(new_n1064), .A4(new_n972), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1027), .A2(new_n1062), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1065), .A2(new_n1063), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1066), .B(new_n1067), .C1(KEYINPUT123), .C2(G301), .ZN(new_n1068));
  AOI21_X1  g643(.A(G301), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT54), .B(new_n1068), .C1(new_n1070), .C2(KEYINPUT123), .ZN(new_n1071));
  INV_X1    g646(.A(G2090), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1023), .B(new_n1072), .C1(new_n1026), .C2(new_n1024), .ZN(new_n1073));
  INV_X1    g648(.A(G1971), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1044), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1042), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G305), .A2(G1981), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT49), .ZN(new_n1083));
  INV_X1    g658(.A(G1981), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n562), .A2(new_n569), .A3(new_n1084), .A4(new_n573), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1083), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1004), .A2(KEYINPUT108), .A3(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT108), .B1(new_n1004), .B2(G8), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n1086), .A2(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n779), .A2(G1976), .A3(new_n780), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT109), .B(G1976), .Z(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(G288), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1091), .B(new_n1093), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1091), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT52), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1081), .A2(new_n1090), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT111), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n975), .A2(new_n976), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1023), .A2(new_n1072), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1042), .B1(new_n1100), .B2(new_n1075), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1098), .B1(new_n1101), .B2(new_n1080), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1079), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(new_n1077), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n977), .A2(new_n978), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1105), .A2(new_n1072), .B1(new_n1074), .B2(new_n1044), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT111), .B(new_n1104), .C1(new_n1106), .C2(new_n1042), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1097), .A2(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1110));
  AND3_X1   g685(.A1(new_n1066), .A2(G301), .A3(new_n1067), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1110), .B1(new_n1111), .B2(new_n1069), .ZN(new_n1112));
  AND4_X1   g687(.A1(new_n1061), .A2(new_n1071), .A3(new_n1109), .A4(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1039), .A2(new_n1040), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT110), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1096), .A2(new_n1090), .A3(new_n1094), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n1081), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1085), .ZN(new_n1118));
  NOR2_X1   g693(.A1(G288), .A2(G1976), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1090), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1115), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  OAI221_X1 g698(.A(KEYINPUT110), .B1(new_n1120), .B2(new_n1121), .C1(new_n1116), .C2(new_n1081), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1046), .A2(G168), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT63), .B1(new_n1109), .B2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1126), .B(KEYINPUT63), .C1(new_n1080), .C2(new_n1076), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(new_n1097), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1125), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1058), .A2(new_n1131), .A3(new_n1060), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1097), .A2(new_n1108), .A3(new_n1070), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1061), .A2(KEYINPUT62), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1130), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1114), .A2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n580), .B(G1986), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n943), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n954), .A2(new_n961), .A3(new_n1139), .A4(new_n963), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT124), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1143), .B(new_n1140), .C1(new_n1114), .C2(new_n1136), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n969), .B1(new_n1142), .B2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g720(.A(G319), .B1(new_n633), .B2(new_n634), .ZN(new_n1147));
  NOR2_X1   g721(.A1(G227), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g722(.A(new_n1148), .B(KEYINPUT127), .ZN(new_n1149));
  NOR2_X1   g723(.A1(G229), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g724(.A1(new_n934), .A2(new_n1150), .A3(new_n859), .ZN(G225));
  INV_X1    g725(.A(G225), .ZN(G308));
endmodule


