//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT2), .B(G113), .Z(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT68), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT2), .B(G113), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT67), .B(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G116), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT66), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n197), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(new_n194), .B2(G119), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n189), .B(new_n192), .C1(new_n201), .C2(KEYINPUT66), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT4), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT79), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n205), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n204), .B1(new_n209), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n199), .A2(new_n202), .B1(new_n203), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n209), .A2(new_n204), .A3(new_n213), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n218), .A2(KEYINPUT4), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n216), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n201), .A2(KEYINPUT5), .ZN(new_n223));
  INV_X1    g037(.A(G113), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT5), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n200), .B2(new_n225), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n223), .A2(new_n226), .B1(new_n201), .B2(new_n188), .ZN(new_n227));
  OAI21_X1  g041(.A(G101), .B1(new_n208), .B2(new_n211), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n218), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n222), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G110), .B(G122), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n233), .B(KEYINPUT84), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n215), .A2(new_n221), .B1(new_n230), .B2(new_n227), .ZN(new_n236));
  INV_X1    g050(.A(new_n234), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(KEYINPUT6), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G143), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  OR2_X1    g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n244), .B1(new_n247), .B2(new_n245), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G125), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n241), .A2(KEYINPUT1), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n244), .A2(new_n252), .A3(G128), .ZN(new_n253));
  INV_X1    g067(.A(G128), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n241), .B(new_n243), .C1(KEYINPUT1), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n257), .A2(KEYINPUT86), .A3(G125), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT86), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n259), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n251), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT87), .B(G224), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(G953), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n262), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT85), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n237), .B1(new_n222), .B2(new_n231), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR4_X1   g083(.A1(new_n236), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n237), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n239), .B(new_n265), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT88), .B(KEYINPUT7), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n262), .B1(new_n264), .B2(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n234), .B(KEYINPUT8), .Z(new_n274));
  INV_X1    g088(.A(new_n231), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n227), .A2(new_n230), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n264), .B(KEYINPUT89), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n278), .A2(KEYINPUT7), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n251), .C1(new_n258), .C2(new_n261), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n273), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n281), .B2(new_n238), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n271), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(G210), .B1(G237), .B2(G902), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n271), .A2(new_n282), .A3(new_n284), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G214), .B1(G237), .B2(G902), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(KEYINPUT83), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(G113), .B(G122), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(new_n210), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT90), .ZN(new_n295));
  INV_X1    g109(.A(G214), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n296), .A2(G237), .A3(G953), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n295), .B1(new_n297), .B2(G143), .ZN(new_n298));
  INV_X1    g112(.A(G237), .ZN(new_n299));
  INV_X1    g113(.A(G953), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(G214), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT90), .A3(new_n242), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n298), .A2(new_n302), .B1(G143), .B2(new_n297), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT18), .A2(G131), .ZN(new_n304));
  XNOR2_X1  g118(.A(G125), .B(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n240), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n305), .A2(new_n240), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n303), .A2(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n298), .A2(new_n302), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n297), .A2(G143), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT18), .A3(G131), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n305), .A2(KEYINPUT16), .ZN(new_n315));
  OR3_X1    g129(.A1(new_n260), .A2(KEYINPUT16), .A3(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(G146), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT19), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n305), .B(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n317), .B1(new_n319), .B2(G146), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n311), .A2(G131), .ZN(new_n321));
  INV_X1    g135(.A(G131), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n303), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n294), .B1(new_n314), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT17), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n321), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n317), .ZN(new_n328));
  AOI21_X1  g142(.A(G146), .B1(new_n315), .B2(new_n316), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n321), .B2(new_n326), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n293), .B(new_n313), .C1(new_n327), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT91), .ZN(new_n334));
  NOR2_X1   g148(.A1(G475), .A2(G902), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT91), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n325), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT20), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT20), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n325), .B2(new_n332), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n313), .B1(new_n327), .B2(new_n331), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n294), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n332), .ZN(new_n346));
  INV_X1    g160(.A(G902), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n339), .A2(new_n343), .B1(G475), .B2(new_n348), .ZN(new_n349));
  XOR2_X1   g163(.A(KEYINPUT73), .B(G902), .Z(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n194), .A2(G122), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n353));
  AND2_X1   g167(.A1(KEYINPUT92), .A2(G122), .ZN(new_n354));
  NOR2_X1   g168(.A1(KEYINPUT92), .A2(G122), .ZN(new_n355));
  OAI21_X1  g169(.A(G116), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n352), .B2(KEYINPUT14), .ZN(new_n357));
  OAI21_X1  g171(.A(G107), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(KEYINPUT64), .A2(G134), .ZN(new_n359));
  NOR2_X1   g173(.A1(KEYINPUT64), .A2(G134), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n242), .A2(G128), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n254), .A2(G143), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n363), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT64), .B(G134), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n367), .A3(KEYINPUT93), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n352), .A2(new_n206), .A3(new_n356), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n364), .A2(new_n367), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n358), .B(new_n370), .C1(KEYINPUT93), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n363), .A2(KEYINPUT13), .ZN(new_n373));
  MUX2_X1   g187(.A(KEYINPUT13), .B(new_n373), .S(new_n362), .Z(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G134), .ZN(new_n375));
  INV_X1    g189(.A(new_n369), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n206), .B1(new_n352), .B2(new_n356), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n375), .B(new_n364), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(KEYINPUT9), .B(G234), .Z(new_n380));
  XOR2_X1   g194(.A(KEYINPUT74), .B(G217), .Z(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n300), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT94), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n383), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n372), .A2(new_n385), .A3(new_n378), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n351), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G478), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(KEYINPUT15), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n386), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n385), .B1(new_n372), .B2(new_n378), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n350), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT15), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G478), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT95), .B(G952), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(G953), .ZN(new_n396));
  NAND2_X1  g210(.A1(G234), .A2(G237), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n351), .A2(G953), .A3(new_n397), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT21), .B(G898), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n389), .A2(new_n394), .A3(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n288), .A2(new_n291), .A3(new_n349), .A4(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n230), .A2(new_n405), .A3(KEYINPUT10), .A4(new_n257), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n218), .A2(new_n255), .A3(new_n253), .A4(new_n228), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT81), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n214), .A2(new_n203), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n411), .A2(new_n249), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n221), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n407), .A2(new_n408), .ZN(new_n414));
  INV_X1    g228(.A(G137), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n415), .A2(KEYINPUT11), .A3(G134), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(new_n361), .B2(G137), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n359), .B2(new_n360), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT11), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n420), .A3(new_n322), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT65), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n417), .A2(new_n420), .A3(KEYINPUT65), .A4(new_n322), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n420), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n423), .A2(new_n424), .B1(G131), .B2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n410), .A2(new_n413), .A3(new_n414), .A4(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT12), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n426), .B2(KEYINPUT82), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n424), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(G131), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n229), .A2(new_n256), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n430), .A2(new_n431), .B1(new_n407), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n429), .A2(new_n433), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n427), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G140), .ZN(new_n438));
  INV_X1    g252(.A(G227), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(G953), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n438), .B(new_n440), .Z(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n410), .A2(new_n413), .A3(new_n414), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n430), .A2(new_n431), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n427), .A3(new_n441), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n443), .A2(G469), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(G469), .A2(G902), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n427), .A3(new_n442), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT12), .B1(new_n445), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n433), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n410), .A2(new_n413), .A3(new_n414), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n454), .A2(new_n434), .B1(new_n455), .B2(new_n426), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n450), .B(new_n350), .C1(new_n456), .C2(new_n442), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n448), .B(new_n449), .C1(G469), .C2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G221), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n380), .B2(new_n347), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n187), .B1(new_n404), .B2(new_n462), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n271), .A2(new_n284), .A3(new_n282), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n284), .B1(new_n271), .B2(new_n282), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n291), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n348), .A2(G475), .ZN(new_n467));
  INV_X1    g281(.A(new_n337), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n336), .B1(new_n325), .B2(new_n332), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n340), .B1(new_n470), .B2(new_n335), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n467), .B(new_n403), .C1(new_n471), .C2(new_n342), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n458), .A2(new_n461), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT96), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n445), .A2(new_n249), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n199), .A2(new_n202), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n415), .A2(G134), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n366), .B2(new_n415), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n255), .B(new_n253), .C1(new_n481), .C2(new_n322), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n430), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n477), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT28), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT71), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n250), .B1(new_n430), .B2(new_n431), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n482), .B1(new_n423), .B2(new_n424), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n488), .B(new_n478), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n484), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n490), .A2(KEYINPUT69), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n494), .A2(new_n477), .A3(new_n479), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n488), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n477), .A2(new_n484), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n478), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n492), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n487), .B1(new_n500), .B2(new_n486), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n299), .A2(new_n300), .A3(G210), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n502), .B(KEYINPUT27), .Z(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT26), .B(G101), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n503), .B(new_n504), .Z(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n490), .A2(KEYINPUT69), .ZN(new_n510));
  AOI211_X1 g324(.A(new_n493), .B(new_n482), .C1(new_n423), .C2(new_n424), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n510), .A2(new_n489), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n509), .B1(new_n512), .B2(KEYINPUT30), .ZN(new_n513));
  OAI22_X1  g327(.A1(new_n426), .A2(new_n250), .B1(new_n490), .B2(KEYINPUT69), .ZN(new_n514));
  NOR4_X1   g328(.A1(new_n514), .A2(KEYINPUT70), .A3(new_n507), .A4(new_n511), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n478), .B(new_n508), .C1(new_n513), .C2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n505), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n496), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT29), .B1(new_n506), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n478), .B1(new_n514), .B2(new_n511), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n496), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n521), .A2(KEYINPUT28), .B1(KEYINPUT72), .B2(new_n487), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT72), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n523), .B(new_n486), .C1(new_n520), .C2(new_n496), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT29), .A3(new_n505), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n350), .ZN(new_n527));
  OAI21_X1  g341(.A(G472), .B1(new_n519), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(G472), .A2(G902), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n516), .A2(new_n496), .A3(new_n505), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n531), .A2(KEYINPUT31), .B1(new_n501), .B2(new_n517), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n516), .A2(new_n533), .A3(new_n496), .A4(new_n505), .ZN(new_n534));
  AOI211_X1 g348(.A(KEYINPUT32), .B(new_n530), .C1(new_n532), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT32), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(KEYINPUT31), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n501), .A2(new_n517), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n539), .B2(new_n529), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n528), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT22), .B(G137), .Z(new_n542));
  INV_X1    g356(.A(G234), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n459), .A2(new_n543), .A3(G953), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n542), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT76), .B(KEYINPUT23), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n254), .A2(G119), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n254), .A2(KEYINPUT23), .A3(G119), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n549), .A2(KEYINPUT75), .B1(new_n196), .B2(G128), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT77), .ZN(new_n553));
  OR3_X1    g367(.A1(new_n552), .A2(new_n553), .A3(G110), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n553), .B1(new_n552), .B2(G110), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n196), .A2(G128), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n547), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT24), .B(G110), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n317), .A2(new_n306), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n557), .A2(new_n558), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n330), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n552), .A2(G110), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n560), .A2(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n545), .B1(new_n566), .B2(KEYINPUT78), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(KEYINPUT78), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n569), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n567), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n350), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT25), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n381), .B1(new_n351), .B2(new_n543), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n351), .B1(new_n570), .B2(new_n572), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n576), .A2(new_n347), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n575), .A2(new_n579), .B1(new_n580), .B2(new_n573), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n476), .A2(new_n541), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  NAND2_X1  g397(.A1(new_n539), .A2(new_n350), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G472), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n539), .A2(new_n529), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n289), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n286), .B2(new_n287), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n402), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n467), .B1(new_n471), .B2(new_n342), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n387), .A2(new_n388), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT97), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n595), .B(KEYINPUT33), .C1(new_n390), .C2(new_n391), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n595), .A2(KEYINPUT33), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(KEYINPUT33), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n384), .A2(new_n386), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n351), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n594), .B1(new_n600), .B2(new_n388), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT98), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n594), .B(new_n603), .C1(new_n600), .C2(new_n388), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n593), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n592), .A2(KEYINPUT99), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n591), .B2(new_n605), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n581), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n462), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n588), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  NAND3_X1  g429(.A1(new_n612), .A2(new_n586), .A3(new_n585), .ZN(new_n616));
  INV_X1    g430(.A(new_n470), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n339), .B1(new_n617), .B2(new_n341), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n389), .A2(new_n394), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n618), .A2(new_n619), .A3(new_n467), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n592), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT35), .B(G107), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  NAND2_X1  g438(.A1(new_n575), .A2(new_n579), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n545), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n566), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n580), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n463), .A2(new_n475), .A3(new_n630), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n631), .A2(new_n587), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT100), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  OAI21_X1  g449(.A(new_n398), .B1(new_n399), .B2(G900), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n590), .A2(new_n630), .A3(new_n620), .A4(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n541), .A2(new_n474), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G128), .ZN(G30));
  INV_X1    g453(.A(new_n629), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n575), .B2(new_n579), .ZN(new_n641));
  INV_X1    g455(.A(new_n619), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n349), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n641), .A2(new_n289), .A3(new_n643), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n644), .A2(KEYINPUT101), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(KEYINPUT101), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n288), .B(KEYINPUT38), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n636), .B(KEYINPUT39), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n474), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT40), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n521), .A2(new_n517), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n531), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(G472), .B1(new_n653), .B2(G902), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n654), .B1(new_n535), .B2(new_n540), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n648), .A2(new_n651), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n242), .ZN(G45));
  NAND4_X1  g472(.A1(new_n593), .A2(new_n602), .A3(new_n604), .A4(new_n636), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n289), .B1(new_n464), .B2(new_n465), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n659), .A2(new_n641), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n541), .A2(new_n474), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G146), .ZN(G48));
  NAND2_X1  g477(.A1(KEYINPUT102), .A2(G469), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n457), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n437), .A2(new_n441), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n667), .A2(new_n450), .A3(new_n350), .A4(new_n664), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n461), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT103), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n610), .A2(new_n541), .A3(new_n581), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT104), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  INV_X1    g488(.A(new_n621), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n541), .A2(new_n581), .A3(new_n675), .A4(new_n670), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G116), .ZN(G18));
  AND3_X1   g491(.A1(new_n666), .A2(new_n461), .A3(new_n668), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n590), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT105), .B1(new_n660), .B2(new_n669), .ZN(new_n681));
  AOI211_X1 g495(.A(new_n472), .B(new_n641), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT106), .B1(new_n682), .B2(new_n541), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(KEYINPUT106), .A3(new_n541), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G119), .ZN(G21));
  OAI21_X1  g501(.A(new_n517), .B1(new_n522), .B2(new_n524), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n537), .A2(new_n534), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n529), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n585), .A2(new_n581), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n643), .A2(new_n590), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n670), .A2(new_n693), .A3(new_n402), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G122), .ZN(G24));
  INV_X1    g510(.A(new_n659), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n679), .B1(new_n590), .B2(new_n678), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n660), .A2(new_n669), .A3(KEYINPUT105), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n351), .B1(new_n532), .B2(new_n534), .ZN(new_n701));
  INV_X1    g515(.A(G472), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n690), .B(new_n630), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n260), .ZN(G27));
  NOR2_X1   g519(.A1(new_n288), .A2(new_n589), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n461), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n447), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n447), .A2(new_n708), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n709), .A2(new_n443), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n457), .A2(G469), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n712), .A2(new_n713), .A3(new_n449), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n707), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n541), .A2(new_n581), .A3(new_n697), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT42), .ZN(new_n718));
  AOI21_X1  g532(.A(KEYINPUT42), .B1(new_n716), .B2(new_n717), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G131), .ZN(G33));
  AND2_X1   g535(.A1(new_n620), .A2(new_n636), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n541), .A2(new_n581), .A3(new_n722), .A4(new_n715), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G134), .ZN(G36));
  NAND3_X1  g538(.A1(new_n349), .A2(new_n602), .A3(new_n604), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g541(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n727), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT111), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n587), .A3(new_n630), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n443), .A2(new_n447), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n711), .A2(KEYINPUT45), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(G469), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n449), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n735), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n739), .A2(KEYINPUT109), .A3(KEYINPUT46), .A4(new_n449), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n741), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n742), .A2(new_n713), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n745), .A2(new_n461), .A3(new_n649), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n733), .A2(new_n706), .A3(new_n734), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G137), .ZN(G39));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n461), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n706), .ZN(new_n752));
  OR4_X1    g566(.A1(new_n581), .A2(new_n541), .A3(new_n659), .A4(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G140), .ZN(G42));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n641), .A2(new_n461), .A3(new_n636), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n758), .A2(new_n714), .A3(new_n692), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n655), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n662), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n586), .A2(KEYINPUT32), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n539), .A2(new_n536), .A3(new_n529), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n462), .B1(new_n764), .B2(new_n528), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n704), .B1(new_n765), .B2(new_n637), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n761), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n703), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n659), .B1(new_n680), .B2(new_n681), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n638), .A2(new_n662), .A3(new_n771), .A4(new_n760), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT114), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n768), .A2(KEYINPUT52), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(new_n768), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n769), .A2(new_n697), .A3(new_n715), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n642), .A2(new_n467), .A3(new_n636), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n618), .A2(new_n630), .A3(new_n706), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n541), .A2(new_n474), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n723), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n718), .A2(new_n719), .A3(new_n781), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n476), .A2(new_n541), .A3(new_n581), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n605), .B1(new_n593), .B2(new_n642), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n288), .A2(new_n291), .A3(new_n402), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OAI22_X1  g601(.A1(new_n616), .A2(new_n787), .B1(new_n631), .B2(new_n587), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT112), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n616), .A2(new_n787), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(new_n632), .A3(new_n791), .A4(new_n582), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n685), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n683), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n671), .A2(new_n695), .A3(new_n676), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n782), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n757), .B1(new_n776), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n757), .B1(new_n789), .B2(new_n792), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n671), .A2(new_n695), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n686), .A2(new_n801), .A3(new_n802), .A4(new_n676), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT116), .B1(new_n795), .B2(new_n796), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n782), .A2(new_n800), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n768), .A2(new_n773), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n638), .A2(new_n771), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT113), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n638), .A2(new_n771), .A3(new_n811), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n810), .A2(new_n812), .B1(new_n765), .B2(new_n661), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n807), .B1(new_n655), .B2(new_n759), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n808), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n805), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n799), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n798), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT53), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n768), .A2(new_n773), .A3(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n808), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n820), .A3(KEYINPUT53), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n823), .A2(KEYINPUT115), .A3(new_n820), .A4(KEYINPUT53), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n821), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n819), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n729), .A2(new_n398), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n581), .A3(new_n585), .A4(new_n690), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n680), .A2(new_n681), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n666), .A2(new_n668), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n707), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n611), .A2(new_n398), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n656), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI221_X1 g652(.A(new_n396), .B1(new_n832), .B2(new_n834), .C1(new_n605), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n831), .A2(new_n836), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT118), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n541), .A2(new_n581), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n844), .B(KEYINPUT48), .Z(new_n845));
  NOR2_X1   g659(.A1(new_n832), .A2(new_n752), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n835), .A2(new_n461), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n751), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT51), .B1(new_n848), .B2(KEYINPUT119), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n832), .A2(new_n289), .A3(new_n647), .A4(new_n669), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT50), .ZN(new_n851));
  INV_X1    g665(.A(new_n838), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n593), .B1(new_n602), .B2(new_n604), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n841), .A2(new_n769), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n848), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n839), .B(new_n845), .C1(new_n849), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(new_n849), .B2(new_n855), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n830), .A2(new_n857), .B1(G952), .B2(G953), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n581), .A2(new_n461), .A3(new_n291), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n835), .B(KEYINPUT49), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n647), .A2(new_n859), .A3(new_n860), .A4(new_n725), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n656), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n858), .A2(new_n862), .ZN(G75));
  NOR2_X1   g677(.A1(new_n300), .A2(G952), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n239), .B1(new_n269), .B2(new_n270), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(new_n265), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT55), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT53), .B1(new_n823), .B2(new_n820), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n806), .A2(new_n807), .B1(new_n813), .B2(new_n814), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n800), .A2(new_n803), .A3(new_n804), .A4(new_n782), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n351), .B(new_n285), .C1(new_n868), .C2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT56), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n867), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n351), .B1(new_n868), .B2(new_n871), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT120), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n877), .B(new_n351), .C1(new_n868), .C2(new_n871), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n285), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n867), .A2(new_n873), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n864), .B(new_n874), .C1(new_n879), .C2(new_n880), .ZN(G51));
  XOR2_X1   g695(.A(new_n449), .B(KEYINPUT57), .Z(new_n882));
  INV_X1    g696(.A(new_n818), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n868), .A2(new_n871), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n818), .B1(new_n799), .B2(new_n817), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n667), .A3(new_n450), .ZN(new_n887));
  INV_X1    g701(.A(new_n739), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n876), .A2(new_n888), .A3(new_n878), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n864), .B1(new_n887), .B2(new_n889), .ZN(G54));
  NAND2_X1  g704(.A1(KEYINPUT58), .A2(G475), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT121), .Z(new_n892));
  NAND3_X1  g706(.A1(new_n876), .A2(new_n878), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n617), .ZN(new_n894));
  INV_X1    g708(.A(new_n864), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n876), .A2(new_n470), .A3(new_n878), .A4(new_n892), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G60));
  NAND2_X1  g711(.A1(new_n596), .A2(new_n599), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT59), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n830), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n899), .A2(new_n901), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n883), .B1(new_n868), .B2(new_n871), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(new_n819), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n904), .B1(new_n908), .B2(new_n864), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n905), .B1(new_n884), .B2(new_n885), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(KEYINPUT122), .A3(new_n895), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n899), .A2(new_n903), .B1(new_n909), .B2(new_n911), .ZN(G63));
  XOR2_X1   g726(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n913));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT60), .Z(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n799), .B2(new_n817), .ZN(new_n917));
  OAI211_X1 g731(.A(KEYINPUT124), .B(new_n895), .C1(new_n917), .C2(new_n573), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n628), .B(new_n915), .C1(new_n868), .C2(new_n871), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n915), .B1(new_n868), .B2(new_n871), .ZN(new_n921));
  INV_X1    g735(.A(new_n573), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT124), .B1(new_n923), .B2(new_n895), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n913), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n895), .B1(new_n917), .B2(new_n573), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n864), .B1(new_n921), .B2(new_n922), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n930), .A2(KEYINPUT125), .A3(KEYINPUT61), .A4(new_n919), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n925), .A2(new_n932), .ZN(G66));
  NAND2_X1  g747(.A1(new_n793), .A2(new_n797), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n300), .ZN(new_n935));
  OAI21_X1  g749(.A(G953), .B1(new_n263), .B2(new_n400), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n865), .B1(G898), .B2(new_n300), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  NOR2_X1   g753(.A1(new_n513), .A2(new_n515), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n507), .B2(new_n498), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n319), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n746), .A2(new_n843), .A3(new_n693), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n755), .A2(new_n723), .A3(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n720), .A3(new_n747), .A4(new_n813), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n300), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n439), .A2(G900), .A3(G953), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n942), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n657), .B1(new_n950), .B2(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n813), .A2(new_n951), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n952), .A2(new_n950), .A3(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n784), .A2(new_n706), .ZN(new_n954));
  OR3_X1    g768(.A1(new_n842), .A2(new_n650), .A3(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n747), .A2(new_n755), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n952), .B1(new_n950), .B2(KEYINPUT62), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n953), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n949), .B1(new_n958), .B2(G953), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n948), .B1(new_n959), .B2(new_n942), .ZN(G72));
  XNOR2_X1  g774(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n702), .A2(new_n347), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n961), .B(new_n962), .Z(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n958), .B2(new_n934), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n517), .B1(new_n516), .B2(new_n496), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n964), .B1(new_n945), .B2(new_n934), .ZN(new_n968));
  INV_X1    g782(.A(new_n518), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(new_n895), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n828), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n969), .A2(new_n966), .A3(new_n963), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G57));
endmodule


