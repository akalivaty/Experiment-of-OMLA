

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U555 ( .A(n633), .Z(n634) );
  NOR2_X1 U556 ( .A1(n557), .A2(G2104), .ZN(n558) );
  NOR2_X2 U557 ( .A1(n786), .A2(n787), .ZN(n726) );
  NOR2_X1 U558 ( .A1(n714), .A2(n715), .ZN(n703) );
  NAND2_X1 U559 ( .A1(n696), .A2(n695), .ZN(n786) );
  XNOR2_X1 U560 ( .A(KEYINPUT89), .B(n821), .ZN(n521) );
  AND2_X1 U561 ( .A1(n561), .A2(n560), .ZN(n522) );
  NOR2_X1 U562 ( .A1(n952), .A2(KEYINPUT33), .ZN(n523) );
  AND2_X1 U563 ( .A1(n771), .A2(n770), .ZN(n524) );
  AND2_X1 U564 ( .A1(n701), .A2(n700), .ZN(n525) );
  INV_X1 U565 ( .A(n927), .ZN(n702) );
  NAND2_X1 U566 ( .A1(n525), .A2(n702), .ZN(n714) );
  NOR2_X1 U567 ( .A1(n736), .A2(n735), .ZN(n737) );
  INV_X1 U568 ( .A(KEYINPUT101), .ZN(n741) );
  AND2_X1 U569 ( .A1(n523), .A2(n760), .ZN(n761) );
  INV_X1 U570 ( .A(n694), .ZN(n696) );
  NAND2_X1 U571 ( .A1(n658), .A2(G66), .ZN(n604) );
  NAND2_X1 U572 ( .A1(n822), .A2(n521), .ZN(n823) );
  NOR2_X1 U573 ( .A1(G543), .A2(n530), .ZN(n531) );
  INV_X1 U574 ( .A(G651), .ZN(n530) );
  INV_X1 U575 ( .A(G2105), .ZN(n557) );
  NOR2_X1 U576 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U577 ( .A(KEYINPUT73), .B(KEYINPUT15), .ZN(n608) );
  AND2_X1 U578 ( .A1(n557), .A2(G2104), .ZN(n901) );
  XNOR2_X1 U579 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n552) );
  XNOR2_X1 U580 ( .A(n609), .B(n608), .ZN(n944) );
  NOR2_X1 U581 ( .A1(G651), .A2(n647), .ZN(n656) );
  XNOR2_X1 U582 ( .A(n553), .B(n552), .ZN(n555) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n657) );
  NAND2_X1 U584 ( .A1(n657), .A2(G89), .ZN(n526) );
  XNOR2_X1 U585 ( .A(n526), .B(KEYINPUT4), .ZN(n528) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n647) );
  NOR2_X1 U587 ( .A1(n647), .A2(n530), .ZN(n661) );
  NAND2_X1 U588 ( .A1(G76), .A2(n661), .ZN(n527) );
  NAND2_X1 U589 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U590 ( .A(n529), .B(KEYINPUT5), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n656), .A2(G51), .ZN(n534) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n531), .Z(n532) );
  XNOR2_X2 U593 ( .A(n532), .B(KEYINPUT66), .ZN(n658) );
  NAND2_X1 U594 ( .A1(G63), .A2(n658), .ZN(n533) );
  NAND2_X1 U595 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U596 ( .A(KEYINPUT6), .B(n535), .Z(n536) );
  NAND2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U598 ( .A(n538), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U599 ( .A(G168), .B(KEYINPUT8), .Z(n539) );
  XNOR2_X1 U600 ( .A(KEYINPUT74), .B(n539), .ZN(G286) );
  NAND2_X1 U601 ( .A1(G85), .A2(n657), .ZN(n541) );
  NAND2_X1 U602 ( .A1(G60), .A2(n658), .ZN(n540) );
  NAND2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n545) );
  NAND2_X1 U604 ( .A1(G72), .A2(n661), .ZN(n543) );
  NAND2_X1 U605 ( .A1(G47), .A2(n656), .ZN(n542) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U607 ( .A1(n545), .A2(n544), .ZN(G290) );
  NAND2_X1 U608 ( .A1(G88), .A2(n657), .ZN(n547) );
  NAND2_X1 U609 ( .A1(G75), .A2(n661), .ZN(n546) );
  NAND2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n656), .A2(G50), .ZN(n549) );
  NAND2_X1 U612 ( .A1(G62), .A2(n658), .ZN(n548) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U614 ( .A1(n551), .A2(n550), .ZN(G166) );
  INV_X1 U615 ( .A(G166), .ZN(G303) );
  NAND2_X1 U616 ( .A1(G101), .A2(n901), .ZN(n553) );
  AND2_X1 U617 ( .A1(G2104), .A2(G2105), .ZN(n896) );
  NAND2_X1 U618 ( .A1(G113), .A2(n896), .ZN(n554) );
  AND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n698) );
  NOR2_X1 U620 ( .A1(G2104), .A2(G2105), .ZN(n556) );
  XOR2_X1 U621 ( .A(KEYINPUT17), .B(n556), .Z(n633) );
  NAND2_X1 U622 ( .A1(n633), .A2(G137), .ZN(n561) );
  XNOR2_X1 U623 ( .A(n558), .B(KEYINPUT64), .ZN(n572) );
  INV_X1 U624 ( .A(n572), .ZN(n559) );
  INV_X1 U625 ( .A(n559), .ZN(n897) );
  NAND2_X1 U626 ( .A1(G125), .A2(n897), .ZN(n560) );
  AND2_X1 U627 ( .A1(n698), .A2(n522), .ZN(G160) );
  XOR2_X1 U628 ( .A(G2438), .B(G2454), .Z(n563) );
  XNOR2_X1 U629 ( .A(G2435), .B(G2430), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U631 ( .A(n564), .B(G2427), .Z(n566) );
  XNOR2_X1 U632 ( .A(G1348), .B(G1341), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n570) );
  XOR2_X1 U634 ( .A(G2443), .B(G2446), .Z(n568) );
  XNOR2_X1 U635 ( .A(KEYINPUT106), .B(G2451), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U637 ( .A(n570), .B(n569), .Z(n571) );
  AND2_X1 U638 ( .A1(G14), .A2(n571), .ZN(G401) );
  NAND2_X1 U639 ( .A1(n572), .A2(G126), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G114), .A2(n896), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n575), .B(KEYINPUT86), .ZN(n579) );
  NAND2_X1 U643 ( .A1(G102), .A2(n901), .ZN(n577) );
  NAND2_X1 U644 ( .A1(G138), .A2(n633), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n581) );
  INV_X1 U647 ( .A(KEYINPUT87), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n581), .B(n580), .ZN(n694) );
  BUF_X1 U649 ( .A(n694), .Z(G164) );
  NAND2_X1 U650 ( .A1(n656), .A2(G52), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G64), .A2(n658), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G90), .A2(n657), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G77), .A2(n661), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U656 ( .A(KEYINPUT9), .B(n586), .Z(n587) );
  NOR2_X1 U657 ( .A1(n588), .A2(n587), .ZN(G171) );
  AND2_X1 U658 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U659 ( .A(G57), .ZN(G237) );
  INV_X1 U660 ( .A(G132), .ZN(G219) );
  INV_X1 U661 ( .A(G82), .ZN(G220) );
  NAND2_X1 U662 ( .A1(G7), .A2(G661), .ZN(n589) );
  XOR2_X1 U663 ( .A(n589), .B(KEYINPUT10), .Z(n842) );
  NAND2_X1 U664 ( .A1(n842), .A2(G567), .ZN(n590) );
  XOR2_X1 U665 ( .A(KEYINPUT11), .B(n590), .Z(G234) );
  INV_X1 U666 ( .A(G860), .ZN(n850) );
  NAND2_X1 U667 ( .A1(n657), .A2(G81), .ZN(n591) );
  XNOR2_X1 U668 ( .A(n591), .B(KEYINPUT12), .ZN(n593) );
  NAND2_X1 U669 ( .A1(G68), .A2(n661), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n595) );
  XOR2_X1 U671 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n594) );
  XNOR2_X1 U672 ( .A(n595), .B(n594), .ZN(n598) );
  NAND2_X1 U673 ( .A1(G56), .A2(n658), .ZN(n596) );
  XOR2_X1 U674 ( .A(KEYINPUT14), .B(n596), .Z(n597) );
  NOR2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n656), .A2(G43), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n927) );
  NOR2_X1 U678 ( .A1(n850), .A2(n927), .ZN(n601) );
  XNOR2_X1 U679 ( .A(n601), .B(KEYINPUT71), .ZN(G153) );
  XOR2_X1 U680 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U681 ( .A1(G868), .A2(G301), .ZN(n611) );
  NAND2_X1 U682 ( .A1(G92), .A2(n657), .ZN(n603) );
  NAND2_X1 U683 ( .A1(G79), .A2(n661), .ZN(n602) );
  NAND2_X1 U684 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n656), .A2(G54), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n609) );
  INV_X1 U688 ( .A(n944), .ZN(n715) );
  INV_X1 U689 ( .A(G868), .ZN(n674) );
  NAND2_X1 U690 ( .A1(n715), .A2(n674), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(G284) );
  NAND2_X1 U692 ( .A1(n656), .A2(G53), .ZN(n613) );
  NAND2_X1 U693 ( .A1(G65), .A2(n658), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U695 ( .A(KEYINPUT69), .B(n614), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G91), .A2(n657), .ZN(n615) );
  XNOR2_X1 U697 ( .A(n615), .B(KEYINPUT67), .ZN(n618) );
  NAND2_X1 U698 ( .A1(G78), .A2(n661), .ZN(n616) );
  XOR2_X1 U699 ( .A(KEYINPUT68), .B(n616), .Z(n617) );
  NOR2_X1 U700 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(G299) );
  NOR2_X1 U702 ( .A1(G286), .A2(n674), .ZN(n621) );
  XOR2_X1 U703 ( .A(KEYINPUT75), .B(n621), .Z(n623) );
  NOR2_X1 U704 ( .A1(G868), .A2(G299), .ZN(n622) );
  NOR2_X1 U705 ( .A1(n623), .A2(n622), .ZN(G297) );
  NAND2_X1 U706 ( .A1(n850), .A2(G559), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n624), .A2(n944), .ZN(n625) );
  XNOR2_X1 U708 ( .A(n625), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U709 ( .A1(n715), .A2(n674), .ZN(n626) );
  XOR2_X1 U710 ( .A(KEYINPUT76), .B(n626), .Z(n627) );
  NOR2_X1 U711 ( .A1(G559), .A2(n627), .ZN(n629) );
  NOR2_X1 U712 ( .A1(G868), .A2(n927), .ZN(n628) );
  NOR2_X1 U713 ( .A1(n629), .A2(n628), .ZN(G282) );
  NAND2_X1 U714 ( .A1(G111), .A2(n896), .ZN(n631) );
  NAND2_X1 U715 ( .A1(G99), .A2(n901), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n631), .A2(n630), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G123), .A2(n897), .ZN(n632) );
  XNOR2_X1 U718 ( .A(n632), .B(KEYINPUT18), .ZN(n636) );
  NAND2_X1 U719 ( .A1(G135), .A2(n634), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n1005) );
  XNOR2_X1 U722 ( .A(G2096), .B(n1005), .ZN(n639) );
  INV_X1 U723 ( .A(G2100), .ZN(n860) );
  NAND2_X1 U724 ( .A1(n639), .A2(n860), .ZN(G156) );
  NAND2_X1 U725 ( .A1(G86), .A2(n657), .ZN(n641) );
  NAND2_X1 U726 ( .A1(G61), .A2(n658), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n661), .A2(G73), .ZN(n642) );
  XOR2_X1 U729 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n656), .A2(G48), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U733 ( .A1(G87), .A2(n647), .ZN(n649) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n648) );
  NAND2_X1 U735 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U736 ( .A1(n658), .A2(n650), .ZN(n652) );
  NAND2_X1 U737 ( .A1(n656), .A2(G49), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U739 ( .A1(G559), .A2(n944), .ZN(n653) );
  XOR2_X1 U740 ( .A(n927), .B(n653), .Z(n849) );
  XNOR2_X1 U741 ( .A(KEYINPUT19), .B(KEYINPUT80), .ZN(n655) );
  XNOR2_X1 U742 ( .A(G288), .B(KEYINPUT79), .ZN(n654) );
  XNOR2_X1 U743 ( .A(n655), .B(n654), .ZN(n671) );
  NAND2_X1 U744 ( .A1(G55), .A2(n656), .ZN(n666) );
  NAND2_X1 U745 ( .A1(G93), .A2(n657), .ZN(n660) );
  NAND2_X1 U746 ( .A1(G67), .A2(n658), .ZN(n659) );
  NAND2_X1 U747 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U748 ( .A1(G80), .A2(n661), .ZN(n662) );
  XNOR2_X1 U749 ( .A(KEYINPUT77), .B(n662), .ZN(n663) );
  NOR2_X1 U750 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U751 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U752 ( .A(n667), .B(KEYINPUT78), .ZN(n851) );
  XOR2_X1 U753 ( .A(G299), .B(n851), .Z(n669) );
  XOR2_X1 U754 ( .A(G290), .B(G303), .Z(n668) );
  XNOR2_X1 U755 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U756 ( .A(n671), .B(n670), .Z(n672) );
  XNOR2_X1 U757 ( .A(G305), .B(n672), .ZN(n916) );
  XNOR2_X1 U758 ( .A(n849), .B(n916), .ZN(n673) );
  NOR2_X1 U759 ( .A1(n674), .A2(n673), .ZN(n676) );
  NOR2_X1 U760 ( .A1(n851), .A2(G868), .ZN(n675) );
  NOR2_X1 U761 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U762 ( .A(KEYINPUT81), .B(n677), .Z(G295) );
  NAND2_X1 U763 ( .A1(G2084), .A2(G2078), .ZN(n679) );
  XOR2_X1 U764 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n678) );
  XNOR2_X1 U765 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U766 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U767 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U768 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XOR2_X1 U769 ( .A(KEYINPUT83), .B(G44), .Z(n683) );
  XNOR2_X1 U770 ( .A(KEYINPUT3), .B(n683), .ZN(G218) );
  NOR2_X1 U771 ( .A1(G220), .A2(G219), .ZN(n684) );
  XNOR2_X1 U772 ( .A(KEYINPUT22), .B(n684), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n685), .A2(G96), .ZN(n686) );
  NOR2_X1 U774 ( .A1(G218), .A2(n686), .ZN(n687) );
  XOR2_X1 U775 ( .A(KEYINPUT84), .B(n687), .Z(n854) );
  NAND2_X1 U776 ( .A1(n854), .A2(G2106), .ZN(n691) );
  NAND2_X1 U777 ( .A1(G69), .A2(G120), .ZN(n688) );
  NOR2_X1 U778 ( .A1(G237), .A2(n688), .ZN(n689) );
  NAND2_X1 U779 ( .A1(G108), .A2(n689), .ZN(n853) );
  NAND2_X1 U780 ( .A1(G567), .A2(n853), .ZN(n690) );
  NAND2_X1 U781 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U782 ( .A(KEYINPUT85), .B(n692), .Z(n848) );
  NAND2_X1 U783 ( .A1(G661), .A2(G483), .ZN(n693) );
  NOR2_X1 U784 ( .A1(n848), .A2(n693), .ZN(n847) );
  NAND2_X1 U785 ( .A1(n847), .A2(G36), .ZN(G176) );
  INV_X1 U786 ( .A(G1384), .ZN(n695) );
  AND2_X1 U787 ( .A1(G40), .A2(n522), .ZN(n697) );
  NAND2_X1 U788 ( .A1(n698), .A2(n697), .ZN(n787) );
  NAND2_X1 U789 ( .A1(n726), .A2(G1996), .ZN(n699) );
  XNOR2_X1 U790 ( .A(n699), .B(KEYINPUT26), .ZN(n701) );
  INV_X2 U791 ( .A(n726), .ZN(n743) );
  NAND2_X1 U792 ( .A1(G1341), .A2(n743), .ZN(n700) );
  XNOR2_X1 U793 ( .A(KEYINPUT98), .B(n703), .ZN(n712) );
  NOR2_X1 U794 ( .A1(n726), .A2(G1348), .ZN(n705) );
  NOR2_X1 U795 ( .A1(G2067), .A2(n743), .ZN(n704) );
  NOR2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n710) );
  INV_X1 U797 ( .A(G299), .ZN(n928) );
  NAND2_X1 U798 ( .A1(n726), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U799 ( .A(KEYINPUT27), .B(n706), .ZN(n709) );
  NAND2_X1 U800 ( .A1(G1956), .A2(n743), .ZN(n707) );
  XNOR2_X1 U801 ( .A(KEYINPUT97), .B(n707), .ZN(n708) );
  NOR2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n721) );
  NAND2_X1 U803 ( .A1(n928), .A2(n721), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n710), .A2(n713), .ZN(n711) );
  NOR2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n719) );
  INV_X1 U806 ( .A(n713), .ZN(n717) );
  NAND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U808 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U810 ( .A(n720), .B(KEYINPUT99), .ZN(n724) );
  OR2_X1 U811 ( .A1(n928), .A2(n721), .ZN(n722) );
  XOR2_X1 U812 ( .A(KEYINPUT28), .B(n722), .Z(n723) );
  NOR2_X1 U813 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U814 ( .A(n725), .B(KEYINPUT29), .ZN(n730) );
  INV_X1 U815 ( .A(G1961), .ZN(n931) );
  NAND2_X1 U816 ( .A1(n743), .A2(n931), .ZN(n728) );
  XNOR2_X1 U817 ( .A(KEYINPUT25), .B(G2078), .ZN(n985) );
  NAND2_X1 U818 ( .A1(n726), .A2(n985), .ZN(n727) );
  NAND2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n734) );
  NAND2_X1 U820 ( .A1(G171), .A2(n734), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n730), .A2(n729), .ZN(n740) );
  NAND2_X1 U822 ( .A1(G8), .A2(n743), .ZN(n782) );
  NOR2_X1 U823 ( .A1(G1966), .A2(n782), .ZN(n754) );
  NOR2_X1 U824 ( .A1(G2084), .A2(n743), .ZN(n751) );
  NOR2_X1 U825 ( .A1(n754), .A2(n751), .ZN(n731) );
  NAND2_X1 U826 ( .A1(G8), .A2(n731), .ZN(n732) );
  XNOR2_X1 U827 ( .A(KEYINPUT30), .B(n732), .ZN(n733) );
  NOR2_X1 U828 ( .A1(G168), .A2(n733), .ZN(n736) );
  NOR2_X1 U829 ( .A1(G171), .A2(n734), .ZN(n735) );
  XOR2_X1 U830 ( .A(n737), .B(KEYINPUT31), .Z(n738) );
  XNOR2_X1 U831 ( .A(n738), .B(KEYINPUT100), .ZN(n739) );
  NAND2_X1 U832 ( .A1(n740), .A2(n739), .ZN(n752) );
  NAND2_X1 U833 ( .A1(n752), .A2(G286), .ZN(n742) );
  XNOR2_X1 U834 ( .A(n742), .B(n741), .ZN(n748) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n782), .ZN(n745) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n743), .ZN(n744) );
  NOR2_X1 U837 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U838 ( .A1(G303), .A2(n746), .ZN(n747) );
  NAND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U840 ( .A1(n749), .A2(G8), .ZN(n750) );
  XNOR2_X1 U841 ( .A(n750), .B(KEYINPUT32), .ZN(n758) );
  NAND2_X1 U842 ( .A1(G8), .A2(n751), .ZN(n756) );
  INV_X1 U843 ( .A(n752), .ZN(n753) );
  NOR2_X1 U844 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n775) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n952) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n759) );
  XNOR2_X1 U849 ( .A(KEYINPUT102), .B(n759), .ZN(n935) );
  INV_X1 U850 ( .A(n935), .ZN(n760) );
  NAND2_X1 U851 ( .A1(n775), .A2(n761), .ZN(n772) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n765) );
  NAND2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n945) );
  INV_X1 U854 ( .A(n945), .ZN(n762) );
  OR2_X1 U855 ( .A1(n762), .A2(n782), .ZN(n763) );
  OR2_X1 U856 ( .A1(KEYINPUT103), .A2(n763), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n771) );
  XOR2_X1 U858 ( .A(n935), .B(KEYINPUT103), .Z(n766) );
  NAND2_X1 U859 ( .A1(n766), .A2(KEYINPUT33), .ZN(n767) );
  NOR2_X1 U860 ( .A1(n782), .A2(n767), .ZN(n769) );
  XOR2_X1 U861 ( .A(G1981), .B(G305), .Z(n939) );
  INV_X1 U862 ( .A(n939), .ZN(n768) );
  NOR2_X1 U863 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U864 ( .A1(n772), .A2(n524), .ZN(n778) );
  NOR2_X1 U865 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U866 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U867 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n776), .A2(n782), .ZN(n777) );
  NAND2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U870 ( .A(KEYINPUT104), .B(n779), .ZN(n785) );
  NOR2_X1 U871 ( .A1(G1981), .A2(G305), .ZN(n780) );
  XOR2_X1 U872 ( .A(n780), .B(KEYINPUT24), .Z(n781) );
  NOR2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U874 ( .A(n783), .B(KEYINPUT96), .ZN(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n824) );
  INV_X1 U876 ( .A(n786), .ZN(n788) );
  NOR2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U878 ( .A(KEYINPUT88), .B(n789), .ZN(n836) );
  XOR2_X1 U879 ( .A(KEYINPUT95), .B(n836), .Z(n808) );
  NAND2_X1 U880 ( .A1(G105), .A2(n901), .ZN(n790) );
  XNOR2_X1 U881 ( .A(n790), .B(KEYINPUT38), .ZN(n797) );
  NAND2_X1 U882 ( .A1(G117), .A2(n896), .ZN(n792) );
  NAND2_X1 U883 ( .A1(G129), .A2(n897), .ZN(n791) );
  NAND2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G141), .A2(n634), .ZN(n793) );
  XNOR2_X1 U886 ( .A(KEYINPUT93), .B(n793), .ZN(n794) );
  NOR2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U889 ( .A(KEYINPUT94), .B(n798), .ZN(n910) );
  NAND2_X1 U890 ( .A1(G1996), .A2(n910), .ZN(n807) );
  NAND2_X1 U891 ( .A1(n901), .A2(G95), .ZN(n800) );
  NAND2_X1 U892 ( .A1(G119), .A2(n897), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n896), .A2(G107), .ZN(n801) );
  XOR2_X1 U895 ( .A(KEYINPUT92), .B(n801), .Z(n802) );
  NOR2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n634), .A2(G131), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n882) );
  NAND2_X1 U899 ( .A1(G1991), .A2(n882), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n1010) );
  NAND2_X1 U901 ( .A1(n808), .A2(n1010), .ZN(n826) );
  INV_X1 U902 ( .A(n836), .ZN(n820) );
  XNOR2_X1 U903 ( .A(G2067), .B(KEYINPUT37), .ZN(n834) );
  NAND2_X1 U904 ( .A1(n901), .A2(G104), .ZN(n809) );
  XNOR2_X1 U905 ( .A(n809), .B(KEYINPUT90), .ZN(n811) );
  NAND2_X1 U906 ( .A1(G140), .A2(n634), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U908 ( .A(KEYINPUT34), .B(n812), .ZN(n817) );
  NAND2_X1 U909 ( .A1(G116), .A2(n896), .ZN(n814) );
  NAND2_X1 U910 ( .A1(G128), .A2(n897), .ZN(n813) );
  NAND2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U912 ( .A(KEYINPUT35), .B(n815), .Z(n816) );
  NOR2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U914 ( .A(n818), .B(KEYINPUT91), .ZN(n819) );
  XOR2_X1 U915 ( .A(n819), .B(KEYINPUT36), .Z(n913) );
  OR2_X1 U916 ( .A1(n834), .A2(n913), .ZN(n1011) );
  OR2_X1 U917 ( .A1(n820), .A2(n1011), .ZN(n832) );
  AND2_X1 U918 ( .A1(n826), .A2(n832), .ZN(n822) );
  XOR2_X1 U919 ( .A(G1986), .B(G290), .Z(n946) );
  NOR2_X1 U920 ( .A1(n820), .A2(n946), .ZN(n821) );
  XNOR2_X1 U921 ( .A(n825), .B(KEYINPUT105), .ZN(n839) );
  NOR2_X1 U922 ( .A1(G1996), .A2(n910), .ZN(n1015) );
  INV_X1 U923 ( .A(n826), .ZN(n829) );
  NOR2_X1 U924 ( .A1(G1986), .A2(G290), .ZN(n827) );
  NOR2_X1 U925 ( .A1(G1991), .A2(n882), .ZN(n1006) );
  NOR2_X1 U926 ( .A1(n827), .A2(n1006), .ZN(n828) );
  NOR2_X1 U927 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U928 ( .A1(n1015), .A2(n830), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n831), .B(KEYINPUT39), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n833), .A2(n832), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n834), .A2(n913), .ZN(n1017) );
  NAND2_X1 U932 ( .A1(n835), .A2(n1017), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U935 ( .A(n840), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U936 ( .A1(n842), .A2(G2106), .ZN(n841) );
  XOR2_X1 U937 ( .A(KEYINPUT107), .B(n841), .Z(G217) );
  INV_X1 U938 ( .A(n842), .ZN(G223) );
  NAND2_X1 U939 ( .A1(G15), .A2(G2), .ZN(n843) );
  XOR2_X1 U940 ( .A(KEYINPUT108), .B(n843), .Z(n844) );
  NAND2_X1 U941 ( .A1(n844), .A2(G661), .ZN(n845) );
  XOR2_X1 U942 ( .A(KEYINPUT109), .B(n845), .Z(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U944 ( .A1(n847), .A2(n846), .ZN(G188) );
  INV_X1 U945 ( .A(n848), .ZN(G319) );
  NAND2_X1 U947 ( .A1(n850), .A2(n849), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n852), .B(n851), .ZN(G145) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  INV_X1 U951 ( .A(G69), .ZN(G235) );
  NOR2_X1 U952 ( .A1(n854), .A2(n853), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  XOR2_X1 U954 ( .A(G2096), .B(G2678), .Z(n856) );
  XNOR2_X1 U955 ( .A(G2090), .B(KEYINPUT43), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U957 ( .A(n857), .B(KEYINPUT42), .Z(n859) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n864) );
  XNOR2_X1 U960 ( .A(KEYINPUT110), .B(n860), .ZN(n862) );
  XNOR2_X1 U961 ( .A(G2084), .B(G2078), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(G227) );
  XOR2_X1 U964 ( .A(G1976), .B(G1971), .Z(n866) );
  XNOR2_X1 U965 ( .A(G1986), .B(G1956), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U967 ( .A(n867), .B(KEYINPUT41), .Z(n869) );
  XNOR2_X1 U968 ( .A(G1966), .B(G1981), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n873) );
  XNOR2_X1 U970 ( .A(G2474), .B(n931), .ZN(n871) );
  XNOR2_X1 U971 ( .A(G1996), .B(G1991), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(G229) );
  NAND2_X1 U974 ( .A1(G100), .A2(n901), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G136), .A2(n634), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n897), .A2(G124), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n876), .B(KEYINPUT44), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G112), .A2(n896), .ZN(n877) );
  XOR2_X1 U980 ( .A(KEYINPUT111), .B(n877), .Z(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U982 ( .A1(n881), .A2(n880), .ZN(G162) );
  XNOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n882), .B(G162), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n895) );
  NAND2_X1 U986 ( .A1(G118), .A2(n896), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G130), .A2(n897), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n893) );
  NAND2_X1 U989 ( .A1(n901), .A2(G106), .ZN(n887) );
  XNOR2_X1 U990 ( .A(n887), .B(KEYINPUT112), .ZN(n889) );
  NAND2_X1 U991 ( .A1(G142), .A2(n634), .ZN(n888) );
  NAND2_X1 U992 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U993 ( .A(KEYINPUT45), .B(n890), .ZN(n891) );
  XNOR2_X1 U994 ( .A(KEYINPUT113), .B(n891), .ZN(n892) );
  NOR2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U996 ( .A(n895), .B(n894), .Z(n908) );
  NAND2_X1 U997 ( .A1(G115), .A2(n896), .ZN(n899) );
  NAND2_X1 U998 ( .A1(G127), .A2(n897), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n900), .B(KEYINPUT47), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(G103), .A2(n901), .ZN(n902) );
  NAND2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n634), .A2(G139), .ZN(n904) );
  XOR2_X1 U1004 ( .A(KEYINPUT114), .B(n904), .Z(n905) );
  NOR2_X1 U1005 ( .A1(n906), .A2(n905), .ZN(n1022) );
  XNOR2_X1 U1006 ( .A(G164), .B(n1022), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1008 ( .A(n909), .B(n1005), .Z(n912) );
  XNOR2_X1 U1009 ( .A(G160), .B(n910), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n915), .ZN(G395) );
  XNOR2_X1 U1013 ( .A(n916), .B(n927), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n917), .B(G286), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n944), .B(G171), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n920), .ZN(n921) );
  XOR2_X1 U1018 ( .A(KEYINPUT115), .B(n921), .Z(G397) );
  NOR2_X1 U1019 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(G401), .A2(n923), .ZN(n924) );
  AND2_X1 U1022 ( .A1(G319), .A2(n924), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G108), .ZN(G238) );
  INV_X1 U1027 ( .A(G16), .ZN(n978) );
  XNOR2_X1 U1028 ( .A(KEYINPUT56), .B(n978), .ZN(n954) );
  XNOR2_X1 U1029 ( .A(n927), .B(G1341), .ZN(n930) );
  XOR2_X1 U1030 ( .A(n928), .B(G1956), .Z(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n937) );
  XOR2_X1 U1032 ( .A(n931), .B(G171), .Z(n933) );
  NAND2_X1 U1033 ( .A1(G1971), .A2(G303), .ZN(n932) );
  NAND2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n943) );
  XOR2_X1 U1037 ( .A(G1966), .B(G168), .Z(n938) );
  XNOR2_X1 U1038 ( .A(KEYINPUT123), .B(n938), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1040 ( .A(KEYINPUT57), .B(n941), .Z(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n950) );
  XOR2_X1 U1042 ( .A(G1348), .B(n944), .Z(n948) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n1034) );
  XOR2_X1 U1048 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n961) );
  XNOR2_X1 U1049 ( .A(G1986), .B(G24), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G23), .B(G1976), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G1971), .B(KEYINPUT125), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(G22), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n961), .B(n960), .ZN(n974) );
  XOR2_X1 U1056 ( .A(G1348), .B(KEYINPUT59), .Z(n962) );
  XNOR2_X1 U1057 ( .A(G4), .B(n962), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(G20), .B(G1956), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(G1341), .B(G19), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(G1981), .B(G6), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n969), .B(KEYINPUT60), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(G1961), .B(KEYINPUT124), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(G5), .B(n970), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(G21), .B(G1966), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(KEYINPUT61), .B(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n980), .A2(G11), .ZN(n1004) );
  XNOR2_X1 U1074 ( .A(KEYINPUT119), .B(G2090), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(n981), .B(G35), .ZN(n996) );
  XNOR2_X1 U1076 ( .A(G2067), .B(G26), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(G33), .B(G2072), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n992) );
  XOR2_X1 U1079 ( .A(G1991), .B(G25), .Z(n984) );
  NAND2_X1 U1080 ( .A1(n984), .A2(G28), .ZN(n990) );
  XOR2_X1 U1081 ( .A(G1996), .B(G32), .Z(n987) );
  XNOR2_X1 U1082 ( .A(n985), .B(G27), .ZN(n986) );
  NAND2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1084 ( .A(KEYINPUT120), .B(n988), .ZN(n989) );
  NOR2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1087 ( .A(KEYINPUT53), .B(n993), .ZN(n994) );
  XOR2_X1 U1088 ( .A(KEYINPUT121), .B(n994), .Z(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(G34), .B(G2084), .ZN(n997) );
  XNOR2_X1 U1091 ( .A(KEYINPUT54), .B(n997), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(KEYINPUT122), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1001), .A2(G29), .ZN(n1002) );
  XOR2_X1 U1095 ( .A(KEYINPUT55), .B(n1002), .Z(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1032) );
  XNOR2_X1 U1097 ( .A(G160), .B(G2084), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT116), .B(n1013), .ZN(n1020) );
  XOR2_X1 U1103 ( .A(G2090), .B(G162), .Z(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1105 ( .A(KEYINPUT51), .B(n1016), .Z(n1018) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1108 ( .A(KEYINPUT117), .B(n1021), .Z(n1028) );
  XOR2_X1 U1109 ( .A(G2072), .B(n1022), .Z(n1023) );
  XNOR2_X1 U1110 ( .A(KEYINPUT118), .B(n1023), .ZN(n1025) );
  XOR2_X1 U1111 ( .A(G164), .B(G2078), .Z(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(KEYINPUT50), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1115 ( .A(KEYINPUT52), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1116 ( .A1(n1030), .A2(G29), .ZN(n1031) );
  NAND2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1118 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1119 ( .A(KEYINPUT127), .B(n1035), .Z(n1036) );
  XOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1036), .Z(G150) );
  INV_X1 U1121 ( .A(G150), .ZN(G311) );
endmodule

