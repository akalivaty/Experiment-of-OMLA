//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n212), .A2(G1), .A3(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n206), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n209), .B(new_n221), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n245), .B(new_n251), .ZN(G351));
  NAND2_X1  g0052(.A1(new_n216), .A2(G33), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT68), .ZN(new_n254));
  XOR2_X1   g0054(.A(KEYINPUT8), .B(G58), .Z(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT67), .B1(new_n206), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT67), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n262), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n215), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n259), .A2(new_n265), .B1(new_n202), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n215), .A2(new_n264), .A3(new_n267), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(G20), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(G50), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT9), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n276), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n278), .B1(new_n282), .B2(G226), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n283), .A2(KEYINPUT66), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G222), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(G223), .A3(G1698), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n287), .B(new_n288), .C1(new_n223), .C2(new_n285), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n214), .A2(new_n279), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n283), .A2(KEYINPUT66), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n284), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n293), .A2(G200), .B1(KEYINPUT71), .B2(KEYINPUT10), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n275), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT71), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n299), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n275), .A2(new_n295), .A3(new_n296), .A4(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n293), .A2(G179), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n293), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n274), .A3(new_n305), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n300), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G97), .ZN(new_n308));
  INV_X1    g0108(.A(G232), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G1698), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(G226), .B2(G1698), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT3), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G33), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n308), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n290), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n278), .B1(new_n282), .B2(G238), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n304), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT14), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(G179), .A3(new_n321), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n322), .B2(new_n323), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT70), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n270), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n215), .A2(new_n264), .A3(KEYINPUT70), .A4(new_n267), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n329), .A2(new_n330), .A3(new_n272), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G68), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n214), .B1(new_n261), .B2(new_n263), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n254), .A2(G77), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n247), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n336), .A2(KEYINPUT11), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(KEYINPUT11), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n268), .A2(new_n247), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT12), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n332), .A2(new_n337), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n327), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n320), .A2(G190), .A3(new_n321), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT72), .ZN(new_n344));
  INV_X1    g0144(.A(G200), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n320), .B2(new_n321), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n255), .ZN(new_n349));
  INV_X1    g0149(.A(new_n257), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT15), .B(G87), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n352), .A2(new_n253), .B1(new_n216), .B2(new_n223), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n265), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT69), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(new_n223), .B2(new_n268), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n331), .A2(G77), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n278), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G232), .A2(G1698), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n286), .A2(G238), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n285), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G107), .B2(new_n285), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n214), .A2(new_n279), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n359), .B1(new_n224), .B2(new_n281), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(G179), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n304), .B2(new_n365), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n358), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n365), .A2(new_n294), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(G200), .B2(new_n365), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n356), .A2(new_n357), .A3(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n307), .A2(new_n342), .A3(new_n348), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT77), .ZN(new_n374));
  MUX2_X1   g0174(.A(G223), .B(G226), .S(G1698), .Z(new_n375));
  NAND2_X1  g0175(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT3), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n378), .A3(G33), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n375), .A2(new_n379), .A3(new_n312), .ZN(new_n380));
  INV_X1    g0180(.A(G87), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n260), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n290), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n278), .B1(new_n282), .B2(G232), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n304), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n364), .B1(new_n380), .B2(new_n383), .ZN(new_n388));
  INV_X1    g0188(.A(G179), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n359), .B1(new_n281), .B2(new_n309), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n374), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(G169), .B1(new_n388), .B2(new_n390), .ZN(new_n393));
  INV_X1    g0193(.A(new_n312), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(G33), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n382), .B1(new_n396), .B2(new_n375), .ZN(new_n397));
  OAI211_X1 g0197(.A(G179), .B(new_n386), .C1(new_n397), .C2(new_n364), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n398), .A3(KEYINPUT77), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n255), .A2(new_n272), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n271), .A2(new_n401), .B1(new_n268), .B2(new_n349), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  AND3_X1   g0203(.A1(KEYINPUT74), .A2(G58), .A3(G68), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT74), .B1(G58), .B2(G68), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n216), .B1(new_n406), .B2(new_n218), .ZN(new_n407));
  INV_X1    g0207(.A(G159), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n350), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n314), .B1(new_n395), .B2(G33), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT7), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(G20), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n315), .A2(new_n216), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n411), .A2(new_n413), .B1(new_n414), .B2(new_n412), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n410), .B1(new_n415), .B2(new_n247), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n333), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT75), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n407), .B2(new_n409), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n404), .A2(new_n405), .A3(new_n201), .ZN(new_n421));
  OAI221_X1 g0221(.A(KEYINPUT75), .B1(new_n408), .B2(new_n350), .C1(new_n421), .C2(new_n216), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT7), .B1(new_n396), .B2(G20), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n379), .A2(new_n312), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(new_n412), .A3(new_n216), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(G68), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n427), .A3(KEYINPUT16), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n403), .B1(new_n418), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n400), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT18), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n416), .A2(new_n417), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n432), .A3(new_n265), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT78), .ZN(new_n434));
  AOI21_X1  g0234(.A(G200), .B1(new_n385), .B2(new_n386), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n388), .A2(G190), .A3(new_n390), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n385), .A2(new_n294), .A3(new_n386), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n345), .B1(new_n388), .B2(new_n390), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(KEYINPUT78), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n433), .A2(new_n437), .A3(new_n440), .A4(new_n402), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n373), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(G257), .A2(G1698), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n226), .B2(G1698), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n379), .A3(new_n312), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n315), .A2(G303), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n364), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G41), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n266), .B(G45), .C1(new_n450), .C2(KEYINPUT5), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT79), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(KEYINPUT5), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n451), .B2(KEYINPUT79), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n280), .A2(G274), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n449), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(G270), .B(new_n280), .C1(new_n453), .C2(new_n455), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n345), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT20), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  INV_X1    g0262(.A(G97), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n216), .C1(G33), .C2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G20), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n461), .B1(new_n333), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n265), .A2(KEYINPUT20), .A3(new_n464), .A4(new_n466), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n465), .B1(new_n266), .B2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n329), .A2(new_n330), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n268), .A2(new_n465), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT80), .B1(new_n460), .B2(new_n474), .ZN(new_n475));
  OR2_X1    g0275(.A1(new_n451), .A2(KEYINPUT79), .ZN(new_n476));
  INV_X1    g0276(.A(new_n456), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n452), .A4(new_n454), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n447), .A2(new_n448), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n459), .B(new_n478), .C1(new_n479), .C2(new_n364), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G200), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT80), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n468), .A2(new_n469), .B1(new_n465), .B2(new_n268), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n472), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n458), .A2(G190), .A3(new_n459), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n475), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n304), .B1(new_n458), .B2(new_n459), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n474), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT21), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n480), .A2(new_n389), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n488), .A2(new_n489), .B1(new_n474), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(new_n474), .A3(KEYINPUT21), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n486), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G264), .B(new_n280), .C1(new_n453), .C2(new_n455), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G250), .A2(G1698), .ZN(new_n496));
  INV_X1    g0296(.A(G257), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(G1698), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n396), .A2(new_n498), .B1(G33), .B2(G294), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n495), .B(new_n478), .C1(new_n499), .C2(new_n364), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n345), .ZN(new_n501));
  INV_X1    g0301(.A(new_n498), .ZN(new_n502));
  INV_X1    g0302(.A(G294), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n425), .A2(new_n502), .B1(new_n260), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n290), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(new_n294), .A3(new_n478), .A4(new_n495), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT22), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(new_n381), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n379), .A2(new_n216), .A3(new_n312), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n216), .A2(G87), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n508), .B1(new_n315), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G116), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G20), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT23), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n216), .B2(G107), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n225), .A2(KEYINPUT23), .A3(G20), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n510), .A2(new_n512), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT24), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT24), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n510), .A2(new_n512), .A3(new_n521), .A4(new_n518), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n333), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n267), .A2(G107), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT25), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n266), .A2(G33), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n333), .A2(new_n267), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n525), .B1(new_n527), .B2(new_n225), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n507), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n500), .A2(new_n304), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n505), .A2(new_n389), .A3(new_n478), .A4(new_n495), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(new_n532), .C1(new_n523), .C2(new_n528), .ZN(new_n533));
  INV_X1    g0333(.A(new_n280), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n266), .A2(G45), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G250), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n534), .A2(new_n536), .B1(new_n277), .B2(new_n535), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(G238), .A2(G1698), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n224), .B2(G1698), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n396), .A2(new_n540), .B1(G33), .B2(G116), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(new_n364), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n304), .ZN(new_n543));
  NOR2_X1   g0343(.A1(G97), .A2(G107), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(new_n381), .B1(new_n308), .B2(new_n216), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G97), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n545), .A2(new_n546), .B1(new_n253), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n379), .A2(new_n216), .A3(G68), .A4(new_n312), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(new_n265), .B1(new_n268), .B2(new_n352), .ZN(new_n551));
  INV_X1    g0351(.A(new_n352), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n271), .A2(new_n526), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n540), .A2(new_n379), .A3(new_n312), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n364), .B1(new_n555), .B2(new_n513), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n537), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n389), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n543), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(G190), .B(new_n538), .C1(new_n541), .C2(new_n364), .ZN(new_n560));
  OAI21_X1  g0360(.A(G200), .B1(new_n556), .B2(new_n537), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n271), .A2(G87), .A3(new_n526), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n551), .A4(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n530), .A2(new_n533), .A3(new_n559), .A4(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n267), .A2(G97), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n527), .B2(new_n463), .ZN(new_n567));
  XNOR2_X1  g0367(.A(G97), .B(G107), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT6), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n569), .A2(new_n463), .A3(G107), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n415), .B2(new_n225), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n567), .B1(new_n575), .B2(new_n265), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n286), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n577), .A2(new_n462), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n224), .A2(G1698), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n425), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n364), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(G257), .B(new_n280), .C1(new_n453), .C2(new_n455), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n478), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n584), .A2(new_n586), .A3(G190), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n585), .A2(new_n478), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT4), .B1(new_n396), .B2(new_n581), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n577), .A2(new_n462), .A3(new_n578), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n290), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(G200), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n576), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n567), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n411), .A2(new_n413), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n412), .B1(new_n285), .B2(G20), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n225), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n571), .B1(new_n569), .B2(new_n568), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n598), .A2(new_n216), .B1(new_n223), .B2(new_n350), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n265), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n588), .A2(new_n591), .A3(new_n389), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n304), .B1(new_n584), .B2(new_n586), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n593), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n564), .A2(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n444), .A2(new_n494), .A3(new_n606), .ZN(G372));
  INV_X1    g0407(.A(new_n306), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n423), .A2(KEYINPUT16), .A3(new_n427), .ZN(new_n609));
  OAI22_X1  g0409(.A1(new_n421), .A2(new_n216), .B1(new_n408), .B2(new_n350), .ZN(new_n610));
  INV_X1    g0410(.A(new_n314), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n376), .A2(new_n378), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(new_n260), .ZN(new_n613));
  INV_X1    g0413(.A(new_n413), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n596), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n610), .B1(new_n615), .B2(G68), .ZN(new_n616));
  INV_X1    g0416(.A(new_n417), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n265), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n402), .B1(new_n609), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n393), .A2(new_n398), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g0421(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n342), .ZN(new_n625));
  INV_X1    g0425(.A(new_n368), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n348), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n442), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n300), .A2(new_n302), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n608), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n444), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n543), .A2(new_n554), .A3(new_n558), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n560), .A2(new_n561), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n551), .A2(new_n562), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT81), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT81), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n551), .A2(new_n562), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n633), .B1(new_n634), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n559), .A2(new_n563), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT26), .B1(new_n644), .B2(new_n604), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n643), .A2(new_n559), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n593), .A2(new_n604), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT82), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n647), .A2(new_n640), .A3(new_n648), .A4(new_n530), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n593), .A2(new_n530), .A3(new_n604), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n551), .A2(new_n562), .A3(new_n637), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n637), .B1(new_n551), .B2(new_n562), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n634), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n559), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT82), .B1(new_n650), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n491), .A2(new_n492), .A3(new_n533), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n649), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n646), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n631), .B1(new_n632), .B2(new_n658), .ZN(G369));
  NAND3_X1  g0459(.A1(new_n266), .A2(new_n216), .A3(G13), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n474), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g0466(.A(new_n666), .B(KEYINPUT84), .Z(new_n667));
  INV_X1    g0467(.A(KEYINPUT85), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n493), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n668), .B2(new_n493), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n488), .A2(new_n489), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n490), .A2(new_n474), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n492), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n665), .B1(new_n523), .B2(new_n528), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n530), .A2(new_n533), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT86), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n530), .A2(KEYINPUT86), .A3(new_n533), .A4(new_n676), .ZN(new_n680));
  INV_X1    g0480(.A(new_n665), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n679), .B(new_n680), .C1(new_n533), .C2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n675), .A2(G330), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n533), .A2(new_n665), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n673), .A2(new_n681), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n683), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n207), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR4_X1   g0492(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n219), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n505), .A2(new_n495), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT87), .B1(new_n697), .B2(new_n542), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n584), .A2(new_n586), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT87), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n557), .A2(new_n700), .A3(new_n505), .A4(new_n495), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n698), .A2(new_n490), .A3(new_n699), .A4(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n480), .A2(new_n389), .A3(new_n542), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n500), .B1(new_n584), .B2(new_n586), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n702), .B2(new_n703), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n681), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT31), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT88), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(KEYINPUT88), .A3(KEYINPUT31), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n494), .A2(new_n606), .A3(new_n681), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n709), .B1(new_n715), .B2(KEYINPUT31), .ZN(new_n716));
  OAI21_X1  g0516(.A(G330), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n644), .A2(new_n604), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n633), .B1(new_n719), .B2(new_n641), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT89), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT26), .B1(new_n654), .B2(new_n604), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n656), .A2(new_n647), .A3(new_n530), .A4(new_n640), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n721), .B1(new_n720), .B2(new_n722), .ZN(new_n726));
  OAI211_X1 g0526(.A(KEYINPUT90), .B(new_n681), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n642), .A2(new_n641), .A3(new_n559), .A4(new_n563), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n559), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT89), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n723), .A3(new_n724), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT90), .B1(new_n733), .B2(new_n681), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT29), .B1(new_n728), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n665), .B1(new_n646), .B2(new_n657), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(KEYINPUT29), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n718), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n696), .B1(new_n739), .B2(G1), .ZN(G364));
  AOI21_X1  g0540(.A(new_n215), .B1(G20), .B2(new_n304), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n216), .A2(new_n294), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n345), .A2(G179), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G303), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n315), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n389), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n216), .A2(G190), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n743), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G322), .A2(new_n749), .B1(new_n752), .B2(G283), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n747), .A2(new_n750), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n755), .A2(G311), .B1(new_n758), .B2(G329), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n216), .B1(new_n756), .B2(G190), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n746), .B(new_n760), .C1(G294), .C2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT93), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n294), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G326), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n765), .A2(G190), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(KEYINPUT33), .B(G317), .Z(new_n770));
  OAI211_X1 g0570(.A(new_n763), .B(new_n767), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT94), .Z(new_n772));
  OAI21_X1  g0572(.A(new_n285), .B1(new_n744), .B2(new_n381), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n751), .A2(new_n225), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n761), .A2(new_n463), .ZN(new_n775));
  OR3_X1    g0575(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(G50), .B2(new_n766), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n247), .B2(new_n769), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G58), .A2(new_n749), .B1(new_n755), .B2(G77), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(KEYINPUT92), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n779), .A2(KEYINPUT92), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n757), .A2(new_n408), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT32), .Z(new_n783));
  NOR4_X1   g0583(.A1(new_n778), .A2(new_n780), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n741), .B1(new_n772), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n216), .A2(G13), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n266), .B1(new_n786), .B2(G45), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n691), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n690), .A2(new_n315), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n791), .A2(G355), .B1(new_n465), .B2(new_n690), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n396), .A2(new_n690), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(G45), .B2(new_n219), .ZN(new_n794));
  INV_X1    g0594(.A(G45), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n251), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n792), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT91), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n741), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n797), .B2(new_n798), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n790), .B1(new_n799), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n802), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n785), .B(new_n806), .C1(new_n675), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G330), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n670), .B2(new_n674), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(new_n789), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n675), .A2(G330), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n808), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT95), .Z(G396));
  NOR2_X1   g0614(.A1(new_n368), .A2(new_n665), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n358), .A2(new_n665), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n371), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n815), .B1(new_n368), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n736), .B(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n789), .B1(new_n819), .B2(new_n717), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n717), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n741), .A2(new_n800), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n789), .B1(new_n823), .B2(G77), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n225), .A2(new_n744), .B1(new_n748), .B2(new_n503), .ZN(new_n825));
  INV_X1    g0625(.A(G311), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n751), .A2(new_n381), .B1(new_n757), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n315), .B1(new_n754), .B2(new_n465), .ZN(new_n828));
  NOR4_X1   g0628(.A1(new_n825), .A2(new_n827), .A3(new_n828), .A4(new_n775), .ZN(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  INV_X1    g0630(.A(new_n766), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n830), .B2(new_n769), .C1(new_n745), .C2(new_n831), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G143), .A2(new_n749), .B1(new_n755), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(G150), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n769), .B2(new_n834), .C1(new_n835), .C2(new_n831), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n752), .A2(G68), .ZN(new_n839));
  INV_X1    g0639(.A(new_n744), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G50), .A2(new_n840), .B1(new_n758), .B2(G132), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n425), .B1(G58), .B2(new_n762), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n838), .A2(new_n839), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n836), .A2(new_n837), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n832), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n824), .B1(new_n845), .B2(new_n741), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n818), .B2(new_n801), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT96), .Z(new_n848));
  AND2_X1   g0648(.A1(new_n821), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n786), .A2(new_n266), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n341), .A2(new_n665), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n342), .A2(new_n348), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n327), .A2(new_n341), .A3(new_n665), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n710), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n855), .B(new_n818), .C1(new_n716), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT98), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n400), .B2(new_n429), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n393), .A2(new_n398), .A3(KEYINPUT77), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT77), .B1(new_n393), .B2(new_n398), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n619), .A3(KEYINPUT98), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT99), .B1(new_n429), .B2(new_n663), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT99), .ZN(new_n867));
  INV_X1    g0667(.A(new_n663), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n619), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n441), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n865), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT100), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT100), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n865), .A2(new_n870), .A3(new_n872), .A4(new_n875), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n441), .A2(KEYINPUT101), .B1(new_n619), .B2(new_n620), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n870), .B(new_n877), .C1(KEYINPUT101), .C2(new_n441), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n874), .A2(new_n876), .B1(KEYINPUT37), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n870), .B1(new_n624), .B2(new_n442), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n858), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT97), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n617), .B1(new_n423), .B2(new_n427), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n883), .B2(new_n333), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n428), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n883), .A2(new_n882), .A3(new_n333), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n402), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n393), .A2(new_n398), .A3(new_n663), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n441), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n441), .A2(new_n871), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n869), .B2(new_n866), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n875), .B1(new_n893), .B2(new_n865), .ZN(new_n894));
  AND4_X1   g0694(.A1(new_n875), .A2(new_n865), .A3(new_n870), .A4(new_n872), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n887), .A2(new_n868), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n431), .B2(new_n442), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(KEYINPUT38), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n857), .B1(new_n881), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n874), .A2(new_n876), .B1(KEYINPUT37), .B2(new_n890), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n903), .A2(new_n858), .A3(new_n898), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n896), .B2(new_n899), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n709), .ZN(new_n907));
  NOR4_X1   g0707(.A1(new_n493), .A2(new_n564), .A3(new_n605), .A4(new_n665), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT31), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n710), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n911), .A2(new_n902), .A3(new_n818), .A4(new_n855), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n901), .A2(new_n902), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT103), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n444), .A2(new_n911), .ZN(new_n915));
  OAI21_X1  g0715(.A(G330), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n916), .A2(KEYINPUT104), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(KEYINPUT104), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n914), .A2(new_n915), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n881), .A2(new_n900), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT102), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT102), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n881), .A2(new_n900), .A3(new_n924), .A4(new_n921), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT39), .B1(new_n904), .B2(new_n905), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n625), .A2(new_n681), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n736), .A2(new_n818), .ZN(new_n931));
  INV_X1    g0731(.A(new_n815), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n855), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n906), .A2(new_n934), .B1(new_n624), .B2(new_n868), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n735), .A2(new_n444), .A3(new_n738), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n631), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n851), .B1(new_n920), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n940), .B2(new_n920), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n943), .A2(G116), .A3(new_n217), .A4(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT36), .Z(new_n946));
  NAND3_X1  g0746(.A1(new_n220), .A2(G77), .A3(new_n406), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n266), .B(G13), .C1(new_n947), .C2(new_n246), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n942), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT105), .Z(G367));
  NAND2_X1  g0751(.A1(new_n766), .A2(G143), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n952), .B1(new_n247), .B2(new_n761), .C1(new_n834), .C2(new_n748), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT113), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n285), .B1(new_n757), .B2(new_n835), .ZN(new_n956));
  INV_X1    g0756(.A(G58), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n744), .A2(new_n957), .B1(new_n754), .B2(new_n202), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n956), .B(new_n958), .C1(G77), .C2(new_n752), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n955), .B(new_n959), .C1(new_n408), .C2(new_n769), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n953), .A2(new_n954), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n744), .A2(new_n465), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(KEYINPUT46), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT112), .Z(new_n964));
  INV_X1    g0764(.A(G317), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n757), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n751), .A2(new_n463), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(G303), .C2(new_n749), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n396), .B1(new_n962), .B2(KEYINPUT46), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n964), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n754), .A2(new_n830), .B1(new_n761), .B2(new_n225), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT111), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n503), .B2(new_n769), .C1(new_n826), .C2(new_n831), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n960), .A2(new_n961), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT114), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n741), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n804), .B1(new_n690), .B2(new_n552), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n241), .A2(new_n793), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n790), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n636), .A2(new_n638), .A3(new_n665), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n640), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n559), .B2(new_n981), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n977), .B(new_n980), .C1(new_n807), .C2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n739), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n686), .B1(new_n679), .B2(new_n680), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n682), .B2(new_n687), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n810), .B(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT29), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n681), .B1(new_n725), .B2(new_n726), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT90), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n990), .B1(new_n993), .B2(new_n727), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n989), .B(new_n717), .C1(new_n994), .C2(new_n737), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n601), .A2(new_n665), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n647), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n642), .A2(new_n665), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n688), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1001), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n688), .A2(new_n999), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT108), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT44), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n688), .A2(new_n999), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n999), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(new_n986), .C2(new_n684), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1008), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1005), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n683), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1005), .A2(new_n1013), .A3(new_n683), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(KEYINPUT109), .B1(new_n995), .B2(new_n1018), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n1005), .A2(new_n1013), .A3(new_n683), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n683), .B1(new_n1005), .B2(new_n1013), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT109), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1022), .A2(new_n739), .A3(new_n1023), .A4(new_n989), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n985), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n691), .B(KEYINPUT41), .Z(new_n1026));
  OAI21_X1  g0826(.A(new_n787), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n986), .A2(new_n999), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n1028), .A2(KEYINPUT106), .A3(KEYINPUT42), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT106), .B1(new_n1028), .B2(KEYINPUT42), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n533), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n647), .A2(new_n1031), .A3(new_n996), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n665), .B1(new_n1032), .B2(new_n604), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n1028), .B2(KEYINPUT42), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1029), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1037), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n683), .A2(new_n1009), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1041), .B(new_n1043), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n1027), .A2(new_n1044), .A3(KEYINPUT110), .ZN(new_n1045));
  AOI21_X1  g0845(.A(KEYINPUT110), .B1(new_n1027), .B2(new_n1044), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n984), .B1(new_n1045), .B2(new_n1046), .ZN(G387));
  OR2_X1    g0847(.A1(new_n682), .A2(new_n807), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n791), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1049), .A2(new_n693), .B1(G107), .B2(new_n207), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n238), .A2(new_n795), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n693), .B(new_n795), .C1(new_n247), .C2(new_n223), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT50), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n349), .B2(G50), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n255), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n793), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1050), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n789), .B1(new_n1059), .B2(new_n804), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G159), .A2(new_n766), .B1(new_n768), .B2(new_n255), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n744), .A2(new_n223), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n761), .A2(new_n352), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n967), .A2(new_n1062), .A3(new_n1063), .A4(new_n425), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n748), .A2(new_n202), .B1(new_n754), .B2(new_n247), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G150), .B2(new_n758), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1061), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n840), .A2(G294), .B1(new_n762), .B2(G283), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n748), .A2(new_n965), .B1(new_n754), .B2(new_n745), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT115), .Z(new_n1070));
  XOR2_X1   g0870(.A(KEYINPUT116), .B(G322), .Z(new_n1071));
  NAND2_X1  g0871(.A1(new_n766), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(new_n826), .C2(new_n769), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT48), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1068), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n1074), .B2(new_n1073), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(KEYINPUT117), .B(KEYINPUT49), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1076), .B(new_n1077), .Z(new_n1078));
  AOI22_X1  g0878(.A1(new_n752), .A2(G116), .B1(new_n758), .B2(G326), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n425), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1067), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1060), .B1(new_n1081), .B2(new_n741), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n989), .A2(new_n788), .B1(new_n1048), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n995), .A2(new_n691), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n739), .A2(new_n989), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(G393));
  AND2_X1   g0886(.A1(new_n995), .A2(new_n1018), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n692), .B(new_n1087), .C1(new_n1024), .C2(new_n1019), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n803), .B1(new_n463), .B2(new_n207), .C1(new_n245), .C2(new_n1057), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n789), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n285), .B(new_n774), .C1(G116), .C2(new_n762), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n768), .A2(G303), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n840), .A2(G283), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G294), .A2(new_n755), .B1(new_n758), .B2(new_n1071), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n766), .A2(G317), .B1(G311), .B2(new_n749), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n766), .A2(G150), .B1(G159), .B2(new_n749), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT51), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n768), .A2(G50), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n255), .A2(new_n755), .B1(new_n752), .B2(G87), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G68), .A2(new_n840), .B1(new_n758), .B2(G143), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n425), .B1(G77), .B2(new_n762), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1095), .A2(new_n1097), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1090), .B1(new_n1105), .B2(new_n741), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n999), .B2(new_n807), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1018), .B2(new_n787), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1088), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(G390));
  OAI21_X1  g0910(.A(new_n789), .B1(new_n823), .B2(new_n255), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n315), .B1(new_n761), .B2(new_n223), .C1(new_n381), .C2(new_n744), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n839), .B1(new_n465), .B2(new_n748), .C1(new_n503), .C2(new_n757), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(G283), .C2(new_n766), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n769), .A2(new_n225), .B1(new_n463), .B2(new_n754), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT121), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1119), .A2(KEYINPUT122), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(KEYINPUT122), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G128), .A2(new_n766), .B1(new_n768), .B2(G137), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1123), .A2(new_n754), .B1(new_n751), .B2(new_n202), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G125), .B2(new_n758), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n744), .A2(new_n834), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  INV_X1    g0927(.A(G132), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n285), .B1(new_n748), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G159), .B2(new_n762), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1122), .A2(new_n1125), .A3(new_n1127), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1120), .A2(new_n1121), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1111), .B1(new_n1132), .B2(new_n741), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n927), .B2(new_n801), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT123), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(KEYINPUT123), .B(new_n1133), .C1(new_n927), .C2(new_n801), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n815), .B1(new_n736), .B2(new_n818), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n855), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n928), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n923), .A2(new_n925), .A3(new_n926), .A4(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n929), .B1(new_n881), .B2(new_n900), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n993), .A2(new_n727), .A3(new_n932), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n817), .A2(new_n368), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1143), .B1(new_n1146), .B2(new_n1140), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n911), .A2(G330), .A3(new_n818), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1149), .A2(new_n1140), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(G330), .B(new_n818), .C1(new_n714), .C2(new_n716), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1152), .A2(new_n1140), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1142), .A2(new_n1147), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1138), .B1(new_n1155), .B2(new_n787), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT120), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1149), .A2(new_n1140), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT119), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1149), .A2(KEYINPUT119), .A3(new_n1140), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1161), .A2(new_n1146), .A3(new_n1153), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT118), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1152), .A2(new_n1164), .A3(new_n1140), .ZN(new_n1165));
  OAI21_X1  g0965(.A(KEYINPUT118), .B1(new_n1149), .B2(new_n1140), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1152), .A2(new_n1140), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n933), .B(new_n1165), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n444), .A2(G330), .A3(new_n911), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n938), .A2(new_n631), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n692), .B1(new_n1155), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1171), .B1(new_n1168), .B2(new_n1163), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1151), .A2(new_n1175), .A3(new_n1154), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1158), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1142), .A2(new_n1147), .A3(new_n1153), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1150), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1173), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  AND4_X1   g0981(.A1(new_n1158), .A2(new_n1181), .A3(new_n691), .A4(new_n1176), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1157), .B1(new_n1177), .B2(new_n1182), .ZN(G378));
  NAND2_X1  g0983(.A1(new_n274), .A2(new_n868), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n307), .B(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1185), .B(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n901), .A2(new_n902), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n858), .B1(new_n903), .B2(new_n898), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n912), .B1(new_n900), .B2(new_n1190), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1188), .B(G330), .C1(new_n1189), .C2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1188), .B1(new_n913), .B2(G330), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n937), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1188), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n857), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n894), .B2(new_n895), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n869), .B(new_n866), .C1(new_n628), .C2(new_n623), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT38), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1197), .B1(new_n904), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1190), .A2(new_n900), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n857), .A2(KEYINPUT40), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1202), .A2(KEYINPUT40), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1196), .B1(new_n1205), .B2(new_n809), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n935), .B1(new_n927), .B2(new_n929), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1207), .A3(new_n1192), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1195), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1196), .A2(new_n800), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n396), .A2(G41), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G50), .B(new_n1211), .C1(new_n260), .C2(new_n450), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n744), .A2(new_n223), .B1(new_n754), .B2(new_n352), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n751), .A2(new_n957), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G283), .B2(new_n758), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n225), .B2(new_n748), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1213), .B(new_n1216), .C1(G68), .C2(new_n762), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G97), .A2(new_n768), .B1(new_n766), .B2(G116), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1211), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT58), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1212), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1220), .B2(new_n1219), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n744), .A2(new_n1123), .ZN(new_n1223));
  INV_X1    g1023(.A(G128), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n748), .A2(new_n1224), .B1(new_n754), .B2(new_n835), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G150), .C2(new_n762), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n766), .A2(G125), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n1128), .C2(new_n769), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n752), .A2(G159), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G33), .B(G41), .C1(new_n758), .C2(G124), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n741), .B1(new_n1222), .B2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT124), .Z(new_n1236));
  AOI211_X1 g1036(.A(new_n790), .B(new_n1236), .C1(new_n202), .C2(new_n822), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1209), .A2(new_n788), .B1(new_n1210), .B2(new_n1237), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1206), .A2(new_n1207), .A3(new_n1192), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1207), .B1(new_n1192), .B2(new_n1206), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1171), .B1(new_n1242), .B2(new_n1169), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n691), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1176), .A2(new_n1172), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT57), .B1(new_n1245), .B2(new_n1209), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1238), .B1(new_n1244), .B2(new_n1246), .ZN(G375));
  INV_X1    g1047(.A(new_n1169), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1171), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1026), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n1173), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n748), .A2(new_n830), .B1(new_n754), .B2(new_n225), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n744), .A2(new_n463), .B1(new_n757), .B2(new_n745), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n315), .B1(new_n751), .B2(new_n223), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .A4(new_n1063), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n465), .B2(new_n769), .C1(new_n503), .C2(new_n831), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n425), .B(new_n1214), .C1(G150), .C2(new_n755), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n748), .A2(new_n835), .B1(new_n757), .B2(new_n1224), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G159), .B2(new_n840), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1257), .B(new_n1259), .C1(new_n202), .C2(new_n761), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1128), .A2(new_n831), .B1(new_n769), .B2(new_n1123), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1256), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1262), .A2(KEYINPUT125), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(KEYINPUT125), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n741), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n790), .B1(new_n822), .B2(new_n247), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1265), .B(new_n1266), .C1(new_n855), .C2(new_n801), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1248), .B2(new_n787), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1251), .A2(new_n1269), .ZN(G381));
  NAND2_X1  g1070(.A1(new_n1210), .A2(new_n1237), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1272), .B2(new_n787), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1245), .A2(new_n1209), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT57), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1195), .B2(new_n1208), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n692), .B1(new_n1277), .B2(new_n1245), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1273), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1156), .B1(new_n1176), .B2(new_n1174), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  OR2_X1    g1081(.A1(G393), .A2(G396), .ZN(new_n1282));
  OR3_X1    g1082(.A1(G390), .A2(G384), .A3(new_n1282), .ZN(new_n1283));
  OR4_X1    g1083(.A1(G387), .A2(new_n1281), .A3(G381), .A4(new_n1283), .ZN(G407));
  OAI211_X1 g1084(.A(G407), .B(G213), .C1(G343), .C2(new_n1281), .ZN(G409));
  NAND4_X1  g1085(.A1(new_n1171), .A2(new_n1163), .A3(new_n1168), .A4(KEYINPUT60), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n691), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1173), .A2(KEYINPUT60), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1287), .B1(new_n1288), .B2(new_n1249), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n849), .B1(new_n1289), .B2(new_n1268), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(KEYINPUT60), .B2(new_n1173), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G384), .B(new_n1269), .C1(new_n1292), .C2(new_n1287), .ZN(new_n1293));
  INV_X1    g1093(.A(G213), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1294), .A2(G343), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(G2897), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1290), .A2(new_n1293), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1296), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1238), .B1(new_n1026), .B2(new_n1274), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n1279), .A2(G378), .B1(new_n1280), .B2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1302), .B2(new_n1295), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1245), .A2(new_n1209), .A3(new_n1250), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1280), .B1(new_n1304), .B2(new_n1273), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1181), .A2(new_n691), .A3(new_n1176), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(KEYINPUT120), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1174), .A2(new_n1158), .A3(new_n1176), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1156), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1305), .B1(G375), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1295), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .A4(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1303), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1279), .A2(G378), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1295), .B1(new_n1318), .B2(new_n1305), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1311), .B1(new_n1319), .B2(new_n1314), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(G387), .A2(new_n1109), .ZN(new_n1322));
  XOR2_X1   g1122(.A(G393), .B(G396), .Z(new_n1323));
  OAI211_X1 g1123(.A(G390), .B(new_n984), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1322), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1323), .B1(new_n1322), .B2(new_n1324), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1299), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1297), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1329), .B1(new_n1312), .B2(new_n1310), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1327), .B(new_n1316), .C1(new_n1330), .C2(KEYINPUT126), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1310), .A2(new_n1312), .A3(new_n1314), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1300), .B(KEYINPUT126), .C1(new_n1302), .C2(new_n1295), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1310), .A2(KEYINPUT63), .A3(new_n1312), .A4(new_n1314), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1334), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  OAI22_X1  g1137(.A1(new_n1321), .A2(new_n1327), .B1(new_n1331), .B2(new_n1337), .ZN(G405));
  NAND2_X1  g1138(.A1(new_n1314), .A2(KEYINPUT127), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(G375), .A2(new_n1280), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(new_n1318), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT127), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1313), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1313), .A2(new_n1342), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1339), .A2(new_n1340), .A3(new_n1318), .A4(new_n1344), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1343), .A2(new_n1327), .A3(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1327), .B1(new_n1343), .B2(new_n1345), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(G402));
endmodule


