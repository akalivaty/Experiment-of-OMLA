//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  INV_X1    g040(.A(G113), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  OAI22_X1  g042(.A1(new_n464), .A2(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G2105), .B1(G101), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n472), .B1(new_n462), .B2(new_n463), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(KEYINPUT65), .A3(new_n472), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n464), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n464), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n483), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n462), .B2(new_n463), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT66), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n476), .A2(new_n494), .A3(new_n491), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n492), .A2(KEYINPUT66), .A3(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n496), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT67), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT67), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(G543), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n508), .A2(new_n511), .B1(KEYINPUT5), .B2(new_n507), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n512), .A2(new_n516), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(G166));
  INV_X1    g097(.A(new_n520), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT68), .B(KEYINPUT7), .ZN(new_n525));
  AND3_X1   g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n517), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT69), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n527), .A2(new_n528), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(G89), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n529), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n514), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(G543), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n520), .A2(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n538), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  AOI22_X1  g119(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n514), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT70), .B(G81), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n520), .A2(new_n547), .B1(new_n548), .B2(new_n541), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT71), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI211_X1 g133(.A(KEYINPUT72), .B(new_n557), .C1(new_n541), .C2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n512), .A2(G91), .A3(new_n516), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n558), .B1(new_n561), .B2(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n557), .A2(KEYINPUT72), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n516), .A2(new_n562), .A3(G543), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n512), .A2(G65), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n514), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n565), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  OAI221_X1 g145(.A(new_n518), .B1(new_n520), .B2(new_n519), .C1(new_n513), .C2(new_n514), .ZN(G303));
  NAND2_X1  g146(.A1(new_n508), .A2(new_n511), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n572), .A2(G87), .A3(new_n573), .A4(new_n516), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n572), .A2(new_n573), .ZN(new_n580));
  INV_X1    g155(.A(G74), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n514), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n574), .A2(new_n575), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT73), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G288));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  INV_X1    g162(.A(G48), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n520), .A2(new_n587), .B1(new_n588), .B2(new_n541), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n512), .A2(G61), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n514), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT74), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n596));
  NOR3_X1   g171(.A1(new_n596), .A2(KEYINPUT74), .A3(new_n514), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n595), .B2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n517), .A2(G47), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n512), .A2(G85), .A3(new_n516), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT75), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT75), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n599), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G72), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n580), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n602), .A2(new_n604), .B1(G651), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G301), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n520), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n512), .A2(KEYINPUT10), .A3(G92), .A4(new_n516), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n580), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n619), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT76), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n616), .A2(new_n620), .A3(KEYINPUT76), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n611), .B1(new_n625), .B2(new_n610), .ZN(G284));
  AOI21_X1  g201(.A(new_n611), .B1(new_n625), .B2(new_n610), .ZN(G321));
  NOR2_X1   g202(.A1(G299), .A2(G868), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g204(.A(new_n628), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n625), .B1(new_n631), .B2(G860), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT77), .ZN(G148));
  AND3_X1   g208(.A1(new_n616), .A2(new_n620), .A3(KEYINPUT76), .ZN(new_n634));
  AOI21_X1  g209(.A(KEYINPUT76), .B1(new_n616), .B2(new_n620), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n631), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n637), .B(KEYINPUT78), .C1(G868), .C2(new_n550), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(KEYINPUT78), .B2(new_n637), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n476), .A2(new_n469), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT80), .B(G2100), .Z(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI22_X1  g221(.A1(G123), .A2(new_n484), .B1(new_n481), .B2(G135), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n483), .A2(KEYINPUT81), .A3(G111), .ZN(new_n648));
  OAI21_X1  g223(.A(KEYINPUT81), .B1(new_n483), .B2(G111), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n649), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n647), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n644), .A2(new_n645), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n646), .A2(new_n652), .A3(new_n653), .ZN(G156));
  XOR2_X1   g229(.A(KEYINPUT15), .B(G2435), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2438), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2443), .B(G2446), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT83), .ZN(new_n665));
  XOR2_X1   g240(.A(G2451), .B(G2454), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1341), .B(G1348), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT85), .ZN(new_n671));
  OAI21_X1  g246(.A(G14), .B1(new_n668), .B2(new_n669), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2067), .B(G2678), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT86), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT18), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n676), .B(KEYINPUT17), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n681), .B(new_n678), .C1(new_n675), .C2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n675), .A3(new_n677), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G2100), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT87), .B(G2096), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G227));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1961), .B(G1966), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT20), .Z(new_n696));
  AND2_X1   g271(.A1(new_n692), .A2(new_n693), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT88), .ZN(new_n699));
  NOR3_X1   g274(.A1(new_n691), .A2(new_n694), .A3(new_n697), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1991), .B(G1996), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT89), .B(KEYINPUT90), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1981), .B(G1986), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n703), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(G229));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n711), .A2(G6), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G305), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT32), .B(G1981), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n711), .ZN(new_n718));
  INV_X1    g293(.A(G1971), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n713), .A2(new_n715), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n711), .A2(G23), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n582), .A2(new_n583), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n711), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT33), .B(G1976), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  AND4_X1   g301(.A1(new_n716), .A2(new_n720), .A3(new_n721), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n481), .A2(G131), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n484), .A2(G119), .ZN(new_n734));
  OR2_X1    g309(.A1(G95), .A2(G2105), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n735), .B(G2104), .C1(G107), .C2(new_n483), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n732), .B1(new_n738), .B2(new_n731), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n608), .A2(new_n711), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n711), .B2(G24), .ZN(new_n743));
  INV_X1    g318(.A(G1986), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n744), .B2(new_n743), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n729), .A2(new_n730), .A3(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT36), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n711), .A2(G21), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G168), .B2(new_n711), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(G1966), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(G1966), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n731), .A2(G26), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n481), .A2(G140), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n484), .A2(G128), .ZN(new_n756));
  OR2_X1    g331(.A1(G104), .A2(G2105), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n757), .B(G2104), .C1(G116), .C2(new_n483), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n754), .B1(new_n760), .B2(new_n731), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT91), .B(G2067), .Z(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT30), .B(G28), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n765), .A2(new_n731), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n651), .B2(new_n731), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n763), .A2(new_n764), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n731), .A2(G27), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G164), .B2(new_n731), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(new_n443), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n751), .A2(new_n752), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G1348), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n625), .A2(new_n711), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G4), .B2(new_n711), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n774), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n711), .A2(G20), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT23), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n565), .A2(new_n568), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n711), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT98), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT97), .B(G1956), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n778), .B(new_n785), .C1(new_n775), .C2(new_n777), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n481), .A2(G141), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT95), .Z(new_n788));
  AND2_X1   g363(.A1(new_n469), .A2(G105), .ZN(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT26), .ZN(new_n791));
  AOI211_X1 g366(.A(new_n789), .B(new_n791), .C1(G129), .C2(new_n484), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G32), .B(new_n793), .S(G29), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT27), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1996), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n797));
  INV_X1    g372(.A(G34), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n731), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n798), .B2(new_n797), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n479), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2084), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n731), .A2(G35), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G162), .B2(new_n731), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT29), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n802), .B1(new_n806), .B2(G2090), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n711), .A2(G5), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G171), .B2(new_n711), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1961), .ZN(new_n810));
  NOR2_X1   g385(.A1(G29), .A2(G33), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT92), .Z(new_n812));
  AOI22_X1  g387(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(new_n483), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n818));
  NAND2_X1  g393(.A1(G103), .A2(G2104), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(G2105), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n483), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n481), .A2(G139), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n816), .A2(new_n817), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n812), .B1(new_n823), .B2(new_n731), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n442), .ZN(new_n825));
  NOR2_X1   g400(.A1(G16), .A2(G19), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n550), .B2(G16), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1341), .ZN(new_n828));
  NOR4_X1   g403(.A1(new_n807), .A2(new_n810), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n806), .A2(G2090), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT96), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n796), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n748), .A2(new_n786), .A3(new_n832), .ZN(G311));
  INV_X1    g408(.A(G311), .ZN(G150));
  NAND2_X1  g409(.A1(new_n625), .A2(G559), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT38), .Z(new_n836));
  AOI22_X1  g411(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n837), .A2(new_n514), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT99), .B(G93), .Z(new_n839));
  INV_X1    g414(.A(G55), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n520), .A2(new_n839), .B1(new_n840), .B2(new_n541), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n550), .A2(new_n842), .ZN(new_n843));
  OAI22_X1  g418(.A1(new_n546), .A2(new_n549), .B1(new_n838), .B2(new_n841), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n836), .B(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  INV_X1    g422(.A(G860), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n842), .A2(new_n848), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(G145));
  XNOR2_X1  g428(.A(new_n651), .B(new_n488), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n479), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n481), .A2(G142), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT100), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n484), .A2(G130), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n483), .A2(G118), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n737), .B(new_n643), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n760), .B(new_n505), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n823), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(new_n793), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n793), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n865), .A2(new_n866), .B1(new_n870), .B2(new_n871), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n855), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n867), .A2(new_n872), .ZN(new_n876));
  INV_X1    g451(.A(new_n855), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n876), .B(new_n877), .C1(new_n872), .C2(new_n863), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n875), .A2(new_n878), .A3(KEYINPUT102), .A4(new_n879), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n882), .A2(KEYINPUT40), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT40), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(G395));
  NAND2_X1  g461(.A1(G305), .A2(new_n608), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(G166), .B1(new_n582), .B2(new_n583), .ZN(new_n889));
  NAND2_X1  g464(.A1(G303), .A2(new_n723), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(G305), .A2(new_n608), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n888), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n597), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT74), .B1(new_n596), .B2(new_n514), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n589), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(G290), .A2(new_n896), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n897), .A2(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT106), .B1(new_n893), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n891), .B1(new_n888), .B2(new_n892), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n897), .A2(new_n887), .A3(new_n889), .A4(new_n890), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(KEYINPUT42), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n900), .A2(new_n901), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(KEYINPUT106), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n843), .A2(new_n844), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n636), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n625), .A2(new_n631), .A3(new_n845), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(G299), .A2(new_n616), .A3(new_n620), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n621), .A2(KEYINPUT103), .A3(new_n781), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT103), .B1(new_n621), .B2(new_n781), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT104), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n914), .A4(new_n915), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n913), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n916), .B2(new_n917), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n919), .A2(KEYINPUT41), .A3(new_n914), .A4(new_n915), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n911), .A2(new_n912), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n923), .A2(new_n929), .A3(KEYINPUT105), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n932), .A3(new_n928), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n931), .B1(new_n930), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n909), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(new_n933), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT107), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n908), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n610), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n842), .A2(G868), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT108), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n943));
  INV_X1    g518(.A(new_n941), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n935), .A2(new_n909), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n947), .B2(new_n909), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n943), .B(new_n944), .C1(new_n948), .C2(new_n610), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n942), .A2(new_n949), .ZN(G295));
  OAI21_X1  g525(.A(KEYINPUT109), .B1(new_n940), .B2(new_n941), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n952), .B(new_n944), .C1(new_n948), .C2(new_n610), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n951), .A2(new_n953), .ZN(G331));
  NAND2_X1  g529(.A1(G168), .A2(G171), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n531), .A2(G301), .A3(new_n535), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n910), .A3(new_n956), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n531), .A2(G301), .A3(new_n535), .ZN(new_n958));
  AOI21_X1  g533(.A(G301), .B1(new_n531), .B2(new_n535), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n845), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n927), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n960), .B(new_n957), .C1(new_n917), .C2(new_n916), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n905), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n879), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n957), .A2(new_n960), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n922), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(KEYINPUT111), .A3(new_n922), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n925), .A2(new_n926), .A3(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n972), .B(new_n961), .C1(new_n971), .C2(new_n926), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n905), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n965), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT112), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n980), .A3(new_n977), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n905), .B1(new_n962), .B2(new_n963), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT43), .B1(new_n965), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n979), .A2(new_n981), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n962), .A2(new_n963), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n975), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(new_n964), .A3(new_n977), .A4(new_n879), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n977), .B2(new_n976), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n988), .A2(new_n989), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT44), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n985), .A2(new_n993), .ZN(G397));
  INV_X1    g569(.A(KEYINPUT124), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n494), .B1(new_n476), .B2(new_n491), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n503), .B1(new_n497), .B2(new_n996), .ZN(new_n997));
  AOI211_X1 g572(.A(KEYINPUT50), .B(G1384), .C1(new_n997), .C2(new_n496), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n505), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g577(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n1003));
  NAND2_X1  g578(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n465), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n466), .A2(new_n467), .ZN(new_n1006));
  OAI21_X1  g581(.A(G2105), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n469), .A2(G101), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n478), .A2(G40), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n470), .A2(KEYINPUT114), .A3(G40), .A4(new_n478), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1956), .B1(new_n1002), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n1016), .B(G1384), .C1(new_n997), .C2(new_n496), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n505), .B2(new_n1000), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT56), .B(G2072), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NOR4_X1   g595(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n995), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n781), .B(KEYINPUT57), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(new_n1013), .A3(new_n1019), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n498), .A2(new_n502), .A3(new_n499), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1000), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n505), .A2(new_n999), .A3(new_n1000), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n1011), .A3(new_n1012), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1956), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1026), .A2(new_n1034), .A3(KEYINPUT124), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1022), .A2(new_n1024), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1032), .A2(KEYINPUT122), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1013), .A2(new_n1039), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n775), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1384), .B1(new_n997), .B2(new_n496), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1011), .A2(new_n1042), .A3(new_n1012), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1011), .A2(new_n1042), .A3(KEYINPUT121), .A4(new_n1012), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G2067), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1041), .A2(new_n1049), .A3(KEYINPUT123), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT123), .B1(new_n1041), .B2(new_n1049), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1026), .A2(new_n1034), .A3(new_n1023), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1054), .A2(new_n625), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1037), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1054), .A2(KEYINPUT61), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1024), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1054), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT61), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1036), .A2(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT58), .B(G1341), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1029), .A2(new_n1016), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(new_n1011), .A3(new_n1012), .A4(new_n1064), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1047), .A2(new_n1062), .B1(G1996), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n550), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT59), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1069), .A3(new_n550), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n625), .A2(KEYINPUT60), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1041), .A2(new_n1049), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1075), .B2(new_n1050), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n625), .A2(KEYINPUT60), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(KEYINPUT125), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1061), .B(new_n1071), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g654(.A(new_n1078), .B1(KEYINPUT60), .B2(new_n625), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1056), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1961), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1038), .A2(new_n1083), .A3(new_n1040), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1065), .B2(G2078), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1009), .A2(new_n1085), .A3(G2078), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1025), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1084), .A2(G301), .A3(new_n1086), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1084), .A2(new_n1086), .A3(new_n1092), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G171), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1098), .B(KEYINPUT54), .C1(G171), .C2(new_n1089), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n531), .A2(new_n535), .A3(G8), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n1101), .B2(KEYINPUT126), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1015), .A2(new_n998), .A3(new_n1001), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT119), .B(G2084), .ZN(new_n1105));
  INV_X1    g680(.A(G1966), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1104), .A2(new_n1105), .B1(new_n1065), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G8), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1103), .B(new_n1101), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1105), .ZN(new_n1110));
  OAI22_X1  g685(.A1(new_n1087), .A2(G1966), .B1(new_n1032), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(G8), .B(new_n1102), .C1(new_n1111), .C2(G286), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1111), .A2(G8), .A3(G286), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1096), .A2(new_n1099), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT55), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1117), .A2(KEYINPUT115), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(KEYINPUT115), .ZN(new_n1119));
  AOI22_X1  g694(.A1(G303), .A2(G8), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(G8), .B(new_n1119), .C1(new_n515), .C2(new_n521), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G2090), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1104), .A2(new_n1124), .B1(new_n1065), .B2(new_n719), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1125), .B2(new_n1108), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n578), .A2(G1976), .A3(new_n574), .A4(new_n575), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT116), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n576), .A2(new_n1129), .A3(G1976), .A4(new_n578), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1043), .A2(G8), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n585), .A2(G1976), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1132), .B(new_n1133), .C1(KEYINPUT52), .C2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1134), .A2(G8), .A3(new_n1043), .A4(new_n1131), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT52), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1043), .A2(new_n1131), .A3(new_n1133), .A4(G8), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(G1981), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1141), .B(new_n590), .C1(new_n595), .C2(new_n597), .ZN(new_n1142));
  OAI21_X1  g717(.A(G1981), .B1(new_n589), .B2(new_n593), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT118), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT49), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1043), .A2(G8), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT49), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(KEYINPUT118), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1002), .A2(new_n1124), .A3(new_n1013), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1065), .A2(new_n719), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1123), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(G8), .A3(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1126), .A2(new_n1140), .A3(new_n1150), .A4(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1108), .B(new_n1123), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1154), .B1(new_n1153), .B2(G8), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1148), .B1(new_n1144), .B2(KEYINPUT118), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1163), .B(KEYINPUT49), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1165), .A2(new_n1147), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1161), .A2(KEYINPUT127), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1158), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1116), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1082), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1107), .A2(new_n1108), .A3(G286), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1171), .B1(new_n1156), .B2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1161), .A2(KEYINPUT63), .A3(new_n1166), .A4(new_n1172), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OR2_X1    g751(.A1(G288), .A2(G1976), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1142), .B1(new_n1165), .B2(new_n1177), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1166), .A2(new_n1159), .B1(new_n1178), .B2(new_n1147), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1176), .A2(KEYINPUT120), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1090), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1115), .A2(KEYINPUT62), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1186), .A2(new_n1187), .A3(new_n1158), .A4(new_n1167), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1170), .A2(new_n1180), .A3(new_n1183), .A4(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1015), .A2(new_n1063), .ZN(new_n1190));
  INV_X1    g765(.A(G1996), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n793), .B(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n759), .B(new_n1048), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n738), .A2(new_n740), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n738), .A2(new_n740), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n608), .A2(new_n744), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n608), .A2(new_n744), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1190), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1189), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1193), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1190), .B1(new_n1203), .B2(new_n793), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1205));
  AND2_X1   g780(.A1(new_n1205), .A2(KEYINPUT46), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1205), .A2(KEYINPUT46), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1204), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT47), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n1198), .A2(new_n1063), .A3(new_n1015), .ZN(new_n1210));
  AOI22_X1  g785(.A1(new_n1196), .A2(new_n1190), .B1(KEYINPUT48), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1211), .B1(KEYINPUT48), .B2(new_n1210), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1213));
  OAI22_X1  g788(.A1(new_n1213), .A2(new_n1194), .B1(G2067), .B2(new_n759), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1214), .A2(new_n1190), .ZN(new_n1215));
  AND3_X1   g790(.A1(new_n1209), .A2(new_n1212), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1202), .A2(new_n1216), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g792(.A1(new_n979), .A2(new_n981), .A3(new_n984), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n882), .A2(new_n883), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n688), .A2(new_n709), .A3(G319), .ZN(new_n1221));
  NOR2_X1   g795(.A1(G401), .A2(new_n1221), .ZN(new_n1222));
  AND3_X1   g796(.A1(new_n1219), .A2(new_n1220), .A3(new_n1222), .ZN(G308));
  NAND3_X1  g797(.A1(new_n1219), .A2(new_n1220), .A3(new_n1222), .ZN(G225));
endmodule


