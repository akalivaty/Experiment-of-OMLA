//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G43gat), .ZN(new_n204));
  INV_X1    g003(.A(G43gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G50gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT85), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT85), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT14), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n208), .A2(new_n211), .A3(new_n218), .A4(KEYINPUT15), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT15), .B1(new_n209), .B2(new_n210), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT85), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n208), .A2(new_n211), .A3(KEYINPUT86), .A4(KEYINPUT15), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n214), .A2(new_n216), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT89), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT89), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n217), .A3(new_n230), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n203), .A2(KEYINPUT87), .A3(G43gat), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT87), .B1(new_n203), .B2(G43gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n205), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT15), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n231), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n220), .B1(new_n226), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G8gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(G15gat), .B(G22gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT16), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(G1gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT90), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n242), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(G1gat), .B2(new_n243), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI221_X1 g048(.A(new_n245), .B1(new_n246), .B2(new_n242), .C1(G1gat), .C2(new_n243), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n202), .B1(new_n241), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n250), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT15), .ZN(new_n254));
  OR2_X1    g053(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n255));
  AOI21_X1  g054(.A(G43gat), .B1(new_n255), .B2(new_n235), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT87), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n205), .B2(G50gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n203), .A2(KEYINPUT87), .A3(G43gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n254), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n261), .A2(new_n217), .A3(new_n229), .A4(new_n230), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n262), .B1(new_n224), .B2(new_n225), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n253), .B1(new_n263), .B2(new_n220), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n252), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G229gat), .A2(G233gat), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n266), .B(KEYINPUT13), .Z(new_n267));
  INV_X1    g066(.A(new_n241), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(new_n202), .A3(new_n253), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n265), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT92), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT17), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n241), .A2(KEYINPUT17), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n251), .A3(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n275), .A2(KEYINPUT18), .A3(new_n266), .A4(new_n264), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n251), .B1(new_n241), .B2(KEYINPUT17), .ZN(new_n277));
  AOI211_X1 g076(.A(new_n272), .B(new_n220), .C1(new_n226), .C2(new_n240), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n266), .B(new_n264), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT18), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT92), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n265), .A2(new_n282), .A3(new_n269), .A4(new_n267), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n271), .A2(new_n276), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G113gat), .B(G141gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G169gat), .B(G197gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT12), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n271), .A2(new_n276), .A3(new_n283), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n279), .A2(KEYINPUT93), .A3(new_n280), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n290), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT93), .B1(new_n279), .B2(new_n280), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT22), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT68), .B(G211gat), .ZN(new_n300));
  INV_X1    g099(.A(G218gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G211gat), .B(G218gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT3), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(G141gat), .B(G148gat), .Z(new_n312));
  INV_X1    g111(.A(G155gat), .ZN(new_n313));
  INV_X1    g112(.A(G162gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(KEYINPUT2), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n312), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G141gat), .B(G148gat), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n316), .B(new_n315), .C1(new_n320), .C2(KEYINPUT2), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n325), .A2(new_n310), .ZN(new_n326));
  OAI22_X1  g125(.A1(new_n311), .A2(new_n323), .B1(new_n326), .B2(new_n309), .ZN(new_n327));
  INV_X1    g126(.A(new_n308), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n305), .B1(new_n302), .B2(new_n303), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n310), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT75), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G228gat), .A2(G233gat), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n332), .A2(G22gat), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G22gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n326), .B2(new_n309), .ZN(new_n337));
  INV_X1    g136(.A(new_n333), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n327), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n324), .B1(new_n330), .B2(KEYINPUT29), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n341), .A2(new_n322), .B1(new_n331), .B2(new_n330), .ZN(new_n342));
  OAI21_X1  g141(.A(G22gat), .B1(new_n332), .B2(new_n333), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n337), .A2(new_n335), .A3(new_n338), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G78gat), .B(G106gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT31), .B(G50gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT76), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n346), .A2(new_n352), .A3(new_n349), .ZN(new_n353));
  INV_X1    g152(.A(new_n349), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n340), .A2(new_n354), .A3(new_n345), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n340), .A2(KEYINPUT77), .A3(new_n345), .A4(new_n354), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n351), .A2(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT5), .ZN(new_n360));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(G127gat), .B(G134gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G113gat), .B(G120gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n363), .B1(KEYINPUT1), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(KEYINPUT65), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367));
  INV_X1    g166(.A(G120gat), .ZN(new_n368));
  OR3_X1    g167(.A1(new_n368), .A2(KEYINPUT65), .A3(G113gat), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n366), .A2(new_n367), .A3(new_n362), .A4(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n323), .A2(new_n365), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n365), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n322), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n361), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n360), .B1(new_n374), .B2(KEYINPUT74), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(KEYINPUT74), .B2(new_n374), .ZN(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT0), .ZN(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n372), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n323), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(new_n372), .A3(new_n325), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(new_n372), .B2(new_n322), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n361), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n360), .A2(KEYINPUT73), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n376), .B(new_n381), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT81), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n388), .A2(new_n389), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT79), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n371), .A2(new_n361), .A3(new_n373), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT39), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT39), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n407), .A3(new_n380), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(KEYINPUT40), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(KEYINPUT40), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n405), .A2(new_n407), .A3(new_n380), .A4(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n400), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G183gat), .A2(G190gat), .ZN(new_n414));
  INV_X1    g213(.A(G169gat), .ZN(new_n415));
  INV_X1    g214(.A(G176gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT26), .ZN(new_n418));
  NOR2_X1   g217(.A1(G169gat), .A2(G176gat), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT26), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n418), .B(new_n421), .C1(new_n415), .C2(new_n416), .ZN(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT27), .B(G183gat), .ZN(new_n423));
  INV_X1    g222(.A(G190gat), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n423), .A2(KEYINPUT28), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT28), .B1(new_n423), .B2(new_n424), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n414), .B(new_n422), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n419), .A2(KEYINPUT23), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT64), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n419), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT23), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n430), .A2(new_n431), .B1(new_n432), .B2(new_n417), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n414), .ZN(new_n435));
  NAND3_X1  g234(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n435), .A2(new_n436), .B1(G169gat), .B2(G176gat), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT25), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n417), .A2(new_n432), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n439), .A2(KEYINPUT25), .A3(new_n428), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n440), .A2(new_n437), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n427), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n310), .ZN(new_n443));
  NAND2_X1  g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n444), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n448), .A2(new_n330), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT69), .ZN(new_n450));
  INV_X1    g249(.A(new_n447), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n446), .B1(new_n442), .B2(new_n310), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n445), .A2(KEYINPUT69), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n309), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT70), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n449), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT69), .B1(new_n445), .B2(new_n447), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n452), .A2(new_n450), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n330), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT70), .ZN(new_n461));
  XNOR2_X1  g260(.A(G8gat), .B(G36gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT71), .ZN(new_n463));
  XNOR2_X1  g262(.A(G64gat), .B(G92gat), .ZN(new_n464));
  XOR2_X1   g263(.A(new_n463), .B(new_n464), .Z(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n457), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n456), .B(new_n330), .C1(new_n458), .C2(new_n459), .ZN(new_n470));
  INV_X1    g269(.A(new_n449), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n455), .A2(new_n456), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n457), .A2(new_n461), .A3(KEYINPUT30), .A4(new_n466), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n469), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n359), .B1(new_n413), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n472), .A2(new_n473), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT37), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n465), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n478), .A2(new_n479), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT38), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n376), .B1(new_n393), .B2(new_n394), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n380), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n397), .A2(new_n484), .A3(new_n486), .A4(new_n399), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n396), .A2(KEYINPUT6), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n487), .A2(new_n488), .A3(new_n467), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT38), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n453), .A2(new_n309), .A3(new_n454), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT82), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n448), .A2(new_n330), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n491), .A2(KEYINPUT82), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT37), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n480), .A2(new_n490), .A3(new_n465), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n483), .A2(new_n489), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n477), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(G227gat), .A2(G233gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n442), .A2(new_n382), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n372), .B(new_n427), .C1(new_n438), .C2(new_n441), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n503), .A2(new_n504), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n501), .A2(new_n500), .A3(new_n502), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT32), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G43gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(G71gat), .B(G99gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n509), .B1(new_n513), .B2(KEYINPUT33), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT66), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n509), .A2(KEYINPUT33), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n516), .B1(new_n518), .B2(new_n513), .ZN(new_n519));
  AOI211_X1 g318(.A(KEYINPUT66), .B(new_n512), .C1(new_n508), .C2(new_n517), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n507), .B(new_n515), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT67), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n524));
  INV_X1    g323(.A(new_n507), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n521), .A2(new_n522), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n528), .A2(KEYINPUT36), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n526), .A2(new_n521), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT36), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n357), .A2(new_n358), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n352), .B1(new_n346), .B2(new_n349), .ZN(new_n534));
  AOI211_X1 g333(.A(KEYINPUT76), .B(new_n354), .C1(new_n340), .C2(new_n345), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT78), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n474), .A2(new_n475), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT72), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT72), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n474), .A2(new_n475), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n486), .A2(new_n484), .A3(new_n395), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n542), .A2(new_n488), .B1(new_n467), .B2(new_n468), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n499), .A2(new_n532), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT83), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n526), .A2(new_n521), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n359), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n536), .A3(KEYINPUT83), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT35), .B1(new_n551), .B2(new_n544), .ZN(new_n552));
  INV_X1    g351(.A(new_n476), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n487), .A2(new_n488), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n359), .A2(KEYINPUT35), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n528), .A2(new_n553), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n298), .B1(new_n546), .B2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G190gat), .B(G218gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT96), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(KEYINPUT97), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(KEYINPUT8), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n565), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G99gat), .B(G106gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n568), .A2(new_n569), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(new_n571), .A3(new_n565), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n273), .A2(new_n274), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  AND2_X1   g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n268), .A2(new_n578), .B1(KEYINPUT41), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n561), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n560), .A2(KEYINPUT97), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  OR2_X1    g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G57gat), .B(G64gat), .Z(new_n590));
  INV_X1    g389(.A(G71gat), .ZN(new_n591));
  INV_X1    g390(.A(G78gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT9), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n590), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G57gat), .B(G64gat), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n594), .B(new_n593), .C1(new_n599), .C2(new_n596), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  OAI21_X1  g404(.A(new_n251), .B1(new_n602), .B2(new_n601), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT95), .ZN(new_n609));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT94), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n609), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n607), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n589), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n570), .A2(new_n572), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n571), .B1(new_n574), .B2(new_n565), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n601), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n573), .A2(new_n575), .A3(new_n600), .A4(new_n598), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(KEYINPUT98), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n576), .A2(new_n623), .A3(new_n601), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT10), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n617), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n617), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n622), .A2(new_n629), .A3(new_n624), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G120gat), .B(G148gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT99), .ZN(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  OR2_X1    g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n616), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n558), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n542), .A2(new_n488), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g442(.A1(new_n640), .A2(new_n553), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT16), .B(G8gat), .Z(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(KEYINPUT42), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n644), .B(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n648), .A2(new_n645), .ZN(new_n649));
  OAI221_X1 g448(.A(new_n646), .B1(new_n648), .B2(new_n242), .C1(new_n649), .C2(KEYINPUT42), .ZN(G1325gat));
  OAI21_X1  g449(.A(G15gat), .B1(new_n640), .B2(new_n532), .ZN(new_n651));
  INV_X1    g450(.A(new_n528), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n652), .A2(G15gat), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n651), .B1(new_n640), .B2(new_n653), .ZN(G1326gat));
  INV_X1    g453(.A(new_n537), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT101), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT43), .B(G22gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  NOR3_X1   g458(.A1(new_n589), .A2(new_n615), .A3(new_n638), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n558), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n641), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n212), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT45), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n546), .A2(new_n557), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT44), .B1(new_n666), .B2(new_n589), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n552), .A2(KEYINPUT103), .A3(new_n556), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT103), .B1(new_n552), .B2(new_n556), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n546), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n587), .A2(new_n588), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n615), .ZN(new_n675));
  INV_X1    g474(.A(new_n638), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n292), .B2(new_n297), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n284), .A2(new_n291), .ZN(new_n679));
  INV_X1    g478(.A(new_n296), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n290), .A3(new_n294), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n679), .B(KEYINPUT102), .C1(new_n293), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n674), .A2(new_n675), .A3(new_n676), .A4(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(G29gat), .B1(new_n685), .B2(new_n641), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n665), .A2(new_n686), .ZN(G1328gat));
  NOR2_X1   g486(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n553), .A2(G36gat), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n662), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G36gat), .B1(new_n685), .B2(new_n553), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(G1329gat));
  OAI21_X1  g493(.A(new_n205), .B1(new_n661), .B2(new_n652), .ZN(new_n695));
  INV_X1    g494(.A(new_n532), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G43gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n685), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g498(.A1(new_n236), .A2(new_n237), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n685), .B2(new_n536), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n662), .A2(KEYINPUT106), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n537), .B(new_n700), .C1(new_n661), .C2(new_n704), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n702), .B(KEYINPUT48), .C1(new_n703), .C2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n703), .A2(new_n705), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n685), .A2(new_n655), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n708), .B2(new_n701), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n706), .B1(new_n709), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g509(.A1(new_n684), .A2(new_n616), .A3(new_n676), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n670), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n663), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g514(.A1(new_n712), .A2(new_n553), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  AND2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n716), .B2(new_n717), .ZN(G1333gat));
  NAND3_X1  g519(.A1(new_n713), .A2(G71gat), .A3(new_n696), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n591), .B1(new_n712), .B2(new_n652), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n721), .A2(KEYINPUT108), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1334gat));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n655), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(new_n592), .ZN(G1335gat));
  NOR2_X1   g530(.A1(new_n684), .A2(new_n615), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n638), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n667), .B2(new_n673), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735), .B2(new_n641), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n670), .A2(new_n671), .A3(new_n732), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n676), .B1(new_n739), .B2(KEYINPUT109), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(KEYINPUT109), .B2(new_n739), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n663), .A2(new_n563), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n736), .B1(new_n741), .B2(new_n742), .ZN(G1336gat));
  AOI21_X1  g542(.A(new_n564), .B1(new_n734), .B2(new_n476), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n737), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n738), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n737), .A2(new_n747), .A3(KEYINPUT51), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n553), .A2(G92gat), .A3(new_n676), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n744), .B2(new_n745), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT52), .B1(new_n746), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT52), .B1(new_n739), .B2(new_n751), .ZN(new_n755));
  INV_X1    g554(.A(new_n744), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(G1337gat));
  OAI21_X1  g557(.A(G99gat), .B1(new_n735), .B2(new_n532), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n652), .A2(G99gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n741), .B2(new_n760), .ZN(G1338gat));
  NOR3_X1   g560(.A1(new_n536), .A2(G106gat), .A3(new_n676), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n749), .A2(new_n750), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(G106gat), .B1(new_n735), .B2(new_n655), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n749), .A2(KEYINPUT112), .A3(new_n750), .A4(new_n762), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT53), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT53), .B1(new_n739), .B2(new_n762), .ZN(new_n770));
  OAI21_X1  g569(.A(G106gat), .B1(new_n735), .B2(new_n536), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(G1339gat));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n774), .B(new_n617), .C1(new_n625), .C2(new_n627), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n775), .A2(new_n635), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n622), .A2(new_n624), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n626), .ZN(new_n778));
  INV_X1    g577(.A(new_n627), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n629), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n628), .A3(KEYINPUT54), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n776), .A2(KEYINPUT55), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n776), .A2(new_n781), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n776), .A2(KEYINPUT113), .A3(new_n781), .A4(KEYINPUT55), .ZN(new_n788));
  AND4_X1   g587(.A1(new_n636), .A2(new_n784), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n678), .A2(new_n682), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n297), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n266), .B1(new_n275), .B2(new_n264), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n267), .B1(new_n265), .B2(new_n269), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n289), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n638), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n671), .B1(new_n790), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n791), .A2(new_n794), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n788), .A2(new_n636), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n787), .A3(new_n784), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n589), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n675), .B1(new_n796), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n639), .A2(new_n683), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n537), .A2(new_n652), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n476), .A2(new_n641), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(G113gat), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n807), .A2(new_n808), .A3(new_n298), .ZN(new_n809));
  INV_X1    g608(.A(new_n551), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n803), .A2(new_n663), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n641), .B1(new_n801), .B2(new_n802), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(KEYINPUT114), .A3(new_n810), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n476), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n684), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n809), .B1(new_n817), .B2(new_n808), .ZN(G1340gat));
  NOR3_X1   g617(.A1(new_n807), .A2(new_n368), .A3(new_n676), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n638), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n368), .ZN(G1341gat));
  AND3_X1   g620(.A1(new_n806), .A2(G127gat), .A3(new_n615), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n816), .A2(new_n615), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(G127gat), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(G1342gat));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n589), .A2(G134gat), .ZN(new_n829));
  AND4_X1   g628(.A1(KEYINPUT114), .A2(new_n803), .A3(new_n663), .A4(new_n810), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT114), .B1(new_n814), .B2(new_n810), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n553), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT116), .B1(new_n832), .B2(KEYINPUT56), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n816), .A2(new_n834), .A3(new_n835), .A4(new_n829), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(G134gat), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n806), .B2(new_n671), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n832), .A2(new_n842), .A3(KEYINPUT56), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n832), .B2(KEYINPUT56), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n828), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n839), .B1(new_n833), .B2(new_n836), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n847), .B(KEYINPUT118), .C1(new_n844), .C2(new_n843), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1343gat));
  AND2_X1   g648(.A1(new_n532), .A2(new_n805), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n536), .B1(new_n801), .B2(new_n802), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(KEYINPUT57), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n537), .A2(KEYINPUT57), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT55), .B1(new_n785), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n776), .A2(KEYINPUT119), .A3(new_n781), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n798), .A3(new_n784), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT120), .ZN(new_n859));
  INV_X1    g658(.A(new_n298), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n857), .A2(new_n798), .A3(new_n861), .A4(new_n784), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n671), .B1(new_n863), .B2(new_n795), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n675), .B1(new_n864), .B2(new_n800), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n853), .B1(new_n865), .B2(new_n802), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n850), .B1(new_n852), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G141gat), .B1(new_n867), .B2(new_n298), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  AND4_X1   g668(.A1(new_n359), .A2(new_n814), .A3(new_n553), .A4(new_n532), .ZN(new_n870));
  INV_X1    g669(.A(G141gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n871), .A3(new_n860), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n868), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n873), .A2(KEYINPUT121), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(KEYINPUT121), .ZN(new_n875));
  OAI21_X1  g674(.A(G141gat), .B1(new_n867), .B2(new_n683), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(new_n872), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n874), .B(new_n875), .C1(new_n869), .C2(new_n877), .ZN(G1344gat));
  INV_X1    g677(.A(G148gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n870), .A2(new_n879), .A3(new_n638), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n655), .A2(KEYINPUT57), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT122), .B1(new_n864), .B2(new_n800), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884));
  INV_X1    g683(.A(new_n800), .ZN(new_n885));
  INV_X1    g684(.A(new_n795), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n298), .B1(new_n858), .B2(KEYINPUT120), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n862), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n884), .B(new_n885), .C1(new_n888), .C2(new_n671), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n883), .A2(new_n675), .A3(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n616), .A2(new_n860), .A3(new_n638), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n882), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n851), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT57), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n892), .A2(new_n638), .A3(new_n850), .A4(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n881), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n867), .A2(new_n676), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(KEYINPUT59), .A3(new_n879), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n880), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT123), .B(new_n880), .C1(new_n896), .C2(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1345gat));
  OAI21_X1  g702(.A(G155gat), .B1(new_n867), .B2(new_n675), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n870), .A2(new_n313), .A3(new_n615), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  OAI21_X1  g705(.A(G162gat), .B1(new_n867), .B2(new_n589), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n870), .A2(new_n314), .A3(new_n671), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n553), .A2(new_n663), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n803), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(new_n810), .ZN(new_n912));
  AOI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n684), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n911), .A2(new_n804), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n298), .A2(new_n415), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(G1348gat));
  NAND3_X1  g715(.A1(new_n914), .A2(G176gat), .A3(new_n638), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT124), .Z(new_n918));
  AOI21_X1  g717(.A(G176gat), .B1(new_n912), .B2(new_n638), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(G1349gat));
  NAND2_X1  g719(.A1(new_n914), .A2(new_n615), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n615), .A2(new_n423), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n921), .A2(G183gat), .B1(new_n912), .B2(new_n922), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT60), .Z(G1350gat));
  NAND2_X1  g723(.A1(new_n914), .A2(new_n671), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n424), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n912), .A2(new_n424), .A3(new_n671), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(G1351gat));
  AND3_X1   g731(.A1(new_n851), .A2(new_n532), .A3(new_n910), .ZN(new_n933));
  AOI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n684), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n892), .A2(new_n532), .A3(new_n894), .A4(new_n910), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n860), .A2(G197gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1352gat));
  INV_X1    g737(.A(G204gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n933), .A2(new_n939), .A3(new_n638), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT126), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n892), .A2(new_n894), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n532), .A2(new_n910), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n945), .A2(new_n676), .A3(new_n946), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n943), .B(new_n944), .C1(new_n947), .C2(new_n939), .ZN(G1353gat));
  NOR2_X1   g747(.A1(new_n935), .A2(new_n675), .ZN(new_n949));
  INV_X1    g748(.A(G211gat), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(KEYINPUT127), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n951), .A2(KEYINPUT127), .ZN(new_n954));
  OR3_X1    g753(.A1(new_n949), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n949), .B2(new_n953), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n933), .A2(new_n300), .A3(new_n615), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n935), .B2(new_n589), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n933), .A2(new_n301), .A3(new_n671), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1355gat));
endmodule


