//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1212, new_n1213,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1261, new_n1262;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND3_X1  g0009(.A1(new_n207), .A2(G20), .A3(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT0), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n210), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G116), .A2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G50), .A2(G226), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n226), .B(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n225), .B(new_n230), .C1(G97), .C2(G257), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n213), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT1), .Z(new_n233));
  AOI211_X1 g0033(.A(new_n219), .B(new_n233), .C1(new_n218), .C2(new_n217), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  INV_X1    g0043(.A(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT65), .B(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G222), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT66), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n254), .B1(new_n221), .B2(new_n252), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n209), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n264), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT9), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n213), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n208), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n211), .B2(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G50), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n214), .A2(new_n212), .A3(G1), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  XOR2_X1   g0079(.A(KEYINPUT8), .B(G58), .Z(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n212), .A2(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR3_X1   g0084(.A1(KEYINPUT67), .A2(G20), .A3(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n281), .A2(new_n282), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(G20), .B2(new_n203), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n209), .B1(new_n213), .B2(G33), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n277), .B1(G50), .B2(new_n279), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n272), .A2(G190), .B1(new_n273), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT72), .B1(new_n272), .B2(new_n293), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n291), .A2(new_n273), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT72), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n271), .A2(new_n296), .A3(G200), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n292), .A2(new_n294), .A3(new_n295), .A4(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  OR3_X1    g0099(.A1(new_n298), .A2(KEYINPUT73), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT73), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n298), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n276), .A2(G77), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT71), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n278), .A2(new_n221), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT69), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT15), .B(G87), .Z(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n310), .B2(new_n282), .ZN(new_n311));
  INV_X1    g0111(.A(new_n286), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n280), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G20), .A2(G77), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n309), .A2(KEYINPUT69), .A3(new_n212), .A4(G33), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n311), .A2(new_n313), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n316), .A2(KEYINPUT70), .A3(new_n275), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT70), .B1(new_n316), .B2(new_n275), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n306), .B(new_n307), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n252), .A2(G232), .A3(new_n253), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n257), .B2(new_n229), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT68), .B(G107), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n252), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n263), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n266), .A2(G244), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n325), .A2(new_n270), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n319), .B1(G190), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n325), .A2(new_n270), .A3(new_n326), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G200), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G179), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n272), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n333), .B(new_n291), .C1(G169), .C2(new_n272), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n300), .A2(new_n304), .A3(new_n331), .A4(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT17), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT79), .ZN(new_n337));
  INV_X1    g0137(.A(G58), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(new_n228), .ZN(new_n339));
  OAI21_X1  g0139(.A(G20), .B1(new_n339), .B2(new_n201), .ZN(new_n340));
  INV_X1    g0140(.A(G159), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n286), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT3), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT78), .B1(new_n344), .B2(G33), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(G33), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(KEYINPUT78), .A3(G33), .ZN(new_n348));
  AOI21_X1  g0148(.A(G20), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  OAI21_X1  g0150(.A(G68), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI211_X1 g0151(.A(KEYINPUT7), .B(G20), .C1(new_n347), .C2(new_n348), .ZN(new_n352));
  OAI211_X1 g0152(.A(KEYINPUT16), .B(new_n343), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT16), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n350), .B1(new_n252), .B2(G20), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n346), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n228), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n355), .B1(new_n360), .B2(new_n342), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n275), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n337), .B1(new_n354), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n279), .A2(new_n280), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n276), .B2(new_n280), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n353), .A2(KEYINPUT79), .A3(new_n275), .A4(new_n361), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n269), .B1(new_n266), .B2(G232), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n348), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n346), .B2(new_n345), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n371), .A2(KEYINPUT80), .A3(G226), .A4(G1698), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(G223), .A3(new_n253), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n347), .A2(new_n348), .A3(G226), .A4(G1698), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT80), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n372), .A2(new_n373), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n369), .B1(new_n378), .B2(new_n263), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(G200), .ZN(new_n380));
  AOI211_X1 g0180(.A(G190), .B(new_n369), .C1(new_n378), .C2(new_n263), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n336), .B1(new_n367), .B2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n363), .A2(new_n366), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(G200), .B2(new_n379), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n384), .A2(KEYINPUT17), .A3(new_n365), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n378), .A2(new_n263), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(G179), .A3(new_n368), .ZN(new_n390));
  INV_X1    g0190(.A(G169), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(new_n379), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n367), .A2(KEYINPUT18), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT18), .B1(new_n367), .B2(new_n392), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n383), .B(new_n388), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT76), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n269), .B(KEYINPUT74), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n266), .A2(G238), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G97), .ZN(new_n399));
  INV_X1    g0199(.A(G232), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G1698), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(G226), .B2(G1698), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n399), .B1(new_n402), .B2(new_n358), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n263), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n397), .A2(new_n398), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT13), .ZN(new_n406));
  AOI22_X1  g0206(.A1(G238), .A2(new_n266), .B1(new_n403), .B2(new_n263), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT13), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(new_n397), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n391), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n396), .B1(new_n410), .B2(KEYINPUT77), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT14), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n406), .A2(new_n409), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G179), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n410), .B2(new_n396), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n412), .B(new_n415), .C1(new_n411), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n228), .A2(G20), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n419), .B1(new_n221), .B2(new_n282), .C1(new_n286), .C2(new_n202), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(KEYINPUT11), .A3(new_n275), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n276), .A2(G68), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n419), .A2(G1), .A3(new_n214), .ZN(new_n424));
  XOR2_X1   g0224(.A(new_n424), .B(KEYINPUT12), .Z(new_n425));
  AND2_X1   g0225(.A1(new_n420), .A2(new_n275), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n423), .B(new_n425), .C1(KEYINPUT11), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT75), .B1(new_n413), .B2(new_n385), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT75), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n406), .A2(new_n409), .A3(new_n430), .A4(G190), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n427), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n413), .A2(G200), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n327), .A2(new_n332), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n329), .A2(new_n391), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n319), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n428), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n335), .A2(new_n395), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT4), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n347), .A2(new_n348), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n440), .B1(new_n441), .B2(new_n222), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G283), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n253), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT4), .B1(new_n358), .B2(new_n224), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G1698), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n442), .A2(new_n443), .A3(new_n444), .A4(new_n446), .ZN(new_n447));
  XOR2_X1   g0247(.A(KEYINPUT5), .B(G41), .Z(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n262), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n211), .A2(G45), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n262), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n447), .A2(new_n263), .B1(G257), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n211), .A2(G45), .A3(G274), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G200), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n279), .A2(G97), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n290), .B(new_n279), .C1(G1), .C2(new_n260), .ZN(new_n460));
  INV_X1    g0260(.A(G97), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT6), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(G97), .A2(G107), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(KEYINPUT6), .A3(G97), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n212), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n323), .B1(new_n356), .B2(new_n359), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n286), .A2(new_n221), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n459), .B(new_n463), .C1(new_n474), .C2(new_n290), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n453), .A2(G190), .A3(new_n455), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n457), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT81), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n441), .A2(G20), .A3(new_n228), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n399), .A2(KEYINPUT19), .A3(G20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n399), .A2(new_n212), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n223), .A2(new_n461), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n322), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n482), .B1(new_n485), .B2(KEYINPUT19), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n275), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n310), .A2(new_n278), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n260), .A2(new_n261), .ZN(new_n490));
  OAI211_X1 g0290(.A(G250), .B(new_n450), .C1(new_n490), .C2(new_n208), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n454), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(KEYINPUT82), .A3(new_n454), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n229), .A2(new_n253), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n222), .A2(G1698), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n347), .A2(new_n348), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G116), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n263), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G200), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n494), .A2(new_n495), .B1(new_n501), .B2(new_n263), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G190), .ZN(new_n506));
  INV_X1    g0306(.A(new_n460), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G87), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n489), .A2(new_n504), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n487), .B(new_n488), .C1(new_n310), .C2(new_n460), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n505), .A2(new_n332), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n503), .A2(new_n391), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n456), .A2(new_n391), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n453), .A2(new_n332), .A3(new_n455), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n475), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n457), .A2(new_n476), .A3(KEYINPUT81), .A4(new_n477), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n480), .A2(new_n515), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT86), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n278), .B(new_n465), .C1(new_n521), .C2(KEYINPUT25), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(KEYINPUT25), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n460), .A2(new_n465), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n212), .A2(KEYINPUT23), .A3(G107), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT23), .B1(new_n322), .B2(new_n212), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT85), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT85), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n528), .B(KEYINPUT23), .C1(new_n322), .C2(new_n212), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n347), .A2(new_n348), .A3(new_n212), .A4(G87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT22), .ZN(new_n532));
  XOR2_X1   g0332(.A(KEYINPUT84), .B(KEYINPUT22), .Z(new_n533));
  NAND4_X1  g0333(.A1(new_n533), .A2(new_n212), .A3(G87), .A4(new_n252), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n212), .A2(G33), .A3(G116), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT24), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT24), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n530), .A2(new_n535), .A3(new_n539), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n524), .B1(new_n541), .B2(new_n275), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n523), .B1(new_n279), .B2(G107), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(G257), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G1698), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n224), .A2(new_n253), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n347), .A2(new_n348), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G294), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n260), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n263), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n452), .A2(G264), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n455), .A3(new_n552), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n553), .A2(KEYINPUT87), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(KEYINPUT87), .ZN(new_n555));
  OAI21_X1  g0355(.A(G169), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n553), .A2(new_n332), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n544), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n554), .A2(new_n555), .A3(G190), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n553), .A2(new_n293), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n543), .B(new_n542), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n260), .A2(G97), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n212), .A3(new_n443), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n290), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n244), .A2(G20), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n566), .A2(KEYINPUT83), .A3(new_n212), .A4(new_n443), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n568), .A2(KEYINPUT20), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n565), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n275), .A2(new_n572), .A3(new_n569), .A4(new_n570), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT20), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n571), .A2(new_n575), .B1(G116), .B2(new_n507), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n278), .A2(new_n244), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n545), .A2(new_n253), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n371), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n253), .A2(G264), .ZN(new_n581));
  INV_X1    g0381(.A(G303), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n580), .A2(new_n581), .B1(new_n582), .B2(new_n252), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n263), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n452), .A2(G270), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n455), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n578), .A2(new_n332), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n391), .B1(new_n576), .B2(new_n577), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n586), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT21), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(new_n591), .A3(new_n586), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n587), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n586), .A2(G200), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n594), .B(new_n578), .C1(new_n385), .C2(new_n586), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n520), .A2(new_n564), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n439), .A2(new_n597), .ZN(G372));
  INV_X1    g0398(.A(new_n513), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n517), .A2(new_n475), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n515), .A2(KEYINPUT26), .A3(new_n516), .A4(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT26), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n518), .B2(new_n514), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n599), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n542), .A2(new_n543), .B1(new_n556), .B2(new_n558), .ZN(new_n605));
  INV_X1    g0405(.A(new_n586), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n576), .A2(new_n577), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(G179), .A3(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n588), .A2(new_n591), .A3(new_n586), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n591), .B1(new_n588), .B2(new_n586), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n563), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n604), .B1(new_n612), .B2(new_n520), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n439), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n334), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT88), .ZN(new_n616));
  INV_X1    g0416(.A(new_n304), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n302), .B1(new_n298), .B2(new_n303), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n300), .A2(KEYINPUT88), .A3(new_n304), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n434), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n428), .B2(new_n437), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(new_n383), .A3(new_n388), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n393), .A2(new_n394), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n615), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n614), .A2(new_n628), .ZN(G369));
  INV_X1    g0429(.A(new_n596), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n214), .A2(G20), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n211), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n607), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n593), .B2(new_n638), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT89), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G330), .ZN(new_n643));
  INV_X1    g0443(.A(new_n564), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n544), .A2(new_n637), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT90), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n605), .A2(new_n637), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n646), .B(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n593), .A2(new_n637), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n560), .B2(new_n637), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n650), .A2(new_n655), .ZN(G399));
  NOR2_X1   g0456(.A1(new_n215), .A2(G41), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n207), .ZN(new_n658));
  INV_X1    g0458(.A(new_n657), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G1), .ZN(new_n660));
  OR3_X1    g0460(.A1(new_n322), .A2(G116), .A3(new_n484), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT28), .ZN(new_n663));
  INV_X1    g0463(.A(new_n637), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n613), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT29), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n453), .A2(new_n505), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n668), .A2(new_n606), .A3(KEYINPUT30), .A4(new_n557), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT30), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n583), .A2(new_n263), .B1(G270), .B2(new_n452), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n551), .A2(new_n552), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(G179), .A4(new_n455), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n453), .A2(new_n505), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n670), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n456), .A2(new_n332), .A3(new_n586), .A4(new_n553), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n669), .B(new_n675), .C1(new_n505), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n637), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT31), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n680), .A2(KEYINPUT91), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT91), .B1(new_n680), .B2(new_n681), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR4_X1   g0484(.A1(new_n564), .A2(new_n520), .A3(new_n596), .A4(new_n637), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n667), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n663), .B1(new_n690), .B2(G1), .ZN(G364));
  INV_X1    g0491(.A(KEYINPUT92), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n643), .B(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n660), .B1(G45), .B2(new_n631), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n693), .B(new_n695), .C1(G330), .C2(new_n642), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n385), .A2(G20), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT95), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n699), .A2(G179), .A3(new_n293), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT97), .Z(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G283), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT94), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n212), .A2(new_n332), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G190), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n703), .B1(new_n705), .B2(G200), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n705), .A2(new_n703), .A3(G200), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G322), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n705), .A2(new_n293), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n332), .A2(new_n293), .A3(G190), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G20), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n711), .A2(G326), .B1(G294), .B2(new_n713), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n709), .A2(new_n710), .B1(KEYINPUT98), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(KEYINPUT98), .B2(new_n714), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n293), .A2(G179), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(G20), .A3(G190), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G303), .ZN(new_n720));
  INV_X1    g0520(.A(G311), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n704), .A2(new_n385), .A3(new_n293), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n704), .A2(new_n385), .A3(G200), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT33), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(new_n725), .B2(G317), .ZN(new_n726));
  INV_X1    g0526(.A(G317), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(KEYINPUT33), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n358), .B1(new_n721), .B2(new_n722), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n699), .A2(G179), .A3(G200), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(G329), .B2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n702), .A2(new_n716), .A3(new_n720), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(G159), .ZN(new_n733));
  XNOR2_X1  g0533(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n733), .B(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n709), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(G58), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n701), .A2(G107), .ZN(new_n738));
  INV_X1    g0538(.A(new_n711), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n739), .A2(new_n202), .B1(new_n228), .B2(new_n723), .ZN(new_n740));
  INV_X1    g0540(.A(new_n713), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n461), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n718), .A2(new_n223), .ZN(new_n743));
  NOR4_X1   g0543(.A1(new_n740), .A2(new_n742), .A3(new_n743), .A4(new_n358), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n737), .A2(new_n738), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n722), .A2(new_n221), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n732), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XOR2_X1   g0547(.A(KEYINPUT93), .B(G169), .Z(new_n748));
  AOI21_X1  g0548(.A(new_n208), .B1(new_n748), .B2(G20), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n371), .A2(new_n215), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G45), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n755), .B1(new_n756), .B2(new_n207), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n250), .A2(G45), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n757), .A2(new_n758), .B1(new_n244), .B2(new_n215), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n216), .A2(G355), .A3(new_n252), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n747), .A2(new_n749), .B1(new_n753), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n752), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n694), .B(new_n762), .C1(new_n640), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n696), .A2(new_n764), .ZN(G396));
  NAND4_X1  g0565(.A1(new_n435), .A2(new_n319), .A3(new_n436), .A4(new_n664), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n319), .A2(new_n637), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n331), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n767), .B1(new_n770), .B2(new_n437), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n613), .A2(new_n771), .A3(new_n664), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(KEYINPUT101), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n768), .B1(new_n328), .B2(new_n330), .ZN(new_n774));
  INV_X1    g0574(.A(new_n437), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n766), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n665), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT101), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n613), .A2(new_n771), .A3(new_n778), .A4(new_n664), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n773), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n688), .B(new_n780), .Z(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n695), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n701), .A2(G87), .ZN(new_n783));
  INV_X1    g0583(.A(new_n730), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n721), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n722), .A2(new_n244), .B1(new_n723), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n358), .B1(new_n718), .B2(new_n465), .ZN(new_n788));
  NOR4_X1   g0588(.A1(new_n785), .A2(new_n742), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n711), .A2(G303), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n736), .A2(G294), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n783), .A2(new_n789), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n722), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n724), .A2(G150), .B1(new_n793), .B2(G159), .ZN(new_n794));
  INV_X1    g0594(.A(G137), .ZN(new_n795));
  INV_X1    g0595(.A(G143), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n794), .B1(new_n795), .B2(new_n739), .C1(new_n709), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n701), .A2(G68), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n371), .B1(new_n338), .B2(new_n741), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n730), .B2(G132), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n799), .A2(new_n800), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n718), .A2(new_n202), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n792), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n749), .A2(new_n750), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT99), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n806), .A2(new_n749), .B1(new_n221), .B2(new_n808), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n694), .B(new_n809), .C1(new_n771), .C2(new_n751), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n782), .A2(new_n810), .ZN(G384));
  AND3_X1   g0611(.A1(new_n480), .A2(new_n518), .A3(new_n519), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n644), .A2(new_n630), .A3(new_n515), .A4(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n680), .B(new_n681), .C1(new_n813), .C2(new_n637), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n439), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT106), .Z(new_n816));
  INV_X1    g0616(.A(new_n635), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n367), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n395), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT103), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n384), .A2(new_n365), .A3(new_n387), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT37), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n367), .B1(new_n392), .B2(new_n817), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n823), .B1(new_n822), .B2(new_n824), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n395), .A2(KEYINPUT103), .A3(new_n818), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n821), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT38), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n822), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n343), .B1(new_n351), .B2(new_n352), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n355), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n835), .A2(new_n275), .A3(new_n353), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n836), .A2(new_n365), .ZN(new_n837));
  INV_X1    g0637(.A(new_n392), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n838), .B2(new_n635), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT37), .B1(new_n833), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n825), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT102), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n837), .A2(new_n635), .ZN(new_n843));
  AND3_X1   g0643(.A1(new_n395), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n842), .B1(new_n395), .B2(new_n843), .ZN(new_n845));
  OAI211_X1 g0645(.A(KEYINPUT38), .B(new_n841), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n832), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n427), .A2(new_n637), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n428), .A2(new_n434), .A3(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n427), .B(new_n637), .C1(new_n622), .C2(new_n418), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n776), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n680), .A2(new_n681), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n685), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n847), .A2(KEYINPUT40), .A3(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n395), .A2(new_n843), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT102), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n395), .A2(new_n842), .A3(new_n843), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n860), .B2(new_n841), .ZN(new_n861));
  INV_X1    g0661(.A(new_n846), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n854), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT105), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT40), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n831), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n853), .B1(new_n868), .B2(new_n846), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT105), .B1(new_n869), .B2(KEYINPUT40), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n856), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n816), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(G330), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n666), .A2(new_n439), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n628), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT104), .Z(new_n876));
  XNOR2_X1  g0676(.A(new_n873), .B(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n626), .A2(new_n817), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n773), .A2(new_n766), .A3(new_n779), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n849), .A2(new_n850), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n861), .A2(new_n862), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n428), .A2(new_n637), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT39), .B1(new_n832), .B2(new_n846), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(KEYINPUT39), .B2(new_n882), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n878), .B(new_n883), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n877), .B(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n211), .B2(new_n631), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT35), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n212), .B(new_n208), .C1(new_n470), .C2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(G116), .C1(new_n890), .C2(new_n470), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT36), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n207), .B(G77), .C1(new_n338), .C2(new_n228), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(G50), .B2(new_n228), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(G1), .A3(new_n214), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n889), .A2(new_n893), .A3(new_n896), .ZN(G367));
  OAI21_X1  g0697(.A(new_n812), .B1(new_n476), .B2(new_n664), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n654), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT42), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n518), .B1(new_n898), .B2(new_n560), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n664), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n489), .A2(new_n508), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n637), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n515), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n599), .A2(new_n904), .A3(new_n637), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n909));
  XOR2_X1   g0709(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n910));
  NAND3_X1  g0710(.A1(new_n906), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n903), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n911), .B2(new_n903), .ZN(new_n913));
  INV_X1    g0713(.A(new_n650), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n600), .A2(new_n516), .A3(new_n637), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n898), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n913), .B(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n657), .B(KEYINPUT41), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n655), .A2(new_n916), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT45), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n655), .A2(new_n916), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT44), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n914), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n922), .A2(new_n914), .A3(new_n925), .ZN(new_n928));
  INV_X1    g0728(.A(new_n649), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n654), .B1(new_n929), .B2(new_n653), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(new_n643), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n693), .B2(new_n930), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n927), .A2(new_n690), .A3(new_n928), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n920), .B1(new_n933), .B2(new_n690), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n211), .B1(new_n631), .B2(G45), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT108), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n918), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n252), .B1(new_n739), .B2(new_n796), .C1(new_n784), .C2(new_n795), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(G77), .B2(new_n700), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n793), .A2(G50), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n719), .A2(G58), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n741), .A2(new_n228), .B1(new_n723), .B2(new_n341), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n736), .B2(G150), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n739), .A2(new_n721), .B1(new_n323), .B2(new_n741), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n736), .B2(G303), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT46), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n718), .B2(new_n244), .ZN(new_n948));
  AOI22_X1  g0748(.A1(G97), .A2(new_n700), .B1(new_n730), .B2(G317), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n718), .A2(new_n947), .A3(new_n244), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n371), .B(new_n950), .C1(G294), .C2(new_n724), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n946), .A2(new_n948), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n722), .A2(new_n786), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n944), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT47), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n695), .B1(new_n955), .B2(new_n749), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n753), .B1(new_n216), .B2(new_n310), .C1(new_n755), .C2(new_n241), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT109), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n956), .B(new_n958), .C1(new_n763), .C2(new_n908), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n937), .A2(new_n959), .ZN(G387));
  OR2_X1    g0760(.A1(new_n932), .A2(new_n690), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n932), .A2(new_n690), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(new_n657), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n932), .A2(new_n936), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n661), .A2(new_n216), .A3(new_n252), .ZN(new_n965));
  AOI21_X1  g0765(.A(G45), .B1(new_n661), .B2(KEYINPUT110), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(KEYINPUT110), .B2(new_n661), .C1(new_n228), .C2(new_n221), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT111), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n280), .A2(new_n202), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT50), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n754), .B1(new_n238), .B2(new_n756), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n965), .B1(G107), .B2(new_n216), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n695), .B1(new_n973), .B2(new_n753), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT112), .ZN(new_n975));
  INV_X1    g0775(.A(new_n749), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n730), .A2(G326), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G322), .A2(new_n711), .B1(new_n724), .B2(G311), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n582), .B2(new_n722), .C1(new_n709), .C2(new_n727), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT48), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n786), .B2(new_n741), .C1(new_n549), .C2(new_n718), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT49), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n371), .B(new_n977), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n700), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n983), .B1(new_n982), .B2(new_n981), .C1(new_n244), .C2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n310), .A2(new_n741), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n736), .B2(G50), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT114), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n701), .A2(G97), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n722), .A2(new_n228), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n371), .B1(new_n221), .B2(new_n718), .C1(new_n281), .C2(new_n723), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(G150), .C2(new_n730), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n711), .A2(G159), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT113), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n988), .A2(new_n989), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n985), .A2(new_n995), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n975), .B1(new_n976), .B2(new_n996), .C1(new_n929), .C2(new_n763), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n963), .A2(new_n964), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT115), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n963), .A2(KEYINPUT115), .A3(new_n964), .A4(new_n997), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(G393));
  NAND3_X1  g0802(.A1(new_n927), .A2(new_n928), .A3(new_n936), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n916), .A2(new_n752), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n753), .B1(new_n461), .B2(new_n216), .C1(new_n247), .C2(new_n755), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n709), .A2(new_n721), .B1(new_n727), .B2(new_n739), .ZN(new_n1006));
  XOR2_X1   g0806(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n719), .A2(G283), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n358), .B1(new_n723), .B2(new_n582), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n741), .A2(new_n244), .B1(new_n722), .B2(new_n549), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(new_n730), .C2(G322), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n738), .A3(new_n1009), .A4(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n741), .A2(new_n221), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n280), .B2(new_n793), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n202), .B2(new_n723), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n441), .B(new_n1016), .C1(G143), .C2(new_n730), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n709), .A2(new_n341), .B1(new_n287), .B2(new_n739), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT51), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n783), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n718), .A2(new_n228), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1013), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n695), .B1(new_n1024), .B2(new_n749), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1004), .A2(new_n1005), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n928), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n962), .B1(new_n1027), .B2(new_n926), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT117), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n659), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(KEYINPUT117), .B(new_n962), .C1(new_n1027), .C2(new_n926), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n933), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1003), .B(new_n1026), .C1(new_n1031), .C2(new_n1033), .ZN(G390));
  INV_X1    g0834(.A(KEYINPUT118), .ZN(new_n1035));
  INV_X1    g0835(.A(G330), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n776), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n814), .A2(new_n880), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1037), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n684), .B2(new_n686), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1038), .B1(new_n1040), .B2(new_n880), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n879), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n880), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n880), .B1(new_n814), .B2(new_n1037), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n772), .A2(new_n766), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n439), .A2(G330), .A3(new_n814), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n875), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1035), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n885), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n868), .A2(KEYINPUT39), .A3(new_n846), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n884), .B1(new_n879), .B2(new_n880), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n847), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n884), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n880), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n1046), .B2(new_n1060), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1038), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1052), .A2(new_n1053), .B1(new_n881), .B2(new_n1059), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1043), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1051), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1044), .B1(new_n1040), .B2(new_n880), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1069), .A2(new_n1046), .B1(new_n1041), .B2(new_n879), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n874), .B(new_n628), .C1(new_n815), .C2(new_n1036), .ZN(new_n1071));
  OAI21_X1  g0871(.A(KEYINPUT118), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1038), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1062), .B(new_n1043), .C1(new_n886), .C2(new_n1055), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1068), .A2(new_n657), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n936), .ZN(new_n1078));
  INV_X1    g0878(.A(G125), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n252), .B1(new_n984), .B2(new_n202), .C1(new_n1079), .C2(new_n784), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT119), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT53), .B1(new_n718), .B2(new_n287), .ZN(new_n1082));
  INV_X1    g0882(.A(G128), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1082), .B1(new_n739), .B2(new_n1083), .ZN(new_n1084));
  OR3_X1    g0884(.A1(new_n718), .A2(KEYINPUT53), .A3(new_n287), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT54), .B(G143), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1085), .B1(new_n795), .B2(new_n723), .C1(new_n722), .C2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1084), .B(new_n1087), .C1(G132), .C2(new_n736), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1081), .B(new_n1088), .C1(new_n341), .C2(new_n741), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G283), .A2(new_n711), .B1(new_n724), .B2(new_n322), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n461), .B2(new_n722), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1014), .B(new_n1091), .C1(G116), .C2(new_n736), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n743), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n252), .B1(new_n730), .B2(G294), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n801), .A4(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n976), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n695), .B(new_n1096), .C1(new_n281), .C2(new_n808), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT120), .Z(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n886), .B2(new_n751), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1077), .A2(new_n1078), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(G378));
  INV_X1    g0901(.A(KEYINPUT57), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1074), .A2(new_n1075), .A3(new_n1048), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n1050), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n869), .A2(KEYINPUT105), .A3(KEYINPUT40), .ZN(new_n1106));
  OAI211_X1 g0906(.A(G330), .B(new_n855), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n621), .A2(new_n334), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT55), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT55), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n621), .A2(new_n1110), .A3(new_n334), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n291), .A2(new_n817), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT56), .Z(new_n1113));
  NAND3_X1  g0913(.A1(new_n1109), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1113), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1110), .B1(new_n621), .B2(new_n334), .ZN(new_n1116));
  AOI211_X1 g0916(.A(KEYINPUT55), .B(new_n615), .C1(new_n619), .C2(new_n620), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1107), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n871), .A2(G330), .A3(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1120), .A2(new_n887), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n887), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1104), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n878), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(new_n882), .B2(new_n881), .C1(new_n1054), .C2(new_n1059), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1107), .A2(new_n1119), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1121), .B1(new_n871), .B2(G330), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1120), .A2(new_n887), .A3(new_n1122), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(KEYINPUT125), .A3(new_n1104), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1127), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1129), .A2(KEYINPUT123), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1120), .A2(new_n1122), .A3(KEYINPUT123), .A4(new_n1129), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1103), .A2(new_n1050), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1102), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n657), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1138), .A2(new_n936), .A3(new_n1139), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1119), .A2(new_n750), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n807), .A2(new_n202), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n441), .A2(new_n261), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G58), .A2(new_n700), .B1(new_n730), .B2(G283), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n228), .B2(new_n741), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1147), .B(new_n1149), .C1(G77), .C2(new_n719), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n739), .A2(new_n244), .B1(new_n461), .B2(new_n723), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n736), .B2(G107), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(new_n310), .C2(new_n722), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT58), .ZN(new_n1154));
  INV_X1    g0954(.A(G132), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n722), .A2(new_n795), .B1(new_n723), .B2(new_n1155), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n739), .A2(new_n1079), .B1(new_n718), .B2(new_n1086), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(new_n736), .C2(G128), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n287), .B2(new_n741), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n730), .A2(G124), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(G33), .A2(G41), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT121), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n700), .B2(G159), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1147), .A2(new_n202), .A3(new_n1164), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1154), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n695), .B1(new_n1168), .B2(new_n749), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1145), .A2(new_n1146), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT122), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT122), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1145), .A2(new_n1172), .A3(new_n1146), .A4(new_n1169), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT124), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1144), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1144), .B2(new_n1174), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1136), .A2(new_n1143), .B1(new_n1176), .B2(new_n1177), .ZN(G375));
  NAND2_X1  g0978(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n1180), .A3(new_n919), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1060), .A2(new_n750), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1086), .A2(new_n723), .B1(new_n722), .B2(new_n287), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n741), .A2(new_n202), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n736), .C2(G137), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n711), .A2(G132), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n441), .B1(G159), .B2(new_n719), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G58), .A2(new_n700), .B1(new_n730), .B2(G128), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n701), .A2(G77), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n784), .A2(new_n582), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n739), .A2(new_n549), .B1(new_n244), .B2(new_n723), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n358), .B1(new_n718), .B2(new_n461), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n986), .A4(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1190), .B(new_n1194), .C1(new_n786), .C2(new_n709), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n323), .A2(new_n722), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1189), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1197), .A2(new_n749), .B1(new_n228), .B2(new_n808), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1182), .A2(new_n694), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1048), .B2(new_n936), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1181), .A2(new_n1200), .ZN(G381));
  INV_X1    g1001(.A(new_n1026), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1033), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1202), .B1(new_n1203), .B2(new_n1030), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1204), .A2(new_n937), .A3(new_n959), .A4(new_n1003), .ZN(new_n1205));
  INV_X1    g1005(.A(G396), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1000), .A2(new_n1206), .A3(new_n1001), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(G375), .A2(G378), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(G381), .A2(G384), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(G407));
  NAND2_X1  g1011(.A1(new_n636), .A2(G213), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(G375), .A2(G378), .A3(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT126), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1015(.A(KEYINPUT60), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1180), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n1071), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1217), .A2(new_n657), .A3(new_n1179), .A4(new_n1218), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1219), .A2(G384), .A3(new_n1200), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G384), .B1(new_n1219), .B2(new_n1200), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n919), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1134), .A2(new_n936), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1100), .A2(new_n1174), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1212), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G375), .B2(G378), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n636), .A2(G213), .A3(G2897), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1223), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT62), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1177), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1144), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1127), .A2(new_n1142), .A3(new_n1135), .A4(new_n657), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1100), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1222), .B(new_n1229), .C1(new_n1237), .C2(new_n1227), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1231), .A2(new_n1232), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1228), .A2(new_n1222), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT61), .B1(new_n1240), .B2(KEYINPUT62), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT127), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G387), .A2(G390), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1205), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G393), .A2(G396), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1247), .A2(new_n1207), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1207), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n1245), .A3(new_n1205), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1239), .A2(KEYINPUT127), .A3(new_n1241), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1244), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT63), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1252), .B1(new_n1255), .B2(new_n1240), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1231), .A2(KEYINPUT63), .A3(new_n1238), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1254), .A2(new_n1259), .ZN(G405));
  NOR2_X1   g1060(.A1(new_n1209), .A2(new_n1237), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(new_n1222), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(new_n1252), .ZN(G402));
endmodule


