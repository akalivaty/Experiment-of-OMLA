//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(new_n189), .A3(G143), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  XNOR2_X1  g014(.A(G143), .B(G146), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT68), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n201), .A2(KEYINPUT68), .A3(new_n203), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n199), .B(new_n200), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT88), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n196), .A2(new_n210), .B1(new_n201), .B2(new_n208), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(new_n200), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n206), .A2(KEYINPUT88), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G224), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G953), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n217), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n213), .A2(new_n219), .A3(new_n214), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G110), .B(G122), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(KEYINPUT85), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT83), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT2), .B(G113), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT71), .B1(new_n227), .B2(G119), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT70), .B(G116), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G119), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(KEYINPUT70), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G116), .ZN(new_n234));
  AND4_X1   g048(.A1(new_n231), .A2(new_n232), .A3(new_n234), .A4(G119), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n226), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT3), .B1(new_n237), .B2(G107), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n239));
  INV_X1    g053(.A(G107), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(G104), .ZN(new_n241));
  INV_X1    g055(.A(G101), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(G107), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n238), .A2(new_n241), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n237), .A2(G107), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n240), .A2(G104), .ZN(new_n246));
  OAI21_X1  g060(.A(G101), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n236), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT5), .ZN(new_n251));
  INV_X1    g065(.A(G119), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(G116), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G113), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n232), .A2(new_n234), .A3(G119), .ZN(new_n255));
  INV_X1    g069(.A(new_n228), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n232), .A2(new_n234), .A3(new_n231), .A4(G119), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n254), .B1(new_n259), .B2(KEYINPUT5), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n224), .B1(new_n250), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G101), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT4), .A3(new_n244), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n265), .A3(G101), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n230), .A2(new_n235), .A3(new_n226), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n225), .B1(new_n257), .B2(new_n258), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n264), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT5), .B1(new_n230), .B2(new_n235), .ZN(new_n270));
  INV_X1    g084(.A(new_n254), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n248), .B1(new_n259), .B2(new_n226), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT83), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n261), .A2(new_n269), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT84), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n223), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n261), .A2(KEYINPUT84), .A3(new_n274), .A4(new_n269), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT87), .B(KEYINPUT6), .Z(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n274), .A2(new_n269), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT83), .B1(new_n272), .B2(new_n273), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n223), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(KEYINPUT86), .A3(new_n278), .A4(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n261), .A2(new_n269), .A3(new_n274), .A4(new_n222), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n286), .A2(KEYINPUT6), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT86), .B1(new_n277), .B2(new_n278), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n221), .B(new_n280), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT89), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n283), .A2(new_n278), .A3(new_n284), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT86), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n285), .A3(new_n287), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n296), .A2(KEYINPUT89), .A3(new_n221), .A4(new_n280), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT7), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n219), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n218), .A2(new_n220), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n222), .B(KEYINPUT8), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n248), .B1(new_n260), .B2(new_n268), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT90), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n272), .A2(new_n273), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n303), .A2(new_n304), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n213), .A2(new_n299), .A3(new_n219), .A4(new_n214), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n301), .A2(new_n286), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n188), .B1(new_n298), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n188), .ZN(new_n316));
  AOI211_X1 g130(.A(new_n316), .B(new_n313), .C1(new_n292), .C2(new_n297), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n187), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT91), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n199), .B1(new_n204), .B2(new_n205), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT11), .ZN(new_n321));
  INV_X1    g135(.A(G134), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(G137), .ZN(new_n323));
  INV_X1    g137(.A(G137), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT11), .A3(G134), .ZN(new_n325));
  INV_X1    g139(.A(G131), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n322), .A2(G137), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n323), .A2(new_n325), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT66), .ZN(new_n329));
  INV_X1    g143(.A(new_n327), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n322), .A2(G137), .ZN(new_n331));
  OAI21_X1  g145(.A(G131), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n320), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT69), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n320), .A2(new_n329), .A3(KEYINPUT69), .A4(new_n332), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n323), .A2(new_n325), .A3(new_n327), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT67), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n323), .A2(new_n325), .A3(new_n339), .A4(new_n327), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(G131), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n329), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n211), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n335), .A2(new_n336), .A3(new_n343), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT72), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n329), .A2(new_n341), .A3(KEYINPUT72), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n211), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(KEYINPUT30), .A3(new_n333), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n267), .A2(new_n268), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n346), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G237), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT73), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G237), .ZN(new_n358));
  AOI21_X1  g172(.A(G953), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G210), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT27), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT26), .B(G101), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n350), .A2(new_n352), .A3(new_n333), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n354), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT31), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n354), .A2(KEYINPUT31), .A3(new_n364), .A4(new_n365), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT28), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n344), .A2(new_n353), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n350), .A2(KEYINPUT28), .A3(new_n352), .A4(new_n333), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n363), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(G472), .A2(G902), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(KEYINPUT32), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n354), .A2(new_n365), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n363), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n372), .A2(new_n364), .A3(new_n373), .A4(new_n374), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n350), .A2(new_n333), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n353), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n363), .A2(new_n382), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n372), .A2(new_n386), .A3(new_n374), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n312), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT74), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(KEYINPUT74), .A3(new_n312), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n384), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G472), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT32), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n368), .A2(new_n369), .B1(new_n363), .B2(new_n375), .ZN(new_n396));
  INV_X1    g210(.A(new_n378), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n379), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT23), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n252), .B2(G128), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n401), .B(new_n402), .C1(G119), .C2(new_n202), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT77), .B(G110), .Z(new_n404));
  XOR2_X1   g218(.A(KEYINPUT24), .B(G110), .Z(new_n405));
  XNOR2_X1  g219(.A(G119), .B(G128), .ZN(new_n406));
  OAI22_X1  g220(.A1(new_n403), .A2(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT16), .ZN(new_n408));
  INV_X1    g222(.A(G140), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(G125), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(G125), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n200), .A2(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g227(.A(G146), .B(new_n410), .C1(new_n413), .C2(new_n408), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n412), .A3(new_n189), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n407), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT76), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n403), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n403), .A2(new_n417), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n418), .A2(G110), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n410), .B1(new_n413), .B2(new_n408), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n189), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n414), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n405), .A2(new_n406), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n416), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G953), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(G221), .A3(G234), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT78), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT22), .B(G137), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n416), .B(new_n431), .C1(new_n420), .C2(new_n425), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT79), .B(KEYINPUT25), .C1(new_n435), .C2(G902), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n312), .B1(KEYINPUT79), .B2(KEYINPUT25), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n433), .B2(new_n434), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT79), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT25), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(G217), .A2(G902), .ZN(new_n442));
  INV_X1    g256(.A(G217), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(G234), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n444), .B(KEYINPUT75), .Z(new_n445));
  NAND3_X1  g259(.A1(new_n436), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n446), .A2(KEYINPUT80), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(KEYINPUT80), .ZN(new_n448));
  INV_X1    g262(.A(new_n435), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n445), .A2(G902), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n447), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n399), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n454), .B(new_n187), .C1(new_n315), .C2(new_n317), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n357), .A2(G237), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n355), .A2(KEYINPUT73), .ZN(new_n457));
  OAI211_X1 g271(.A(G214), .B(new_n427), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n192), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n359), .A2(G143), .A3(G214), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G131), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT17), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n326), .A3(new_n460), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n326), .B1(new_n459), .B2(new_n460), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n423), .B1(new_n466), .B2(KEYINPUT17), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G113), .B(G122), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(new_n237), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n415), .A2(KEYINPUT92), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT93), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n415), .A2(KEYINPUT92), .A3(KEYINPUT93), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n413), .A2(G146), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n473), .A2(G146), .A3(new_n413), .A4(new_n474), .ZN(new_n478));
  AND2_X1   g292(.A1(KEYINPUT18), .A2(G131), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n459), .B2(new_n460), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n459), .A2(new_n460), .A3(new_n479), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n477), .B(new_n478), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n468), .A2(new_n470), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT94), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n468), .A2(KEYINPUT94), .A3(new_n470), .A4(new_n482), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n468), .A2(new_n482), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n487), .B1(new_n470), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n312), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G475), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n462), .A2(new_n464), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n413), .B(KEYINPUT19), .Z(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n492), .B(new_n414), .C1(G146), .C2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n470), .B1(new_n495), .B2(new_n482), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n496), .B1(new_n485), .B2(new_n486), .ZN(new_n497));
  NOR2_X1   g311(.A1(G475), .A2(G902), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n497), .A2(KEYINPUT20), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT95), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT20), .B1(new_n497), .B2(new_n499), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n496), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n499), .B1(new_n487), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n491), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G469), .ZN(new_n510));
  XNOR2_X1  g324(.A(G110), .B(G140), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n427), .A2(G227), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n511), .B(new_n512), .Z(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n264), .A2(new_n211), .A3(new_n266), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n320), .A2(KEYINPUT10), .A3(new_n249), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n201), .A2(new_n203), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n201), .A2(KEYINPUT68), .A3(new_n203), .ZN(new_n520));
  INV_X1    g334(.A(new_n201), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n198), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n519), .A2(new_n520), .B1(new_n522), .B2(KEYINPUT81), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n522), .A2(KEYINPUT81), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n248), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n515), .B(new_n516), .C1(new_n525), .C2(KEYINPUT10), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n348), .A2(new_n349), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n514), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT82), .ZN(new_n529));
  OR3_X1    g343(.A1(new_n320), .A2(new_n529), .A3(new_n249), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n529), .B1(new_n320), .B2(new_n249), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n525), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n342), .A2(KEYINPUT12), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n348), .A2(new_n349), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n535), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n528), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n526), .A2(new_n527), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n526), .A2(new_n527), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n514), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n510), .B(new_n312), .C1(new_n538), .C2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n510), .A2(new_n312), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n528), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n540), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n526), .A2(new_n527), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(new_n534), .B2(new_n537), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n546), .B1(new_n548), .B2(new_n514), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n542), .B(new_n544), .C1(new_n510), .C2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT9), .B(G234), .ZN(new_n551));
  OAI21_X1  g365(.A(G221), .B1(new_n551), .B2(G902), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT13), .B1(new_n202), .B2(G143), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(new_n322), .ZN(new_n555));
  XNOR2_X1  g369(.A(G128), .B(G143), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT96), .B(G122), .Z(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G116), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n229), .A2(G122), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT97), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(KEYINPUT97), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n240), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n564), .A2(new_n240), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n557), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n560), .A2(KEYINPUT14), .B1(new_n558), .B2(G116), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(KEYINPUT14), .B2(new_n560), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G107), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n556), .B(new_n322), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n565), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n551), .A2(new_n443), .A3(G953), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n568), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n574), .B1(new_n568), .B2(new_n573), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n312), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT15), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(G478), .ZN(new_n580));
  INV_X1    g394(.A(G478), .ZN(new_n581));
  OAI221_X1 g395(.A(new_n312), .B1(KEYINPUT15), .B2(new_n581), .C1(new_n576), .C2(new_n577), .ZN(new_n582));
  NAND2_X1  g396(.A1(G234), .A2(G237), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(G952), .A3(new_n427), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(G902), .A3(G953), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT21), .B(G898), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n580), .A2(new_n582), .A3(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n509), .A2(new_n553), .A3(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n319), .A2(new_n453), .A3(new_n455), .A4(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  NAND2_X1  g408(.A1(new_n578), .A2(new_n581), .ZN(new_n595));
  INV_X1    g409(.A(new_n577), .ZN(new_n596));
  NOR2_X1   g410(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n597));
  AND2_X1   g411(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n596), .B(new_n575), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n576), .A2(new_n577), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n599), .B1(new_n600), .B2(new_n598), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n312), .A2(G478), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n595), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n509), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n318), .A2(new_n589), .A3(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n550), .A2(new_n552), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n377), .B(new_n312), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(KEYINPUT98), .B(G472), .C1(new_n396), .C2(G902), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n606), .A2(new_n609), .A3(new_n452), .A4(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT100), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  AND2_X1   g430(.A1(new_n490), .A2(G475), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n502), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(KEYINPUT102), .B(KEYINPUT20), .C1(new_n497), .C2(new_n499), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n505), .B2(new_n506), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n619), .A2(new_n623), .A3(new_n620), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n617), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n580), .A2(new_n582), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n589), .B(KEYINPUT103), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT104), .B1(new_n630), .B2(new_n318), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n619), .A2(new_n623), .A3(new_n620), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n623), .B1(new_n619), .B2(new_n620), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n491), .B(new_n628), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n629), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n187), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n298), .A2(new_n314), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n316), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n298), .A2(new_n188), .A3(new_n314), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n636), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n631), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n612), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  NOR2_X1   g461(.A1(new_n431), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n426), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n450), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n447), .A2(new_n448), .A3(new_n650), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n609), .A2(new_n610), .A3(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n319), .A2(new_n592), .A3(new_n455), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT105), .B(KEYINPUT106), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  AND3_X1   g471(.A1(new_n399), .A2(new_n606), .A3(new_n651), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n585), .B1(new_n587), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n634), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n658), .A2(new_n641), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XOR2_X1   g477(.A(new_n660), .B(KEYINPUT39), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n606), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT40), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n509), .A2(new_n187), .A3(new_n628), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n365), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n352), .B1(new_n350), .B2(new_n333), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n363), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT107), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n673), .B(new_n363), .C1(new_n669), .C2(new_n670), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n672), .A2(new_n366), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n675), .B2(G902), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n379), .A2(new_n398), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n651), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n668), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n315), .A2(new_n317), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT38), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n192), .ZN(G45));
  INV_X1    g498(.A(new_n660), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n603), .A2(new_n509), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n658), .A2(new_n641), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  NOR2_X1   g503(.A1(new_n604), .A2(new_n589), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n538), .A2(new_n541), .ZN(new_n691));
  OAI21_X1  g505(.A(G469), .B1(new_n691), .B2(G902), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n692), .A2(new_n552), .A3(new_n542), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n453), .A2(new_n641), .A3(new_n690), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NAND3_X1  g510(.A1(new_n399), .A2(new_n452), .A3(new_n693), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n631), .B2(new_n643), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT108), .B(G116), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G18));
  NOR2_X1   g514(.A1(new_n509), .A2(new_n591), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n399), .A2(new_n701), .A3(new_n651), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n187), .B(new_n693), .C1(new_n315), .C2(new_n317), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  NOR2_X1   g520(.A1(new_n681), .A2(new_n667), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n372), .A2(new_n374), .A3(new_n386), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n368), .A2(new_n369), .B1(new_n363), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n378), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT109), .B1(new_n709), .B2(new_n397), .ZN(new_n713));
  OAI21_X1  g527(.A(G472), .B1(new_n396), .B2(G902), .ZN(new_n714));
  AND4_X1   g528(.A1(new_n452), .A2(new_n712), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n693), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n635), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n707), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT110), .B(G122), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G24));
  NAND4_X1  g534(.A1(new_n712), .A2(new_n713), .A3(new_n714), .A4(new_n651), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n686), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n704), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n639), .A2(new_n606), .A3(new_n187), .A4(new_n640), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n399), .A2(new_n452), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT42), .B1(new_n728), .B2(new_n687), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n726), .A2(new_n727), .A3(new_n730), .A4(new_n686), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n725), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n315), .A2(new_n317), .A3(new_n553), .A4(new_n637), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n453), .A3(new_n687), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n730), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n728), .A2(KEYINPUT42), .A3(new_n687), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(KEYINPUT111), .A3(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  NAND3_X1  g553(.A1(new_n733), .A2(new_n453), .A3(new_n661), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT112), .B(G134), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G36));
  NAND2_X1  g556(.A1(new_n502), .A2(new_n501), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n505), .A2(new_n506), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n617), .B1(new_n745), .B2(new_n507), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n603), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT114), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n747), .B(KEYINPUT43), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n678), .B1(new_n609), .B2(new_n610), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n750), .A2(new_n753), .A3(KEYINPUT44), .A4(new_n754), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n549), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n510), .B1(new_n549), .B2(new_n759), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n543), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT46), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(KEYINPUT46), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n542), .B(new_n763), .C1(new_n764), .C2(KEYINPUT113), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n764), .A2(KEYINPUT113), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n552), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n664), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n315), .A2(new_n317), .A3(new_n637), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n757), .A2(new_n758), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  NOR4_X1   g587(.A1(new_n770), .A2(new_n399), .A3(new_n452), .A4(new_n686), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT47), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n767), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n767), .A2(new_n775), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  NAND3_X1  g593(.A1(new_n694), .A2(new_n705), .A3(new_n718), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n698), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n628), .A2(new_n660), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n627), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n658), .A2(new_n783), .A3(new_n769), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n733), .A2(new_n722), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n740), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n781), .A2(new_n732), .A3(new_n737), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n553), .A2(new_n660), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n707), .A2(new_n679), .A3(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n662), .A2(new_n688), .A3(new_n723), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT52), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n399), .A2(new_n606), .A3(new_n651), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n318), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n794), .A2(new_n661), .B1(new_n704), .B2(new_n722), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n688), .A4(new_n790), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n788), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n746), .A2(new_n628), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n635), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n319), .A2(new_n455), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT115), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n319), .A2(new_n804), .A3(new_n455), .A4(new_n801), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n612), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n604), .A2(new_n635), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n319), .A2(new_n612), .A3(new_n455), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n593), .A3(new_n653), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n807), .A2(KEYINPUT116), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n611), .B1(new_n803), .B2(new_n805), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n813), .B1(new_n814), .B2(new_n810), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n799), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n662), .A2(new_n723), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT52), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT53), .B1(new_n799), .B2(new_n816), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT54), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT116), .B1(new_n807), .B2(new_n811), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n814), .A2(new_n813), .A3(new_n810), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n786), .A2(new_n780), .A3(new_n698), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n738), .A2(new_n792), .A3(new_n797), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n818), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n792), .A2(new_n797), .ZN(new_n831));
  INV_X1    g645(.A(new_n697), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n644), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n605), .A2(new_n832), .B1(new_n702), .B2(new_n704), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(KEYINPUT117), .A3(new_n718), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n780), .B2(new_n698), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AND4_X1   g652(.A1(KEYINPUT53), .A2(new_n784), .A3(new_n740), .A4(new_n785), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n735), .A2(new_n736), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n839), .A2(new_n840), .A3(new_n820), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n816), .A2(new_n831), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n829), .A2(new_n830), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n823), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n751), .A2(new_n584), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n715), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n703), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT120), .Z(new_n848));
  NOR2_X1   g662(.A1(new_n770), .A2(new_n716), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n727), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT48), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n452), .A2(new_n585), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n770), .A2(new_n677), .A3(new_n716), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n604), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(G952), .A3(new_n427), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n848), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n776), .A2(new_n777), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n692), .A2(new_n542), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n552), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n846), .A2(new_n770), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n693), .A2(new_n637), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT119), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n845), .A2(new_n682), .A3(new_n715), .A4(new_n866), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT50), .Z(new_n868));
  NOR2_X1   g682(.A1(new_n603), .A2(new_n509), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n854), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n850), .B2(new_n721), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n864), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n861), .A2(new_n552), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT118), .Z(new_n876));
  NAND2_X1  g690(.A1(new_n859), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n871), .B1(new_n877), .B2(new_n863), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n878), .A2(new_n868), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n858), .B(new_n874), .C1(KEYINPUT51), .C2(new_n879), .ZN(new_n880));
  OAI22_X1  g694(.A1(new_n844), .A2(new_n880), .B1(G952), .B2(G953), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n861), .A2(KEYINPUT49), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n452), .A3(new_n187), .A4(new_n552), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n861), .A2(KEYINPUT49), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n883), .A2(new_n677), .A3(new_n884), .A4(new_n747), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n682), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n881), .A2(new_n886), .ZN(G75));
  NAND2_X1  g701(.A1(new_n829), .A2(new_n842), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(G210), .A3(G902), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n296), .A2(new_n280), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(new_n221), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT55), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n889), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n889), .B2(new_n890), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n427), .A2(G952), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G51));
  AND4_X1   g711(.A1(G902), .A2(new_n888), .A3(new_n760), .A4(new_n761), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n831), .A2(new_n838), .A3(new_n841), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n826), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT54), .B1(new_n900), .B2(new_n822), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n843), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n543), .B(KEYINPUT57), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n691), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n898), .B1(new_n904), .B2(KEYINPUT121), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n906));
  INV_X1    g720(.A(new_n903), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n901), .B2(new_n843), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n908), .B2(new_n691), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n896), .B1(new_n905), .B2(new_n909), .ZN(G54));
  NAND4_X1  g724(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n911), .A2(KEYINPUT122), .A3(new_n497), .ZN(new_n912));
  INV_X1    g726(.A(new_n896), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n911), .B2(new_n497), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT122), .B1(new_n911), .B2(new_n497), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(G60));
  INV_X1    g730(.A(new_n601), .ZN(new_n917));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT59), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n844), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n902), .A2(new_n917), .A3(new_n919), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n896), .A3(new_n921), .ZN(G63));
  XNOR2_X1  g736(.A(new_n442), .B(KEYINPUT60), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n888), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n896), .B1(new_n925), .B2(new_n435), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n923), .B1(new_n829), .B2(new_n842), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n927), .A2(KEYINPUT123), .A3(new_n649), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT123), .B1(new_n927), .B2(new_n649), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n926), .B(KEYINPUT61), .C1(new_n928), .C2(new_n929), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(G66));
  OAI21_X1  g748(.A(G953), .B1(new_n588), .B2(new_n216), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n816), .A2(new_n781), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n937), .B2(G953), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n891), .B1(G898), .B2(new_n427), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G69));
  AND2_X1   g754(.A1(new_n772), .A2(new_n778), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n942));
  INV_X1    g756(.A(new_n688), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n819), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n795), .A2(KEYINPUT124), .A3(new_n688), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n767), .A2(new_n768), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n727), .A2(new_n681), .A3(new_n667), .ZN(new_n948));
  AOI22_X1  g762(.A1(new_n947), .A2(new_n948), .B1(new_n661), .B2(new_n728), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n941), .A2(new_n738), .A3(new_n946), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n427), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n346), .A2(new_n351), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(new_n494), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n659), .B2(G953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n683), .B1(new_n944), .B2(new_n945), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n946), .B1(new_n682), .B2(new_n680), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n962), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n665), .B1(new_n604), .B2(new_n800), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n965), .A2(new_n453), .A3(new_n769), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT126), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n772), .A2(new_n778), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n959), .B2(new_n960), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n954), .A2(new_n427), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n956), .B(new_n957), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n964), .B2(new_n969), .ZN(new_n973));
  INV_X1    g787(.A(new_n955), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n950), .B2(new_n427), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT127), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n427), .B1(G227), .B2(G900), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n972), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n972), .B2(new_n976), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(G72));
  INV_X1    g794(.A(new_n380), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n970), .A2(new_n937), .ZN(new_n982));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  AOI211_X1 g798(.A(new_n363), .B(new_n981), .C1(new_n982), .C2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n950), .B2(new_n936), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n363), .A3(new_n981), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n381), .A2(new_n366), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n984), .B(new_n988), .C1(new_n821), .C2(new_n822), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n989), .A3(new_n913), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n985), .A2(new_n990), .ZN(G57));
endmodule


