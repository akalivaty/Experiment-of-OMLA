

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U553 ( .A1(n534), .A2(n520), .ZN(G164) );
  XNOR2_X1 U554 ( .A(n734), .B(KEYINPUT101), .ZN(n767) );
  BUF_X1 U555 ( .A(n560), .Z(n530) );
  NOR2_X1 U556 ( .A1(n524), .A2(n523), .ZN(n903) );
  XNOR2_X1 U557 ( .A(KEYINPUT32), .B(KEYINPUT107), .ZN(n753) );
  NOR2_X2 U558 ( .A1(G2105), .A2(n531), .ZN(n906) );
  AND2_X1 U559 ( .A1(n533), .A2(n532), .ZN(n520) );
  OR2_X1 U560 ( .A1(n763), .A2(n770), .ZN(n521) );
  OR2_X1 U561 ( .A1(n787), .A2(n786), .ZN(n522) );
  INV_X1 U562 ( .A(G8), .ZN(n735) );
  NOR2_X1 U563 ( .A1(n741), .A2(n740), .ZN(n742) );
  OR2_X1 U564 ( .A1(n769), .A2(n776), .ZN(n773) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XNOR2_X1 U566 ( .A(n754), .B(n753), .ZN(n775) );
  OR2_X1 U567 ( .A1(n775), .A2(n774), .ZN(n785) );
  AND2_X1 U568 ( .A1(n690), .A2(G40), .ZN(n691) );
  NOR2_X1 U569 ( .A1(G164), .A2(G1384), .ZN(n810) );
  AND2_X1 U570 ( .A1(n821), .A2(n833), .ZN(n822) );
  NOR2_X1 U571 ( .A1(G651), .A2(n645), .ZN(n654) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n652) );
  XNOR2_X1 U573 ( .A(n527), .B(KEYINPUT93), .ZN(n534) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n902) );
  NAND2_X1 U575 ( .A1(n902), .A2(G114), .ZN(n526) );
  INV_X1 U576 ( .A(G2105), .ZN(n524) );
  XOR2_X1 U577 ( .A(G2104), .B(KEYINPUT65), .Z(n523) );
  NAND2_X1 U578 ( .A1(G126), .A2(n903), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U580 ( .A(n528), .B(KEYINPUT17), .ZN(n529) );
  XNOR2_X1 U581 ( .A(n529), .B(KEYINPUT67), .ZN(n560) );
  NAND2_X1 U582 ( .A1(n530), .A2(G138), .ZN(n533) );
  XNOR2_X1 U583 ( .A(KEYINPUT65), .B(G2104), .ZN(n531) );
  NAND2_X1 U584 ( .A1(G102), .A2(n906), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G89), .A2(n652), .ZN(n535) );
  XNOR2_X1 U586 ( .A(n535), .B(KEYINPUT78), .ZN(n536) );
  XNOR2_X1 U587 ( .A(n536), .B(KEYINPUT4), .ZN(n539) );
  INV_X1 U588 ( .A(G651), .ZN(n541) );
  XOR2_X1 U589 ( .A(KEYINPUT0), .B(G543), .Z(n645) );
  OR2_X1 U590 ( .A1(n541), .A2(n645), .ZN(n537) );
  XOR2_X1 U591 ( .A(KEYINPUT70), .B(n537), .Z(n659) );
  NAND2_X1 U592 ( .A1(G76), .A2(n659), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U594 ( .A(KEYINPUT5), .B(n540), .ZN(n549) );
  XNOR2_X1 U595 ( .A(KEYINPUT6), .B(KEYINPUT80), .ZN(n547) );
  NAND2_X1 U596 ( .A1(n654), .A2(G51), .ZN(n545) );
  NOR2_X1 U597 ( .A1(G543), .A2(n541), .ZN(n542) );
  XOR2_X1 U598 ( .A(KEYINPUT1), .B(n542), .Z(n653) );
  NAND2_X1 U599 ( .A1(n653), .A2(G63), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT79), .B(n543), .Z(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U602 ( .A(n547), .B(n546), .Z(n548) );
  NAND2_X1 U603 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U604 ( .A(KEYINPUT7), .B(n550), .ZN(G168) );
  XOR2_X1 U605 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U606 ( .A1(G77), .A2(n659), .ZN(n551) );
  XOR2_X1 U607 ( .A(KEYINPUT71), .B(n551), .Z(n553) );
  NAND2_X1 U608 ( .A1(n652), .A2(G90), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U610 ( .A(KEYINPUT72), .B(KEYINPUT9), .ZN(n554) );
  XNOR2_X1 U611 ( .A(n555), .B(n554), .ZN(n559) );
  NAND2_X1 U612 ( .A1(G64), .A2(n653), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G52), .A2(n654), .ZN(n556) );
  AND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(G301) );
  INV_X1 U616 ( .A(G301), .ZN(G171) );
  NAND2_X1 U617 ( .A1(n560), .A2(G137), .ZN(n561) );
  XNOR2_X1 U618 ( .A(n561), .B(KEYINPUT68), .ZN(n563) );
  NAND2_X1 U619 ( .A1(G113), .A2(n902), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U621 ( .A(n564), .B(KEYINPUT69), .ZN(n566) );
  NAND2_X1 U622 ( .A1(G125), .A2(n903), .ZN(n565) );
  AND2_X1 U623 ( .A1(n566), .A2(n565), .ZN(n690) );
  NAND2_X1 U624 ( .A1(n906), .A2(G101), .ZN(n567) );
  XNOR2_X1 U625 ( .A(n567), .B(KEYINPUT23), .ZN(n568) );
  XOR2_X1 U626 ( .A(n568), .B(KEYINPUT66), .Z(n692) );
  AND2_X1 U627 ( .A1(n690), .A2(n692), .ZN(G160) );
  AND2_X1 U628 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U629 ( .A1(G65), .A2(n653), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G53), .A2(n654), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G91), .A2(n652), .ZN(n572) );
  NAND2_X1 U633 ( .A1(G78), .A2(n659), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n993) );
  INV_X1 U636 ( .A(n993), .ZN(G299) );
  INV_X1 U637 ( .A(G57), .ZN(G237) );
  INV_X1 U638 ( .A(G82), .ZN(G220) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT10), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT74), .B(n576), .ZN(G223) );
  INV_X1 U642 ( .A(G223), .ZN(n840) );
  NAND2_X1 U643 ( .A1(n840), .A2(G567), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  NAND2_X1 U645 ( .A1(G56), .A2(n653), .ZN(n578) );
  XOR2_X1 U646 ( .A(KEYINPUT14), .B(n578), .Z(n585) );
  NAND2_X1 U647 ( .A1(G81), .A2(n652), .ZN(n579) );
  XOR2_X1 U648 ( .A(KEYINPUT12), .B(n579), .Z(n580) );
  XNOR2_X1 U649 ( .A(n580), .B(KEYINPUT75), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G68), .A2(n659), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U652 ( .A(KEYINPUT13), .B(n583), .Z(n584) );
  NOR2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n654), .A2(G43), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n982) );
  INV_X1 U656 ( .A(n982), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n588), .A2(G860), .ZN(G153) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U659 ( .A1(G66), .A2(n653), .ZN(n589) );
  XNOR2_X1 U660 ( .A(n589), .B(KEYINPUT76), .ZN(n596) );
  NAND2_X1 U661 ( .A1(G92), .A2(n652), .ZN(n591) );
  NAND2_X1 U662 ( .A1(G79), .A2(n659), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U664 ( .A1(G54), .A2(n654), .ZN(n592) );
  XNOR2_X1 U665 ( .A(KEYINPUT77), .B(n592), .ZN(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U668 ( .A(KEYINPUT15), .B(n597), .Z(n705) );
  INV_X1 U669 ( .A(n705), .ZN(n979) );
  OR2_X1 U670 ( .A1(n979), .A2(G868), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n599), .A2(n598), .ZN(G284) );
  XNOR2_X1 U672 ( .A(KEYINPUT81), .B(G868), .ZN(n600) );
  NOR2_X1 U673 ( .A1(G286), .A2(n600), .ZN(n601) );
  XNOR2_X1 U674 ( .A(n601), .B(KEYINPUT82), .ZN(n603) );
  NOR2_X1 U675 ( .A1(G299), .A2(G868), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n603), .A2(n602), .ZN(G297) );
  INV_X1 U677 ( .A(G559), .ZN(n604) );
  NOR2_X1 U678 ( .A1(G860), .A2(n604), .ZN(n605) );
  XNOR2_X1 U679 ( .A(KEYINPUT83), .B(n605), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n606), .A2(n979), .ZN(n607) );
  XNOR2_X1 U681 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U682 ( .A1(G868), .A2(n982), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G868), .A2(n979), .ZN(n608) );
  NOR2_X1 U684 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U685 ( .A1(n610), .A2(n609), .ZN(G282) );
  XOR2_X1 U686 ( .A(KEYINPUT84), .B(KEYINPUT18), .Z(n612) );
  NAND2_X1 U687 ( .A1(G123), .A2(n903), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n612), .B(n611), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G111), .A2(n902), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G99), .A2(n906), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U692 ( .A(KEYINPUT85), .B(n615), .Z(n616) );
  NOR2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n530), .A2(G135), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n941) );
  XOR2_X1 U696 ( .A(G2096), .B(KEYINPUT86), .Z(n620) );
  XNOR2_X1 U697 ( .A(n941), .B(n620), .ZN(n622) );
  INV_X1 U698 ( .A(G2100), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(G156) );
  NAND2_X1 U700 ( .A1(n979), .A2(G559), .ZN(n673) );
  XNOR2_X1 U701 ( .A(n982), .B(n673), .ZN(n623) );
  NOR2_X1 U702 ( .A1(n623), .A2(G860), .ZN(n630) );
  NAND2_X1 U703 ( .A1(G67), .A2(n653), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G55), .A2(n654), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G93), .A2(n652), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G80), .A2(n659), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n668) );
  XNOR2_X1 U710 ( .A(n630), .B(n668), .ZN(G145) );
  NAND2_X1 U711 ( .A1(G62), .A2(n653), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G50), .A2(n654), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U714 ( .A(KEYINPUT88), .B(n633), .ZN(n637) );
  NAND2_X1 U715 ( .A1(G88), .A2(n652), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G75), .A2(n659), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n637), .A2(n636), .ZN(G166) );
  NAND2_X1 U719 ( .A1(G86), .A2(n652), .ZN(n639) );
  NAND2_X1 U720 ( .A1(G48), .A2(n654), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n659), .A2(G73), .ZN(n640) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n640), .Z(n641) );
  NOR2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n653), .A2(G61), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G49), .A2(n654), .ZN(n647) );
  NAND2_X1 U728 ( .A1(G87), .A2(n645), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U730 ( .A1(n653), .A2(n648), .ZN(n651) );
  NAND2_X1 U731 ( .A1(G74), .A2(G651), .ZN(n649) );
  XOR2_X1 U732 ( .A(KEYINPUT87), .B(n649), .Z(n650) );
  NAND2_X1 U733 ( .A1(n651), .A2(n650), .ZN(G288) );
  AND2_X1 U734 ( .A1(n652), .A2(G85), .ZN(n658) );
  NAND2_X1 U735 ( .A1(G60), .A2(n653), .ZN(n656) );
  NAND2_X1 U736 ( .A1(G47), .A2(n654), .ZN(n655) );
  NAND2_X1 U737 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U738 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U739 ( .A1(G72), .A2(n659), .ZN(n660) );
  NAND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(G290) );
  INV_X1 U741 ( .A(G868), .ZN(n662) );
  NAND2_X1 U742 ( .A1(n668), .A2(n662), .ZN(n676) );
  XOR2_X1 U743 ( .A(KEYINPUT89), .B(KEYINPUT19), .Z(n664) );
  XNOR2_X1 U744 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n663) );
  XNOR2_X1 U745 ( .A(n664), .B(n663), .ZN(n667) );
  XNOR2_X1 U746 ( .A(G166), .B(n982), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n665), .B(G305), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n667), .B(n666), .ZN(n670) );
  XNOR2_X1 U749 ( .A(G288), .B(n668), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U751 ( .A(n671), .B(G290), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n672), .B(G299), .ZN(n917) );
  XOR2_X1 U753 ( .A(n917), .B(n673), .Z(n674) );
  NAND2_X1 U754 ( .A1(G868), .A2(n674), .ZN(n675) );
  NAND2_X1 U755 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U756 ( .A(KEYINPUT92), .B(n677), .Z(G295) );
  NAND2_X1 U757 ( .A1(G2084), .A2(G2078), .ZN(n678) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U761 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U763 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U766 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U767 ( .A1(G96), .A2(n684), .ZN(n845) );
  NAND2_X1 U768 ( .A1(n845), .A2(G2106), .ZN(n688) );
  NAND2_X1 U769 ( .A1(G69), .A2(G120), .ZN(n685) );
  NOR2_X1 U770 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U771 ( .A1(G108), .A2(n686), .ZN(n844) );
  NAND2_X1 U772 ( .A1(n844), .A2(G567), .ZN(n687) );
  NAND2_X1 U773 ( .A1(n688), .A2(n687), .ZN(n926) );
  NAND2_X1 U774 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U775 ( .A1(n926), .A2(n689), .ZN(n843) );
  NAND2_X1 U776 ( .A1(n843), .A2(G36), .ZN(G176) );
  XOR2_X1 U777 ( .A(KEYINPUT94), .B(G166), .Z(G303) );
  NAND2_X1 U778 ( .A1(n692), .A2(n691), .ZN(n809) );
  INV_X1 U779 ( .A(n809), .ZN(n693) );
  NAND2_X1 U780 ( .A1(n693), .A2(n810), .ZN(n694) );
  XNOR2_X1 U781 ( .A(n694), .B(KEYINPUT64), .ZN(n733) );
  INV_X1 U782 ( .A(n733), .ZN(n700) );
  NAND2_X1 U783 ( .A1(n700), .A2(G1996), .ZN(n697) );
  INV_X1 U784 ( .A(n697), .ZN(n696) );
  INV_X1 U785 ( .A(KEYINPUT26), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U787 ( .A1(n697), .A2(KEYINPUT26), .ZN(n698) );
  NAND2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n702) );
  INV_X1 U789 ( .A(n700), .ZN(n746) );
  NAND2_X1 U790 ( .A1(n746), .A2(G1341), .ZN(n701) );
  NAND2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n707) );
  NOR2_X1 U792 ( .A1(n982), .A2(n707), .ZN(n703) );
  NOR2_X1 U793 ( .A1(n979), .A2(n703), .ZN(n704) );
  XNOR2_X1 U794 ( .A(n704), .B(KEYINPUT103), .ZN(n714) );
  OR2_X1 U795 ( .A1(n705), .A2(n982), .ZN(n706) );
  OR2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U797 ( .A(KEYINPUT102), .B(n708), .ZN(n712) );
  NOR2_X1 U798 ( .A1(G2067), .A2(n746), .ZN(n710) );
  INV_X1 U799 ( .A(n746), .ZN(n717) );
  NOR2_X1 U800 ( .A1(G1348), .A2(n717), .ZN(n709) );
  NOR2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U804 ( .A(n715), .B(KEYINPUT104), .ZN(n721) );
  NAND2_X1 U805 ( .A1(G2072), .A2(n717), .ZN(n716) );
  XNOR2_X1 U806 ( .A(n716), .B(KEYINPUT27), .ZN(n719) );
  INV_X1 U807 ( .A(G1956), .ZN(n1005) );
  NOR2_X1 U808 ( .A1(n717), .A2(n1005), .ZN(n718) );
  NOR2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U810 ( .A1(n722), .A2(n993), .ZN(n720) );
  NAND2_X1 U811 ( .A1(n721), .A2(n720), .ZN(n725) );
  NOR2_X1 U812 ( .A1(n722), .A2(n993), .ZN(n723) );
  XOR2_X1 U813 ( .A(n723), .B(KEYINPUT28), .Z(n724) );
  NAND2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n727) );
  XNOR2_X1 U815 ( .A(KEYINPUT29), .B(KEYINPUT105), .ZN(n726) );
  XNOR2_X1 U816 ( .A(n727), .B(n726), .ZN(n731) );
  AND2_X1 U817 ( .A1(n746), .A2(G1961), .ZN(n729) );
  XNOR2_X1 U818 ( .A(KEYINPUT25), .B(G2078), .ZN(n957) );
  NOR2_X1 U819 ( .A1(n746), .A2(n957), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n732), .A2(G171), .ZN(n730) );
  NAND2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n745) );
  NOR2_X1 U823 ( .A1(G171), .A2(n732), .ZN(n741) );
  AND2_X1 U824 ( .A1(n733), .A2(G8), .ZN(n734) );
  NOR2_X1 U825 ( .A1(G1966), .A2(n767), .ZN(n758) );
  INV_X1 U826 ( .A(n758), .ZN(n737) );
  NOR2_X1 U827 ( .A1(n746), .A2(G2084), .ZN(n755) );
  NOR2_X1 U828 ( .A1(n755), .A2(n735), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U830 ( .A(KEYINPUT30), .B(n738), .ZN(n739) );
  NOR2_X1 U831 ( .A1(n739), .A2(G168), .ZN(n740) );
  XOR2_X1 U832 ( .A(n742), .B(KEYINPUT106), .Z(n743) );
  XNOR2_X1 U833 ( .A(n743), .B(KEYINPUT31), .ZN(n744) );
  NAND2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n757) );
  NAND2_X1 U835 ( .A1(n757), .A2(G286), .ZN(n751) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n767), .ZN(n748) );
  NOR2_X1 U837 ( .A1(n746), .A2(G2090), .ZN(n747) );
  NOR2_X1 U838 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n749), .A2(G303), .ZN(n750) );
  NAND2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U841 ( .A1(n752), .A2(G8), .ZN(n754) );
  NAND2_X1 U842 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U843 ( .A1(n757), .A2(n756), .ZN(n759) );
  NOR2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n769) );
  NOR2_X1 U845 ( .A1(n775), .A2(n769), .ZN(n762) );
  INV_X1 U846 ( .A(G2090), .ZN(n956) );
  NAND2_X1 U847 ( .A1(G8), .A2(n956), .ZN(n760) );
  NOR2_X1 U848 ( .A1(n760), .A2(G303), .ZN(n761) );
  NOR2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n763) );
  INV_X1 U850 ( .A(n767), .ZN(n770) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XNOR2_X1 U852 ( .A(n764), .B(KEYINPUT24), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n765), .A2(n770), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n521), .A2(n766), .ZN(n787) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n996) );
  INV_X1 U856 ( .A(n996), .ZN(n768) );
  OR2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n776) );
  NOR2_X1 U858 ( .A1(G1976), .A2(G288), .ZN(n778) );
  AND2_X1 U859 ( .A1(n778), .A2(KEYINPUT33), .ZN(n771) );
  AND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U861 ( .A(G1981), .B(G305), .ZN(n988) );
  OR2_X1 U862 ( .A1(n772), .A2(n988), .ZN(n783) );
  OR2_X1 U863 ( .A1(n773), .A2(n783), .ZN(n774) );
  INV_X1 U864 ( .A(n776), .ZN(n780) );
  NOR2_X1 U865 ( .A1(G303), .A2(G1971), .ZN(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n997) );
  INV_X1 U867 ( .A(n997), .ZN(n779) );
  AND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U869 ( .A1(n781), .A2(KEYINPUT33), .ZN(n782) );
  OR2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U872 ( .A(G1986), .B(G290), .Z(n980) );
  NAND2_X1 U873 ( .A1(G105), .A2(n906), .ZN(n790) );
  XOR2_X1 U874 ( .A(KEYINPUT96), .B(KEYINPUT38), .Z(n788) );
  XNOR2_X1 U875 ( .A(KEYINPUT97), .B(n788), .ZN(n789) );
  XNOR2_X1 U876 ( .A(n790), .B(n789), .ZN(n797) );
  NAND2_X1 U877 ( .A1(n902), .A2(G117), .ZN(n792) );
  NAND2_X1 U878 ( .A1(G129), .A2(n903), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U880 ( .A1(n530), .A2(G141), .ZN(n793) );
  XOR2_X1 U881 ( .A(KEYINPUT98), .B(n793), .Z(n794) );
  NOR2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n892) );
  NAND2_X1 U884 ( .A1(G1996), .A2(n892), .ZN(n798) );
  XNOR2_X1 U885 ( .A(KEYINPUT99), .B(n798), .ZN(n807) );
  NAND2_X1 U886 ( .A1(n902), .A2(G107), .ZN(n800) );
  NAND2_X1 U887 ( .A1(G119), .A2(n903), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U889 ( .A1(n530), .A2(G131), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G95), .A2(n906), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  OR2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n895) );
  NAND2_X1 U893 ( .A1(G1991), .A2(n895), .ZN(n805) );
  XNOR2_X1 U894 ( .A(KEYINPUT95), .B(n805), .ZN(n806) );
  NOR2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U896 ( .A(n808), .B(KEYINPUT100), .ZN(n825) );
  NAND2_X1 U897 ( .A1(n980), .A2(n825), .ZN(n811) );
  NOR2_X1 U898 ( .A1(n810), .A2(n809), .ZN(n835) );
  NAND2_X1 U899 ( .A1(n811), .A2(n835), .ZN(n821) );
  XNOR2_X1 U900 ( .A(G2067), .B(KEYINPUT37), .ZN(n823) );
  NAND2_X1 U901 ( .A1(n902), .A2(G116), .ZN(n813) );
  NAND2_X1 U902 ( .A1(G128), .A2(n903), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U904 ( .A(n814), .B(KEYINPUT35), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n530), .A2(G140), .ZN(n816) );
  NAND2_X1 U906 ( .A1(G104), .A2(n906), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U908 ( .A(KEYINPUT34), .B(n817), .Z(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U910 ( .A(n820), .B(KEYINPUT36), .Z(n896) );
  NOR2_X1 U911 ( .A1(n823), .A2(n896), .ZN(n932) );
  NAND2_X1 U912 ( .A1(n835), .A2(n932), .ZN(n833) );
  NAND2_X1 U913 ( .A1(n522), .A2(n822), .ZN(n838) );
  AND2_X1 U914 ( .A1(n823), .A2(n896), .ZN(n824) );
  XOR2_X1 U915 ( .A(KEYINPUT110), .B(n824), .Z(n934) );
  XNOR2_X1 U916 ( .A(KEYINPUT109), .B(KEYINPUT39), .ZN(n831) );
  INV_X1 U917 ( .A(n825), .ZN(n949) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n826) );
  NOR2_X1 U919 ( .A1(G1991), .A2(n895), .ZN(n944) );
  NOR2_X1 U920 ( .A1(n826), .A2(n944), .ZN(n827) );
  NOR2_X1 U921 ( .A1(n949), .A2(n827), .ZN(n829) );
  NOR2_X1 U922 ( .A1(n892), .A2(G1996), .ZN(n828) );
  XNOR2_X1 U923 ( .A(n828), .B(KEYINPUT108), .ZN(n936) );
  NOR2_X1 U924 ( .A1(n829), .A2(n936), .ZN(n830) );
  XOR2_X1 U925 ( .A(n831), .B(n830), .Z(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n934), .A2(n834), .ZN(n836) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U929 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U930 ( .A(n839), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U933 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U935 ( .A1(n843), .A2(n842), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U941 ( .A(n846), .B(KEYINPUT112), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U943 ( .A(G1341), .B(G2454), .ZN(n847) );
  XNOR2_X1 U944 ( .A(n847), .B(G2430), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n848), .B(G1348), .ZN(n854) );
  XOR2_X1 U946 ( .A(G2443), .B(G2427), .Z(n850) );
  XNOR2_X1 U947 ( .A(G2438), .B(G2446), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U949 ( .A(G2451), .B(G2435), .Z(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n855) );
  NAND2_X1 U952 ( .A1(n855), .A2(G14), .ZN(n856) );
  XNOR2_X1 U953 ( .A(KEYINPUT111), .B(n856), .ZN(G401) );
  XOR2_X1 U954 ( .A(G2100), .B(G2096), .Z(n858) );
  XNOR2_X1 U955 ( .A(KEYINPUT42), .B(G2678), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U957 ( .A(KEYINPUT43), .B(G2090), .Z(n860) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U960 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U961 ( .A(G2084), .B(G2078), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(G227) );
  XOR2_X1 U963 ( .A(G1976), .B(G1981), .Z(n866) );
  XNOR2_X1 U964 ( .A(G1986), .B(G1966), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U966 ( .A(G1971), .B(G1956), .Z(n868) );
  XNOR2_X1 U967 ( .A(G1996), .B(G1991), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U969 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U970 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(G2474), .B(n873), .ZN(n874) );
  XOR2_X1 U973 ( .A(n874), .B(G1961), .Z(G229) );
  NAND2_X1 U974 ( .A1(n903), .A2(G124), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n875), .B(KEYINPUT44), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n876), .B(KEYINPUT114), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G112), .A2(n902), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n882) );
  NAND2_X1 U979 ( .A1(n530), .A2(G136), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G100), .A2(n906), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U983 ( .A(KEYINPUT115), .B(n883), .Z(G162) );
  NAND2_X1 U984 ( .A1(n530), .A2(G139), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G103), .A2(n906), .ZN(n884) );
  NAND2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n890) );
  NAND2_X1 U987 ( .A1(n902), .A2(G115), .ZN(n887) );
  NAND2_X1 U988 ( .A1(G127), .A2(n903), .ZN(n886) );
  NAND2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U990 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U992 ( .A(KEYINPUT116), .B(n891), .Z(n927) );
  XNOR2_X1 U993 ( .A(n892), .B(n927), .ZN(n894) );
  XNOR2_X1 U994 ( .A(G164), .B(G160), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n899) );
  XOR2_X1 U996 ( .A(n896), .B(n895), .Z(n897) );
  XNOR2_X1 U997 ( .A(n897), .B(n941), .ZN(n898) );
  XOR2_X1 U998 ( .A(n899), .B(n898), .Z(n901) );
  XNOR2_X1 U999 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n914) );
  NAND2_X1 U1001 ( .A1(n902), .A2(G118), .ZN(n905) );
  NAND2_X1 U1002 ( .A1(G130), .A2(n903), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(n911) );
  NAND2_X1 U1004 ( .A1(n530), .A2(G142), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(G106), .A2(n906), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1007 ( .A(KEYINPUT45), .B(n909), .Z(n910) );
  NOR2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(G162), .B(n912), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n915), .ZN(n916) );
  XOR2_X1 U1012 ( .A(KEYINPUT117), .B(n916), .Z(G395) );
  XOR2_X1 U1013 ( .A(n917), .B(G286), .Z(n919) );
  XNOR2_X1 U1014 ( .A(G171), .B(n979), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n920), .ZN(G397) );
  OR2_X1 U1017 ( .A1(n926), .A2(G401), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(G227), .A2(G229), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(n926), .ZN(G319) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n929) );
  XNOR2_X1 U1027 ( .A(G2072), .B(n927), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(n930), .B(KEYINPUT50), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(n931), .B(KEYINPUT121), .ZN(n952) );
  INV_X1 U1031 ( .A(n932), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n940) );
  XOR2_X1 U1033 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1035 ( .A(KEYINPUT51), .B(n937), .Z(n938) );
  XNOR2_X1 U1036 ( .A(n938), .B(KEYINPUT119), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(G160), .B(G2084), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(n945), .B(KEYINPUT118), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1044 ( .A(KEYINPUT120), .B(n950), .Z(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT52), .B(n953), .ZN(n954) );
  INV_X1 U1047 ( .A(KEYINPUT55), .ZN(n975) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n975), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n955), .A2(G29), .ZN(n1034) );
  XNOR2_X1 U1050 ( .A(G35), .B(n956), .ZN(n973) );
  XOR2_X1 U1051 ( .A(G27), .B(n957), .Z(n966) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(G33), .B(G2072), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n964) );
  XOR2_X1 U1055 ( .A(G1991), .B(G25), .Z(n960) );
  NAND2_X1 U1056 ( .A1(n960), .A2(G28), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G32), .B(G1996), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT122), .B(KEYINPUT53), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n968), .B(n967), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G2084), .B(G34), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(KEYINPUT54), .B(n969), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n975), .B(n974), .ZN(n977) );
  INV_X1 U1068 ( .A(G29), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(G11), .A2(n978), .ZN(n1032) );
  XNOR2_X1 U1071 ( .A(G16), .B(KEYINPUT56), .ZN(n1004) );
  XNOR2_X1 U1072 ( .A(G171), .B(G1961), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(G1348), .B(n979), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G1341), .B(n982), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n992) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G168), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(n987), .B(KEYINPUT123), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(KEYINPUT57), .B(n990), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n1002) );
  XNOR2_X1 U1083 ( .A(n993), .B(G1956), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(G1971), .A2(G303), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n999) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(KEYINPUT124), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1030) );
  INV_X1 U1091 ( .A(G16), .ZN(n1028) );
  XOR2_X1 U1092 ( .A(G5), .B(G1961), .Z(n1025) );
  XNOR2_X1 U1093 ( .A(G20), .B(n1005), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G1341), .B(G19), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G6), .B(G1981), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XOR2_X1 U1098 ( .A(KEYINPUT59), .B(G1348), .Z(n1010) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(KEYINPUT60), .B(n1013), .Z(n1015) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G21), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(KEYINPUT125), .B(n1016), .ZN(n1023) );
  XNOR2_X1 U1105 ( .A(G1971), .B(G22), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(G23), .B(G1976), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(G1986), .B(G24), .Z(n1019) );
  NAND2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1110 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1026), .Z(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1035), .Z(G311) );
  XOR2_X1 U1119 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

