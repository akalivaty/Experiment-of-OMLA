

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578;

  XNOR2_X1 U321 ( .A(n403), .B(n402), .ZN(n519) );
  XNOR2_X1 U322 ( .A(n401), .B(KEYINPUT48), .ZN(n402) );
  AND2_X1 U323 ( .A1(G232GAT), .A2(G233GAT), .ZN(n289) );
  INV_X1 U324 ( .A(KEYINPUT110), .ZN(n401) );
  XNOR2_X1 U325 ( .A(n343), .B(n289), .ZN(n344) );
  XNOR2_X1 U326 ( .A(n415), .B(n344), .ZN(n345) );
  XNOR2_X1 U327 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U328 ( .A(n356), .B(n355), .ZN(n555) );
  XNOR2_X1 U329 ( .A(n443), .B(G176GAT), .ZN(n444) );
  XNOR2_X1 U330 ( .A(n445), .B(n444), .ZN(G1349GAT) );
  XOR2_X1 U331 ( .A(G176GAT), .B(G64GAT), .Z(n329) );
  XOR2_X1 U332 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n291) );
  XNOR2_X1 U333 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n290) );
  XNOR2_X1 U334 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U335 ( .A(n329), .B(n292), .Z(n294) );
  NAND2_X1 U336 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U338 ( .A(G204GAT), .B(KEYINPUT72), .Z(n296) );
  XNOR2_X1 U339 ( .A(G148GAT), .B(KEYINPUT71), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U341 ( .A(G78GAT), .B(n297), .Z(n420) );
  XNOR2_X1 U342 ( .A(n298), .B(n420), .ZN(n303) );
  XOR2_X1 U343 ( .A(G92GAT), .B(G106GAT), .Z(n300) );
  XNOR2_X1 U344 ( .A(G99GAT), .B(G85GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n352) );
  XNOR2_X1 U346 ( .A(G71GAT), .B(G57GAT), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n301), .B(KEYINPUT13), .ZN(n371) );
  XOR2_X1 U348 ( .A(n352), .B(n371), .Z(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n572) );
  XNOR2_X1 U350 ( .A(KEYINPUT41), .B(n572), .ZN(n547) );
  XOR2_X1 U351 ( .A(KEYINPUT102), .B(n547), .Z(n529) );
  XOR2_X1 U352 ( .A(G162GAT), .B(G85GAT), .Z(n305) );
  NAND2_X1 U353 ( .A1(G225GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n308) );
  XOR2_X1 U355 ( .A(KEYINPUT85), .B(KEYINPUT3), .Z(n307) );
  XNOR2_X1 U356 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n421) );
  XOR2_X1 U358 ( .A(n308), .B(n421), .Z(n318) );
  XOR2_X1 U359 ( .A(KEYINPUT79), .B(KEYINPUT0), .Z(n310) );
  XNOR2_X1 U360 ( .A(G134GAT), .B(KEYINPUT80), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U362 ( .A(n311), .B(G127GAT), .Z(n313) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(G120GAT), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n438) );
  XOR2_X1 U365 ( .A(G148GAT), .B(KEYINPUT5), .Z(n315) );
  XNOR2_X1 U366 ( .A(KEYINPUT87), .B(G155GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n438), .B(n316), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n326) );
  XOR2_X1 U370 ( .A(KEYINPUT4), .B(KEYINPUT89), .Z(n320) );
  XNOR2_X1 U371 ( .A(KEYINPUT88), .B(KEYINPUT6), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U373 ( .A(KEYINPUT1), .B(G57GAT), .Z(n322) );
  XNOR2_X1 U374 ( .A(G29GAT), .B(G1GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U376 ( .A(n324), .B(n323), .Z(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n506) );
  XOR2_X1 U378 ( .A(KEYINPUT84), .B(KEYINPUT21), .Z(n328) );
  XNOR2_X1 U379 ( .A(G197GAT), .B(G211GAT), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n418) );
  XOR2_X1 U381 ( .A(n418), .B(n329), .Z(n333) );
  XOR2_X1 U382 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n331) );
  XNOR2_X1 U383 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n426) );
  XOR2_X1 U385 ( .A(G8GAT), .B(G183GAT), .Z(n359) );
  XNOR2_X1 U386 ( .A(n426), .B(n359), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n340) );
  XOR2_X1 U388 ( .A(G36GAT), .B(G190GAT), .Z(n343) );
  XOR2_X1 U389 ( .A(KEYINPUT90), .B(G204GAT), .Z(n335) );
  XNOR2_X1 U390 ( .A(G92GAT), .B(G218GAT), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U392 ( .A(n343), .B(n336), .Z(n338) );
  NAND2_X1 U393 ( .A1(G226GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n485) );
  XOR2_X1 U396 ( .A(KEYINPUT73), .B(G218GAT), .Z(n342) );
  XNOR2_X1 U397 ( .A(G50GAT), .B(G162GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n415) );
  XNOR2_X1 U399 ( .A(n345), .B(KEYINPUT9), .ZN(n356) );
  XOR2_X1 U400 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n347) );
  XNOR2_X1 U401 ( .A(G43GAT), .B(G29GAT), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U403 ( .A(KEYINPUT68), .B(n348), .Z(n378) );
  XOR2_X1 U404 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n350) );
  XNOR2_X1 U405 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n378), .B(n351), .ZN(n354) );
  XOR2_X1 U408 ( .A(n352), .B(KEYINPUT74), .Z(n353) );
  XNOR2_X1 U409 ( .A(n555), .B(KEYINPUT75), .ZN(n561) );
  XNOR2_X1 U410 ( .A(n561), .B(KEYINPUT36), .ZN(n478) );
  XOR2_X1 U411 ( .A(G211GAT), .B(KEYINPUT76), .Z(n358) );
  XNOR2_X1 U412 ( .A(KEYINPUT77), .B(KEYINPUT12), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U414 ( .A(G22GAT), .B(G155GAT), .Z(n411) );
  XOR2_X1 U415 ( .A(G64GAT), .B(n411), .Z(n361) );
  XNOR2_X1 U416 ( .A(G127GAT), .B(n359), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U418 ( .A(n363), .B(n362), .Z(n365) );
  NAND2_X1 U419 ( .A1(G231GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U421 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n367) );
  XNOR2_X1 U422 ( .A(G78GAT), .B(KEYINPUT78), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U424 ( .A(n369), .B(n368), .Z(n373) );
  XNOR2_X1 U425 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n370), .B(G15GAT), .ZN(n379) );
  XNOR2_X1 U427 ( .A(n379), .B(n371), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n393) );
  NAND2_X1 U429 ( .A1(n478), .A2(n393), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n374), .B(KEYINPUT45), .ZN(n392) );
  XOR2_X1 U431 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n376) );
  XNOR2_X1 U432 ( .A(G22GAT), .B(KEYINPUT70), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n389) );
  XOR2_X1 U435 ( .A(G50GAT), .B(G36GAT), .Z(n381) );
  XNOR2_X1 U436 ( .A(G113GAT), .B(n379), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U438 ( .A(n382), .B(G141GAT), .Z(n387) );
  XOR2_X1 U439 ( .A(G197GAT), .B(G8GAT), .Z(n384) );
  NAND2_X1 U440 ( .A1(G229GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(G169GAT), .B(n385), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n567) );
  INV_X1 U445 ( .A(n567), .ZN(n545) );
  INV_X1 U446 ( .A(n572), .ZN(n390) );
  NAND2_X1 U447 ( .A1(n545), .A2(n390), .ZN(n391) );
  NOR2_X1 U448 ( .A1(n392), .A2(n391), .ZN(n400) );
  XOR2_X1 U449 ( .A(KEYINPUT47), .B(KEYINPUT109), .Z(n398) );
  XNOR2_X1 U450 ( .A(KEYINPUT108), .B(n393), .ZN(n559) );
  NOR2_X1 U451 ( .A1(n545), .A2(n547), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n394), .B(KEYINPUT46), .ZN(n395) );
  NOR2_X1 U453 ( .A1(n559), .A2(n395), .ZN(n396) );
  NAND2_X1 U454 ( .A1(n396), .A2(n555), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n399) );
  NOR2_X1 U456 ( .A1(n400), .A2(n399), .ZN(n403) );
  NAND2_X1 U457 ( .A1(n485), .A2(n519), .ZN(n405) );
  XOR2_X1 U458 ( .A(KEYINPUT124), .B(KEYINPUT54), .Z(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n406) );
  NAND2_X1 U460 ( .A1(n506), .A2(n406), .ZN(n407) );
  XNOR2_X1 U461 ( .A(n407), .B(KEYINPUT64), .ZN(n566) );
  XOR2_X1 U462 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n409) );
  XNOR2_X1 U463 ( .A(G106GAT), .B(KEYINPUT22), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U465 ( .A(n411), .B(n410), .Z(n413) );
  NAND2_X1 U466 ( .A1(G228GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U468 ( .A(n414), .B(KEYINPUT23), .Z(n417) );
  XNOR2_X1 U469 ( .A(n415), .B(KEYINPUT83), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U471 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U472 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U473 ( .A(n423), .B(n422), .ZN(n454) );
  NOR2_X1 U474 ( .A1(n566), .A2(n454), .ZN(n425) );
  XNOR2_X1 U475 ( .A(KEYINPUT125), .B(KEYINPUT55), .ZN(n424) );
  XNOR2_X1 U476 ( .A(n425), .B(n424), .ZN(n441) );
  XOR2_X1 U477 ( .A(G190GAT), .B(G99GAT), .Z(n428) );
  XNOR2_X1 U478 ( .A(G176GAT), .B(n426), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U480 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n430) );
  NAND2_X1 U481 ( .A1(G227GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U483 ( .A(n432), .B(n431), .Z(n434) );
  XNOR2_X1 U484 ( .A(G43GAT), .B(KEYINPUT65), .ZN(n433) );
  XNOR2_X1 U485 ( .A(n434), .B(n433), .ZN(n440) );
  XOR2_X1 U486 ( .A(KEYINPUT20), .B(G183GAT), .Z(n436) );
  XNOR2_X1 U487 ( .A(G15GAT), .B(G71GAT), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U489 ( .A(n438), .B(n437), .Z(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n521) );
  NAND2_X1 U491 ( .A1(n441), .A2(n521), .ZN(n442) );
  XOR2_X1 U492 ( .A(KEYINPUT126), .B(n442), .Z(n562) );
  NAND2_X1 U493 ( .A1(n529), .A2(n562), .ZN(n445) );
  XOR2_X1 U494 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n443) );
  XOR2_X1 U495 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n467) );
  NOR2_X1 U496 ( .A1(n572), .A2(n545), .ZN(n481) );
  XOR2_X1 U497 ( .A(KEYINPUT27), .B(n485), .Z(n451) );
  NOR2_X1 U498 ( .A1(n506), .A2(n451), .ZN(n518) );
  XOR2_X1 U499 ( .A(n454), .B(KEYINPUT67), .Z(n446) );
  XNOR2_X1 U500 ( .A(KEYINPUT28), .B(n446), .ZN(n523) );
  NOR2_X1 U501 ( .A1(n521), .A2(n523), .ZN(n447) );
  NAND2_X1 U502 ( .A1(n518), .A2(n447), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n448), .B(KEYINPUT91), .ZN(n460) );
  INV_X1 U504 ( .A(n506), .ZN(n465) );
  INV_X1 U505 ( .A(n521), .ZN(n511) );
  NAND2_X1 U506 ( .A1(n454), .A2(n511), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n449), .B(KEYINPUT26), .ZN(n450) );
  XNOR2_X1 U508 ( .A(KEYINPUT92), .B(n450), .ZN(n565) );
  NOR2_X1 U509 ( .A1(n451), .A2(n565), .ZN(n457) );
  NAND2_X1 U510 ( .A1(n521), .A2(n485), .ZN(n452) );
  XNOR2_X1 U511 ( .A(KEYINPUT93), .B(n452), .ZN(n453) );
  NOR2_X1 U512 ( .A1(n454), .A2(n453), .ZN(n455) );
  XOR2_X1 U513 ( .A(KEYINPUT25), .B(n455), .Z(n456) );
  NOR2_X1 U514 ( .A1(n457), .A2(n456), .ZN(n458) );
  NOR2_X1 U515 ( .A1(n465), .A2(n458), .ZN(n459) );
  NOR2_X1 U516 ( .A1(n460), .A2(n459), .ZN(n476) );
  INV_X1 U517 ( .A(n393), .ZN(n551) );
  NOR2_X1 U518 ( .A1(n551), .A2(n561), .ZN(n461) );
  XOR2_X1 U519 ( .A(KEYINPUT16), .B(n461), .Z(n462) );
  NOR2_X1 U520 ( .A1(n476), .A2(n462), .ZN(n463) );
  XNOR2_X1 U521 ( .A(KEYINPUT94), .B(n463), .ZN(n493) );
  NAND2_X1 U522 ( .A1(n481), .A2(n493), .ZN(n464) );
  XNOR2_X1 U523 ( .A(KEYINPUT95), .B(n464), .ZN(n473) );
  NAND2_X1 U524 ( .A1(n473), .A2(n465), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U526 ( .A(G1GAT), .B(n468), .Z(G1324GAT) );
  NAND2_X1 U527 ( .A1(n485), .A2(n473), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n469), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U529 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n471) );
  NAND2_X1 U530 ( .A1(n473), .A2(n521), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U532 ( .A(G15GAT), .B(n472), .Z(G1326GAT) );
  NAND2_X1 U533 ( .A1(n523), .A2(n473), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(KEYINPUT98), .ZN(n475) );
  XNOR2_X1 U535 ( .A(G22GAT), .B(n475), .ZN(G1327GAT) );
  NOR2_X1 U536 ( .A1(n393), .A2(n476), .ZN(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT99), .B(n477), .Z(n479) );
  NAND2_X1 U538 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n480), .B(KEYINPUT37), .ZN(n505) );
  NAND2_X1 U540 ( .A1(n481), .A2(n505), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT38), .ZN(n490) );
  NOR2_X1 U542 ( .A1(n490), .A2(n506), .ZN(n484) );
  XNOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1328GAT) );
  INV_X1 U545 ( .A(n485), .ZN(n509) );
  NOR2_X1 U546 ( .A1(n509), .A2(n490), .ZN(n486) );
  XOR2_X1 U547 ( .A(G36GAT), .B(n486), .Z(G1329GAT) );
  XNOR2_X1 U548 ( .A(KEYINPUT40), .B(KEYINPUT100), .ZN(n488) );
  NOR2_X1 U549 ( .A1(n511), .A2(n490), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U551 ( .A(G43GAT), .B(n489), .Z(G1330GAT) );
  XNOR2_X1 U552 ( .A(G50GAT), .B(KEYINPUT101), .ZN(n492) );
  INV_X1 U553 ( .A(n523), .ZN(n514) );
  NOR2_X1 U554 ( .A1(n514), .A2(n490), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(G1331GAT) );
  AND2_X1 U556 ( .A1(n545), .A2(n529), .ZN(n504) );
  NAND2_X1 U557 ( .A1(n504), .A2(n493), .ZN(n500) );
  NOR2_X1 U558 ( .A1(n506), .A2(n500), .ZN(n494) );
  XOR2_X1 U559 ( .A(G57GAT), .B(n494), .Z(n495) );
  XNOR2_X1 U560 ( .A(KEYINPUT42), .B(n495), .ZN(G1332GAT) );
  NOR2_X1 U561 ( .A1(n509), .A2(n500), .ZN(n497) );
  XNOR2_X1 U562 ( .A(G64GAT), .B(KEYINPUT103), .ZN(n496) );
  XNOR2_X1 U563 ( .A(n497), .B(n496), .ZN(G1333GAT) );
  NOR2_X1 U564 ( .A1(n511), .A2(n500), .ZN(n498) );
  XOR2_X1 U565 ( .A(KEYINPUT104), .B(n498), .Z(n499) );
  XNOR2_X1 U566 ( .A(G71GAT), .B(n499), .ZN(G1334GAT) );
  NOR2_X1 U567 ( .A1(n514), .A2(n500), .ZN(n502) );
  XNOR2_X1 U568 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U570 ( .A(G78GAT), .B(n503), .Z(G1335GAT) );
  NAND2_X1 U571 ( .A1(n505), .A2(n504), .ZN(n513) );
  NOR2_X1 U572 ( .A1(n506), .A2(n513), .ZN(n507) );
  XOR2_X1 U573 ( .A(KEYINPUT106), .B(n507), .Z(n508) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(n508), .ZN(G1336GAT) );
  NOR2_X1 U575 ( .A1(n509), .A2(n513), .ZN(n510) );
  XOR2_X1 U576 ( .A(G92GAT), .B(n510), .Z(G1337GAT) );
  NOR2_X1 U577 ( .A1(n511), .A2(n513), .ZN(n512) );
  XOR2_X1 U578 ( .A(G99GAT), .B(n512), .Z(G1338GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n516) );
  XNOR2_X1 U580 ( .A(KEYINPUT44), .B(KEYINPUT107), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(n517), .ZN(G1339GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(KEYINPUT111), .ZN(n544) );
  NAND2_X1 U585 ( .A1(n544), .A2(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(KEYINPUT112), .B(n522), .ZN(n524) );
  NOR2_X1 U587 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U588 ( .A(n525), .B(KEYINPUT113), .Z(n538) );
  AND2_X1 U589 ( .A1(n567), .A2(n538), .ZN(n527) );
  XNOR2_X1 U590 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT116), .Z(n531) );
  NAND2_X1 U594 ( .A1(n538), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U596 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(KEYINPUT119), .ZN(n537) );
  XOR2_X1 U599 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n535) );
  NAND2_X1 U600 ( .A1(n538), .A2(n559), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U604 ( .A1(n538), .A2(n561), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n542) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT120), .Z(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  INV_X1 U608 ( .A(n565), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n554) );
  NOR2_X1 U610 ( .A1(n545), .A2(n554), .ZN(n546) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  NOR2_X1 U612 ( .A1(n547), .A2(n554), .ZN(n549) );
  XNOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n551), .A2(n554), .ZN(n552) );
  XOR2_X1 U617 ( .A(KEYINPUT122), .B(n552), .Z(n553) );
  XNOR2_X1 U618 ( .A(G155GAT), .B(n553), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(KEYINPUT123), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n562), .A2(n567), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n562), .A2(n559), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n563), .B(KEYINPUT58), .ZN(n564) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(n564), .ZN(G1351GAT) );
  XOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT59), .Z(n569) );
  NOR2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n576) );
  NAND2_X1 U631 ( .A1(n576), .A2(n567), .ZN(n568) );
  XNOR2_X1 U632 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n570) );
  XNOR2_X1 U634 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U636 ( .A1(n576), .A2(n572), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n576), .A2(n393), .ZN(n575) );
  XNOR2_X1 U639 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n478), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT62), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

