

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U566 ( .A(n902), .Z(n532) );
  XNOR2_X1 U567 ( .A(KEYINPUT64), .B(n538), .ZN(n902) );
  NAND2_X1 U568 ( .A1(n796), .A2(n701), .ZN(n740) );
  AND2_X1 U569 ( .A1(n774), .A2(n773), .ZN(n782) );
  NAND2_X1 U570 ( .A1(n828), .A2(n825), .ZN(n533) );
  XOR2_X1 U571 ( .A(n725), .B(KEYINPUT29), .Z(n534) );
  OR2_X1 U572 ( .A1(G301), .A2(n736), .ZN(n535) );
  OR2_X1 U573 ( .A1(n795), .A2(n794), .ZN(n536) );
  XNOR2_X1 U574 ( .A(n731), .B(KEYINPUT98), .ZN(n784) );
  OR2_X1 U575 ( .A1(n788), .A2(n762), .ZN(n774) );
  OR2_X1 U576 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U577 ( .A(n698), .B(KEYINPUT86), .ZN(n797) );
  NOR2_X1 U578 ( .A1(n782), .A2(n781), .ZN(n795) );
  NOR2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n537) );
  NOR2_X1 U580 ( .A1(n826), .A2(n533), .ZN(n827) );
  NOR2_X1 U581 ( .A1(G651), .A2(n653), .ZN(n662) );
  XNOR2_X1 U582 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  AND2_X1 U583 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U584 ( .A(G132), .ZN(G219) );
  INV_X1 U585 ( .A(G57), .ZN(G237) );
  XOR2_X1 U586 ( .A(KEYINPUT17), .B(n537), .Z(n538) );
  NAND2_X1 U587 ( .A1(G137), .A2(n902), .ZN(n541) );
  INV_X1 U588 ( .A(G2105), .ZN(n542) );
  AND2_X1 U589 ( .A1(n542), .A2(G2104), .ZN(n900) );
  NAND2_X1 U590 ( .A1(G101), .A2(n900), .ZN(n539) );
  XOR2_X1 U591 ( .A(KEYINPUT23), .B(n539), .Z(n540) );
  NAND2_X1 U592 ( .A1(n541), .A2(n540), .ZN(n697) );
  NOR2_X1 U593 ( .A1(G2104), .A2(n542), .ZN(n897) );
  NAND2_X1 U594 ( .A1(G125), .A2(n897), .ZN(n544) );
  AND2_X1 U595 ( .A1(G2104), .A2(G2105), .ZN(n898) );
  NAND2_X1 U596 ( .A1(G113), .A2(n898), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n694) );
  NOR2_X1 U598 ( .A1(n697), .A2(n694), .ZN(G160) );
  INV_X1 U599 ( .A(KEYINPUT85), .ZN(n552) );
  NAND2_X1 U600 ( .A1(G126), .A2(n897), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G138), .A2(n902), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G102), .A2(n900), .ZN(n548) );
  NAND2_X1 U604 ( .A1(G114), .A2(n898), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U607 ( .A(n552), .B(n551), .ZN(G164) );
  NOR2_X1 U608 ( .A1(G543), .A2(G651), .ZN(n656) );
  NAND2_X1 U609 ( .A1(G89), .A2(n656), .ZN(n553) );
  XOR2_X1 U610 ( .A(KEYINPUT4), .B(n553), .Z(n554) );
  XNOR2_X1 U611 ( .A(n554), .B(KEYINPUT73), .ZN(n556) );
  XOR2_X1 U612 ( .A(G543), .B(KEYINPUT0), .Z(n653) );
  INV_X1 U613 ( .A(G651), .ZN(n558) );
  NOR2_X1 U614 ( .A1(n653), .A2(n558), .ZN(n657) );
  NAND2_X1 U615 ( .A1(G76), .A2(n657), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U617 ( .A(n557), .B(KEYINPUT5), .ZN(n565) );
  NAND2_X1 U618 ( .A1(G51), .A2(n662), .ZN(n562) );
  NOR2_X1 U619 ( .A1(G543), .A2(n558), .ZN(n559) );
  XOR2_X1 U620 ( .A(KEYINPUT66), .B(n559), .Z(n560) );
  XNOR2_X1 U621 ( .A(KEYINPUT1), .B(n560), .ZN(n661) );
  NAND2_X1 U622 ( .A1(G63), .A2(n661), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n563), .Z(n564) );
  NAND2_X1 U625 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n566), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U629 ( .A(n567), .B(KEYINPUT10), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT70), .B(n568), .Z(n941) );
  NAND2_X1 U631 ( .A1(n941), .A2(G567), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U633 ( .A1(G56), .A2(n661), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT14), .B(n570), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n656), .A2(G81), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G68), .A2(n657), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT13), .B(n574), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT71), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n662), .A2(G43), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n1044) );
  INV_X1 U644 ( .A(G860), .ZN(n631) );
  OR2_X1 U645 ( .A1(n1044), .A2(n631), .ZN(G153) );
  NAND2_X1 U646 ( .A1(G52), .A2(n662), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(KEYINPUT67), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G90), .A2(n656), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G77), .A2(n657), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U651 ( .A(KEYINPUT9), .B(n583), .Z(n584) );
  NOR2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G64), .A2(n661), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(G301) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n597) );
  NAND2_X1 U656 ( .A1(G66), .A2(n661), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G92), .A2(n656), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G79), .A2(n657), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U660 ( .A1(n662), .A2(G54), .ZN(n590) );
  XOR2_X1 U661 ( .A(KEYINPUT72), .B(n590), .Z(n591) );
  NOR2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U664 ( .A(KEYINPUT15), .B(n595), .ZN(n1028) );
  OR2_X1 U665 ( .A1(n1028), .A2(G868), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(G284) );
  NAND2_X1 U667 ( .A1(G53), .A2(n662), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G65), .A2(n661), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U670 ( .A(KEYINPUT68), .B(n600), .Z(n604) );
  NAND2_X1 U671 ( .A1(G91), .A2(n656), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G78), .A2(n657), .ZN(n601) );
  AND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(G299) );
  INV_X1 U675 ( .A(G868), .ZN(n675) );
  NOR2_X1 U676 ( .A1(G286), .A2(n675), .ZN(n606) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U678 ( .A1(n606), .A2(n605), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n631), .A2(G559), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n607), .A2(n1028), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n608), .B(KEYINPUT16), .ZN(n609) );
  XNOR2_X1 U682 ( .A(KEYINPUT74), .B(n609), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G559), .A2(n675), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n1028), .A2(n610), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n611), .B(KEYINPUT75), .ZN(n613) );
  NOR2_X1 U686 ( .A1(n1044), .A2(G868), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G123), .A2(n897), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n614), .B(KEYINPUT18), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n615), .B(KEYINPUT76), .ZN(n617) );
  NAND2_X1 U691 ( .A1(G99), .A2(n900), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n898), .A2(G111), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G135), .A2(n532), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n1002) );
  XNOR2_X1 U697 ( .A(n1002), .B(G2096), .ZN(n622) );
  INV_X1 U698 ( .A(G2100), .ZN(n852) );
  NAND2_X1 U699 ( .A1(n622), .A2(n852), .ZN(G156) );
  NAND2_X1 U700 ( .A1(G93), .A2(n656), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G80), .A2(n657), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U703 ( .A(KEYINPUT78), .B(n625), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G55), .A2(n662), .ZN(n627) );
  NAND2_X1 U705 ( .A1(G67), .A2(n661), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n628) );
  OR2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n674) );
  NAND2_X1 U708 ( .A1(G559), .A2(n1028), .ZN(n630) );
  XOR2_X1 U709 ( .A(n1044), .B(n630), .Z(n672) );
  NAND2_X1 U710 ( .A1(n631), .A2(n672), .ZN(n632) );
  XNOR2_X1 U711 ( .A(n632), .B(KEYINPUT77), .ZN(n633) );
  XOR2_X1 U712 ( .A(n674), .B(n633), .Z(G145) );
  NAND2_X1 U713 ( .A1(G73), .A2(n657), .ZN(n634) );
  XNOR2_X1 U714 ( .A(n634), .B(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U715 ( .A1(G86), .A2(n656), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G48), .A2(n662), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n661), .A2(G61), .ZN(n637) );
  XOR2_X1 U719 ( .A(KEYINPUT80), .B(n637), .Z(n638) );
  NOR2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U721 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G50), .A2(n662), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G62), .A2(n661), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U725 ( .A(KEYINPUT81), .B(n644), .ZN(n648) );
  NAND2_X1 U726 ( .A1(G88), .A2(n656), .ZN(n646) );
  NAND2_X1 U727 ( .A1(G75), .A2(n657), .ZN(n645) );
  AND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(G303) );
  NAND2_X1 U730 ( .A1(G49), .A2(n662), .ZN(n650) );
  NAND2_X1 U731 ( .A1(G74), .A2(G651), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U733 ( .A1(n661), .A2(n651), .ZN(n652) );
  XOR2_X1 U734 ( .A(KEYINPUT79), .B(n652), .Z(n655) );
  NAND2_X1 U735 ( .A1(n653), .A2(G87), .ZN(n654) );
  NAND2_X1 U736 ( .A1(n655), .A2(n654), .ZN(G288) );
  NAND2_X1 U737 ( .A1(G85), .A2(n656), .ZN(n659) );
  NAND2_X1 U738 ( .A1(G72), .A2(n657), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U740 ( .A(KEYINPUT65), .B(n660), .ZN(n666) );
  NAND2_X1 U741 ( .A1(n661), .A2(G60), .ZN(n664) );
  NAND2_X1 U742 ( .A1(G47), .A2(n662), .ZN(n663) );
  AND2_X1 U743 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U744 ( .A1(n666), .A2(n665), .ZN(G290) );
  XNOR2_X1 U745 ( .A(KEYINPUT19), .B(G305), .ZN(n671) );
  XOR2_X1 U746 ( .A(G299), .B(G303), .Z(n667) );
  XNOR2_X1 U747 ( .A(n667), .B(G288), .ZN(n668) );
  XOR2_X1 U748 ( .A(n674), .B(n668), .Z(n669) );
  XNOR2_X1 U749 ( .A(n669), .B(G290), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n671), .B(n670), .ZN(n919) );
  XNOR2_X1 U751 ( .A(n672), .B(n919), .ZN(n673) );
  NAND2_X1 U752 ( .A1(n673), .A2(G868), .ZN(n677) );
  NAND2_X1 U753 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U759 ( .A1(n681), .A2(G2072), .ZN(n682) );
  XNOR2_X1 U760 ( .A(KEYINPUT82), .B(n682), .ZN(G158) );
  XNOR2_X1 U761 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NAND2_X1 U762 ( .A1(G69), .A2(G120), .ZN(n683) );
  NOR2_X1 U763 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U764 ( .A1(G108), .A2(n684), .ZN(n850) );
  NAND2_X1 U765 ( .A1(G567), .A2(n850), .ZN(n685) );
  XNOR2_X1 U766 ( .A(n685), .B(KEYINPUT83), .ZN(n690) );
  NOR2_X1 U767 ( .A1(G219), .A2(G220), .ZN(n686) );
  XNOR2_X1 U768 ( .A(KEYINPUT22), .B(n686), .ZN(n687) );
  NAND2_X1 U769 ( .A1(n687), .A2(G96), .ZN(n688) );
  OR2_X1 U770 ( .A1(G218), .A2(n688), .ZN(n851) );
  AND2_X1 U771 ( .A1(G2106), .A2(n851), .ZN(n689) );
  NOR2_X1 U772 ( .A1(n690), .A2(n689), .ZN(G319) );
  INV_X1 U773 ( .A(G319), .ZN(n693) );
  NAND2_X1 U774 ( .A1(G661), .A2(G483), .ZN(n691) );
  XNOR2_X1 U775 ( .A(KEYINPUT84), .B(n691), .ZN(n692) );
  NOR2_X1 U776 ( .A1(n693), .A2(n692), .ZN(n848) );
  NAND2_X1 U777 ( .A1(n848), .A2(G36), .ZN(G176) );
  INV_X1 U778 ( .A(G303), .ZN(G166) );
  NOR2_X1 U779 ( .A1(G164), .A2(G1384), .ZN(n796) );
  INV_X1 U780 ( .A(KEYINPUT90), .ZN(n699) );
  INV_X1 U781 ( .A(G40), .ZN(n695) );
  OR2_X1 U782 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U783 ( .A(n699), .B(n797), .ZN(n701) );
  AND2_X1 U784 ( .A1(n796), .A2(n701), .ZN(n727) );
  NAND2_X1 U785 ( .A1(G2067), .A2(n727), .ZN(n700) );
  XNOR2_X1 U786 ( .A(KEYINPUT95), .B(n700), .ZN(n704) );
  NAND2_X1 U787 ( .A1(G1348), .A2(n740), .ZN(n702) );
  XOR2_X1 U788 ( .A(KEYINPUT94), .B(n702), .Z(n703) );
  NOR2_X1 U789 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U790 ( .A(n705), .B(KEYINPUT96), .ZN(n711) );
  INV_X1 U791 ( .A(G1996), .ZN(n942) );
  NOR2_X1 U792 ( .A1(n740), .A2(n942), .ZN(n706) );
  XOR2_X1 U793 ( .A(n706), .B(KEYINPUT26), .Z(n709) );
  AND2_X1 U794 ( .A1(n740), .A2(G1341), .ZN(n707) );
  NOR2_X1 U795 ( .A1(n707), .A2(n1044), .ZN(n708) );
  AND2_X1 U796 ( .A1(n709), .A2(n708), .ZN(n712) );
  AND2_X1 U797 ( .A1(n1028), .A2(n712), .ZN(n710) );
  NOR2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n714) );
  NOR2_X1 U799 ( .A1(n1028), .A2(n712), .ZN(n713) );
  NOR2_X1 U800 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U801 ( .A(KEYINPUT97), .B(n715), .ZN(n720) );
  NAND2_X1 U802 ( .A1(n727), .A2(G2072), .ZN(n716) );
  XNOR2_X1 U803 ( .A(n716), .B(KEYINPUT27), .ZN(n718) );
  INV_X1 U804 ( .A(G1956), .ZN(n861) );
  NOR2_X1 U805 ( .A1(n861), .A2(n727), .ZN(n717) );
  NOR2_X1 U806 ( .A1(n718), .A2(n717), .ZN(n721) );
  INV_X1 U807 ( .A(G299), .ZN(n1027) );
  NAND2_X1 U808 ( .A1(n721), .A2(n1027), .ZN(n719) );
  NAND2_X1 U809 ( .A1(n720), .A2(n719), .ZN(n724) );
  NOR2_X1 U810 ( .A1(n721), .A2(n1027), .ZN(n722) );
  XOR2_X1 U811 ( .A(n722), .B(KEYINPUT28), .Z(n723) );
  NAND2_X1 U812 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U813 ( .A(KEYINPUT25), .B(G2078), .Z(n943) );
  NOR2_X1 U814 ( .A1(n943), .A2(n740), .ZN(n726) );
  XOR2_X1 U815 ( .A(KEYINPUT93), .B(n726), .Z(n730) );
  NOR2_X1 U816 ( .A1(n727), .A2(G1961), .ZN(n728) );
  XNOR2_X1 U817 ( .A(KEYINPUT92), .B(n728), .ZN(n729) );
  NOR2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n736) );
  NAND2_X1 U819 ( .A1(n534), .A2(n535), .ZN(n731) );
  NAND2_X1 U820 ( .A1(G8), .A2(n740), .ZN(n732) );
  XNOR2_X1 U821 ( .A(KEYINPUT91), .B(n732), .ZN(n792) );
  INV_X1 U822 ( .A(n792), .ZN(n776) );
  NOR2_X1 U823 ( .A1(G1966), .A2(n776), .ZN(n757) );
  NOR2_X1 U824 ( .A1(G2084), .A2(n740), .ZN(n756) );
  NOR2_X1 U825 ( .A1(n757), .A2(n756), .ZN(n733) );
  NAND2_X1 U826 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U827 ( .A(KEYINPUT30), .B(n734), .ZN(n735) );
  NOR2_X1 U828 ( .A1(G168), .A2(n735), .ZN(n738) );
  AND2_X1 U829 ( .A1(G301), .A2(n736), .ZN(n737) );
  NOR2_X1 U830 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U831 ( .A(KEYINPUT31), .B(n739), .Z(n783) );
  INV_X1 U832 ( .A(G8), .ZN(n746) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n740), .ZN(n741) );
  XNOR2_X1 U834 ( .A(KEYINPUT99), .B(n741), .ZN(n744) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n776), .ZN(n742) );
  NOR2_X1 U836 ( .A1(G166), .A2(n742), .ZN(n743) );
  NAND2_X1 U837 ( .A1(n744), .A2(n743), .ZN(n745) );
  OR2_X1 U838 ( .A1(n746), .A2(n745), .ZN(n748) );
  AND2_X1 U839 ( .A1(n783), .A2(n748), .ZN(n747) );
  NAND2_X1 U840 ( .A1(n784), .A2(n747), .ZN(n752) );
  INV_X1 U841 ( .A(n748), .ZN(n750) );
  AND2_X1 U842 ( .A1(G286), .A2(G8), .ZN(n749) );
  OR2_X1 U843 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U844 ( .A1(n752), .A2(n751), .ZN(n754) );
  INV_X1 U845 ( .A(KEYINPUT32), .ZN(n753) );
  XNOR2_X1 U846 ( .A(n754), .B(n753), .ZN(n788) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n1024) );
  AND2_X1 U848 ( .A1(n783), .A2(n1024), .ZN(n755) );
  AND2_X1 U849 ( .A1(n784), .A2(n755), .ZN(n761) );
  NAND2_X1 U850 ( .A1(G8), .A2(n756), .ZN(n759) );
  INV_X1 U851 ( .A(n757), .ZN(n758) );
  NAND2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n785) );
  AND2_X1 U853 ( .A1(n1024), .A2(n785), .ZN(n760) );
  NOR2_X1 U854 ( .A1(n761), .A2(n760), .ZN(n762) );
  INV_X1 U855 ( .A(n1024), .ZN(n764) );
  NOR2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n765) );
  NOR2_X1 U857 ( .A1(G1971), .A2(G303), .ZN(n763) );
  NOR2_X1 U858 ( .A1(n765), .A2(n763), .ZN(n1036) );
  OR2_X1 U859 ( .A1(n764), .A2(n1036), .ZN(n769) );
  AND2_X1 U860 ( .A1(n765), .A2(KEYINPUT33), .ZN(n766) );
  AND2_X1 U861 ( .A1(n766), .A2(n792), .ZN(n767) );
  XNOR2_X1 U862 ( .A(G1981), .B(G305), .ZN(n1040) );
  OR2_X1 U863 ( .A1(n767), .A2(n1040), .ZN(n775) );
  INV_X1 U864 ( .A(n775), .ZN(n768) );
  NAND2_X1 U865 ( .A1(n768), .A2(KEYINPUT33), .ZN(n778) );
  AND2_X1 U866 ( .A1(n769), .A2(n778), .ZN(n772) );
  NOR2_X1 U867 ( .A1(G1981), .A2(G305), .ZN(n770) );
  XNOR2_X1 U868 ( .A(n770), .B(KEYINPUT24), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n771), .A2(n792), .ZN(n780) );
  AND2_X1 U870 ( .A1(n772), .A2(n780), .ZN(n773) );
  OR2_X1 U871 ( .A1(n776), .A2(n775), .ZN(n777) );
  AND2_X1 U872 ( .A1(n778), .A2(n777), .ZN(n779) );
  AND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n786) );
  NOR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G166), .A2(G8), .ZN(n789) );
  NOR2_X1 U878 ( .A1(G2090), .A2(n789), .ZN(n790) );
  NOR2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n793) );
  NOR2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U881 ( .A1(n797), .A2(n796), .ZN(n840) );
  NAND2_X1 U882 ( .A1(G140), .A2(n532), .ZN(n798) );
  XOR2_X1 U883 ( .A(KEYINPUT87), .B(n798), .Z(n800) );
  NAND2_X1 U884 ( .A1(n900), .A2(G104), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U886 ( .A(KEYINPUT34), .B(n801), .ZN(n807) );
  NAND2_X1 U887 ( .A1(G128), .A2(n897), .ZN(n803) );
  NAND2_X1 U888 ( .A1(G116), .A2(n898), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U890 ( .A(KEYINPUT88), .B(n804), .Z(n805) );
  XNOR2_X1 U891 ( .A(KEYINPUT35), .B(n805), .ZN(n806) );
  NOR2_X1 U892 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n808), .ZN(n884) );
  XNOR2_X1 U894 ( .A(G2067), .B(KEYINPUT37), .ZN(n837) );
  NOR2_X1 U895 ( .A1(n884), .A2(n837), .ZN(n1001) );
  NAND2_X1 U896 ( .A1(n840), .A2(n1001), .ZN(n835) );
  INV_X1 U897 ( .A(n835), .ZN(n826) );
  NAND2_X1 U898 ( .A1(G119), .A2(n897), .ZN(n810) );
  NAND2_X1 U899 ( .A1(G131), .A2(n532), .ZN(n809) );
  NAND2_X1 U900 ( .A1(n810), .A2(n809), .ZN(n814) );
  NAND2_X1 U901 ( .A1(G95), .A2(n900), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G107), .A2(n898), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n813) );
  OR2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n880) );
  NAND2_X1 U905 ( .A1(n880), .A2(G1991), .ZN(n823) );
  NAND2_X1 U906 ( .A1(G129), .A2(n897), .ZN(n816) );
  NAND2_X1 U907 ( .A1(G141), .A2(n532), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n819) );
  NAND2_X1 U909 ( .A1(n900), .A2(G105), .ZN(n817) );
  XOR2_X1 U910 ( .A(KEYINPUT38), .B(n817), .Z(n818) );
  NOR2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U912 ( .A1(n898), .A2(G117), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n913) );
  NAND2_X1 U914 ( .A1(G1996), .A2(n913), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U916 ( .A(n824), .B(KEYINPUT89), .Z(n997) );
  NAND2_X1 U917 ( .A1(n997), .A2(n840), .ZN(n828) );
  XNOR2_X1 U918 ( .A(G1986), .B(G290), .ZN(n1026) );
  NAND2_X1 U919 ( .A1(n840), .A2(n1026), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n536), .A2(n827), .ZN(n843) );
  NOR2_X1 U921 ( .A1(G1996), .A2(n913), .ZN(n1010) );
  INV_X1 U922 ( .A(n828), .ZN(n831) );
  NOR2_X1 U923 ( .A1(G1986), .A2(G290), .ZN(n829) );
  NOR2_X1 U924 ( .A1(G1991), .A2(n880), .ZN(n1003) );
  NOR2_X1 U925 ( .A1(n829), .A2(n1003), .ZN(n830) );
  NOR2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U927 ( .A(n832), .B(KEYINPUT100), .ZN(n833) );
  NOR2_X1 U928 ( .A1(n1010), .A2(n833), .ZN(n834) );
  XNOR2_X1 U929 ( .A(n834), .B(KEYINPUT39), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n836), .A2(n835), .ZN(n838) );
  NAND2_X1 U931 ( .A1(n884), .A2(n837), .ZN(n1012) );
  NAND2_X1 U932 ( .A1(n838), .A2(n1012), .ZN(n839) );
  NAND2_X1 U933 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U934 ( .A(KEYINPUT101), .B(n841), .Z(n842) );
  NAND2_X1 U935 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U936 ( .A(n844), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n941), .ZN(G217) );
  NAND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n845) );
  XNOR2_X1 U939 ( .A(KEYINPUT105), .B(n845), .ZN(n846) );
  NAND2_X1 U940 ( .A1(n846), .A2(G661), .ZN(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n847) );
  XNOR2_X1 U942 ( .A(KEYINPUT106), .B(n847), .ZN(n849) );
  NAND2_X1 U943 ( .A1(n849), .A2(n848), .ZN(G188) );
  INV_X1 U945 ( .A(G120), .ZN(G236) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  INV_X1 U947 ( .A(G69), .ZN(G235) );
  NOR2_X1 U948 ( .A1(n851), .A2(n850), .ZN(G325) );
  INV_X1 U949 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U950 ( .A(n852), .B(G2096), .ZN(n854) );
  XNOR2_X1 U951 ( .A(KEYINPUT42), .B(G2678), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U953 ( .A(KEYINPUT43), .B(G2090), .Z(n856) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U956 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U957 ( .A(G2078), .B(G2084), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(G227) );
  XNOR2_X1 U959 ( .A(G1981), .B(n861), .ZN(n863) );
  XNOR2_X1 U960 ( .A(G1991), .B(G1966), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U962 ( .A(G1986), .B(G1976), .Z(n865) );
  XNOR2_X1 U963 ( .A(G1961), .B(G1971), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U965 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U966 ( .A(G2474), .B(KEYINPUT107), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U968 ( .A(KEYINPUT41), .B(n870), .ZN(n871) );
  XOR2_X1 U969 ( .A(n871), .B(G1996), .Z(G229) );
  NAND2_X1 U970 ( .A1(n897), .A2(G124), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n872), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G136), .A2(n532), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U974 ( .A(KEYINPUT108), .B(n875), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G100), .A2(n900), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G112), .A2(n898), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U978 ( .A1(n879), .A2(n878), .ZN(G162) );
  XNOR2_X1 U979 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n882) );
  XNOR2_X1 U980 ( .A(n880), .B(G164), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U982 ( .A(KEYINPUT48), .B(n883), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n884), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n894) );
  NAND2_X1 U985 ( .A1(n900), .A2(G103), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G139), .A2(n532), .ZN(n887) );
  NAND2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G127), .A2(n897), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G115), .A2(n898), .ZN(n889) );
  NAND2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n992) );
  XOR2_X1 U993 ( .A(n894), .B(n992), .Z(n896) );
  XNOR2_X1 U994 ( .A(G160), .B(G162), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n915) );
  NAND2_X1 U996 ( .A1(G130), .A2(n897), .ZN(n910) );
  NAND2_X1 U997 ( .A1(n898), .A2(G118), .ZN(n899) );
  XNOR2_X1 U998 ( .A(KEYINPUT109), .B(n899), .ZN(n908) );
  NAND2_X1 U999 ( .A1(n900), .A2(G106), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n901), .B(KEYINPUT110), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(G142), .A2(n532), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(KEYINPUT45), .B(n905), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(KEYINPUT111), .B(n906), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n911), .B(n1002), .ZN(n912) );
  XOR2_X1 U1008 ( .A(n913), .B(n912), .Z(n914) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n916), .ZN(G395) );
  XOR2_X1 U1011 ( .A(KEYINPUT114), .B(G286), .Z(n918) );
  XOR2_X1 U1012 ( .A(G301), .B(n1028), .Z(n917) );
  XNOR2_X1 U1013 ( .A(n918), .B(n917), .ZN(n921) );
  XOR2_X1 U1014 ( .A(n1044), .B(n919), .Z(n920) );
  XNOR2_X1 U1015 ( .A(n921), .B(n920), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n922), .ZN(G397) );
  XOR2_X1 U1017 ( .A(G2435), .B(KEYINPUT104), .Z(n924) );
  XNOR2_X1 U1018 ( .A(G2454), .B(G2438), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(n924), .B(n923), .ZN(n928) );
  XOR2_X1 U1020 ( .A(G2446), .B(KEYINPUT103), .Z(n926) );
  XNOR2_X1 U1021 ( .A(G2451), .B(G2427), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(n926), .B(n925), .ZN(n927) );
  XOR2_X1 U1023 ( .A(n928), .B(n927), .Z(n930) );
  XNOR2_X1 U1024 ( .A(KEYINPUT102), .B(G2443), .ZN(n929) );
  XNOR2_X1 U1025 ( .A(n930), .B(n929), .ZN(n933) );
  XOR2_X1 U1026 ( .A(G1341), .B(G1348), .Z(n931) );
  XNOR2_X1 U1027 ( .A(G2430), .B(n931), .ZN(n932) );
  XOR2_X1 U1028 ( .A(n933), .B(n932), .Z(n934) );
  NAND2_X1 U1029 ( .A1(G14), .A2(n934), .ZN(n940) );
  NAND2_X1 U1030 ( .A1(G319), .A2(n940), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(G227), .A2(G229), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(KEYINPUT49), .B(n935), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(G395), .A2(G397), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(G225) );
  INV_X1 U1036 ( .A(G225), .ZN(G308) );
  INV_X1 U1037 ( .A(G108), .ZN(G238) );
  INV_X1 U1038 ( .A(n940), .ZN(G401) );
  INV_X1 U1039 ( .A(n941), .ZN(G223) );
  INV_X1 U1040 ( .A(G301), .ZN(G171) );
  XOR2_X1 U1041 ( .A(KEYINPUT123), .B(G29), .Z(n966) );
  XOR2_X1 U1042 ( .A(n942), .B(G32), .Z(n945) );
  XNOR2_X1 U1043 ( .A(n943), .B(G27), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(KEYINPUT120), .B(n946), .ZN(n952) );
  XOR2_X1 U1046 ( .A(G1991), .B(G25), .Z(n947) );
  NAND2_X1 U1047 ( .A1(n947), .A2(G28), .ZN(n950) );
  XOR2_X1 U1048 ( .A(KEYINPUT119), .B(G2067), .Z(n948) );
  XNOR2_X1 U1049 ( .A(G26), .B(n948), .ZN(n949) );
  NOR2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(n956), .B(KEYINPUT121), .ZN(n960) );
  XOR2_X1 U1056 ( .A(KEYINPUT122), .B(G34), .Z(n958) );
  XNOR2_X1 U1057 ( .A(G2084), .B(KEYINPUT54), .ZN(n957) );
  XNOR2_X1 U1058 ( .A(n958), .B(n957), .ZN(n959) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n963) );
  XNOR2_X1 U1060 ( .A(KEYINPUT118), .B(G2090), .ZN(n961) );
  XNOR2_X1 U1061 ( .A(G35), .B(n961), .ZN(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1063 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n1017) );
  XNOR2_X1 U1064 ( .A(n964), .B(n1017), .ZN(n965) );
  NOR2_X1 U1065 ( .A1(n966), .A2(n965), .ZN(n991) );
  XOR2_X1 U1066 ( .A(G20), .B(G1956), .Z(n970) );
  XNOR2_X1 U1067 ( .A(G1341), .B(G19), .ZN(n968) );
  XNOR2_X1 U1068 ( .A(G6), .B(G1981), .ZN(n967) );
  NOR2_X1 U1069 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1071 ( .A(KEYINPUT59), .B(G1348), .Z(n971) );
  XNOR2_X1 U1072 ( .A(G4), .B(n971), .ZN(n972) );
  NOR2_X1 U1073 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1074 ( .A(KEYINPUT60), .B(n974), .ZN(n978) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G21), .ZN(n976) );
  XNOR2_X1 U1076 ( .A(G1961), .B(G5), .ZN(n975) );
  NOR2_X1 U1077 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1078 ( .A1(n978), .A2(n977), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G1976), .B(G23), .ZN(n980) );
  XNOR2_X1 U1080 ( .A(G1986), .B(G24), .ZN(n979) );
  NOR2_X1 U1081 ( .A1(n980), .A2(n979), .ZN(n983) );
  XNOR2_X1 U1082 ( .A(G1971), .B(KEYINPUT127), .ZN(n981) );
  XNOR2_X1 U1083 ( .A(n981), .B(G22), .ZN(n982) );
  NAND2_X1 U1084 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1085 ( .A(KEYINPUT58), .B(n984), .ZN(n985) );
  NOR2_X1 U1086 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1087 ( .A(KEYINPUT61), .B(n987), .ZN(n988) );
  INV_X1 U1088 ( .A(G16), .ZN(n1022) );
  NAND2_X1 U1089 ( .A1(n988), .A2(n1022), .ZN(n989) );
  NAND2_X1 U1090 ( .A1(n989), .A2(G11), .ZN(n990) );
  NOR2_X1 U1091 ( .A1(n991), .A2(n990), .ZN(n1021) );
  XOR2_X1 U1092 ( .A(G2072), .B(n992), .Z(n994) );
  XOR2_X1 U1093 ( .A(G164), .B(G2078), .Z(n993) );
  NOR2_X1 U1094 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1095 ( .A(KEYINPUT116), .B(n995), .ZN(n996) );
  XNOR2_X1 U1096 ( .A(n996), .B(KEYINPUT50), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(G160), .B(G2084), .ZN(n999) );
  INV_X1 U1098 ( .A(n997), .ZN(n998) );
  NAND2_X1 U1099 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1100 ( .A1(n1001), .A2(n1000), .ZN(n1005) );
  NOR2_X1 U1101 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1102 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1103 ( .A(KEYINPUT115), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1104 ( .A1(n1008), .A2(n1007), .ZN(n1015) );
  XOR2_X1 U1105 ( .A(G2090), .B(G162), .Z(n1009) );
  NOR2_X1 U1106 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1107 ( .A(KEYINPUT51), .B(n1011), .Z(n1013) );
  NAND2_X1 U1108 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1109 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1110 ( .A(KEYINPUT52), .B(n1016), .ZN(n1018) );
  NAND2_X1 U1111 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1112 ( .A1(n1019), .A2(G29), .ZN(n1020) );
  NAND2_X1 U1113 ( .A1(n1021), .A2(n1020), .ZN(n1051) );
  XNOR2_X1 U1114 ( .A(n1022), .B(KEYINPUT56), .ZN(n1049) );
  NAND2_X1 U1115 ( .A1(G1971), .A2(G303), .ZN(n1023) );
  NAND2_X1 U1116 ( .A1(n1024), .A2(n1023), .ZN(n1034) );
  XOR2_X1 U1117 ( .A(G1961), .B(G171), .Z(n1025) );
  NOR2_X1 U1118 ( .A1(n1026), .A2(n1025), .ZN(n1032) );
  XOR2_X1 U1119 ( .A(n1027), .B(G1956), .Z(n1030) );
  XOR2_X1 U1120 ( .A(n1028), .B(G1348), .Z(n1029) );
  NOR2_X1 U1121 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1122 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1123 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1124 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1125 ( .A(KEYINPUT125), .B(n1037), .ZN(n1043) );
  XOR2_X1 U1126 ( .A(G1966), .B(G168), .Z(n1038) );
  XNOR2_X1 U1127 ( .A(KEYINPUT124), .B(n1038), .ZN(n1039) );
  NOR2_X1 U1128 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1129 ( .A(KEYINPUT57), .B(n1041), .Z(n1042) );
  NAND2_X1 U1130 ( .A1(n1043), .A2(n1042), .ZN(n1046) );
  XNOR2_X1 U1131 ( .A(G1341), .B(n1044), .ZN(n1045) );
  NOR2_X1 U1132 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  XNOR2_X1 U1133 ( .A(KEYINPUT126), .B(n1047), .ZN(n1048) );
  NOR2_X1 U1134 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  NOR2_X1 U1135 ( .A1(n1051), .A2(n1050), .ZN(n1052) );
  XOR2_X1 U1136 ( .A(n1052), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1137 ( .A(G150), .ZN(G311) );
endmodule

