

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  INV_X1 U323 ( .A(G190GAT), .ZN(n298) );
  XNOR2_X1 U324 ( .A(n374), .B(n300), .ZN(n301) );
  XNOR2_X1 U325 ( .A(n399), .B(n398), .ZN(n404) );
  AND2_X1 U326 ( .A1(G230GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U327 ( .A(n406), .B(KEYINPUT46), .ZN(n423) );
  NOR2_X1 U328 ( .A1(n555), .A2(n424), .ZN(n426) );
  XNOR2_X1 U329 ( .A(n389), .B(n291), .ZN(n391) );
  XNOR2_X1 U330 ( .A(n391), .B(n409), .ZN(n392) );
  XNOR2_X1 U331 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U332 ( .A(n397), .B(n396), .ZN(n398) );
  INV_X1 U333 ( .A(KEYINPUT102), .ZN(n427) );
  XNOR2_X1 U334 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n448) );
  XNOR2_X1 U335 ( .A(n427), .B(KEYINPUT36), .ZN(n428) );
  NOR2_X1 U336 ( .A1(n516), .A2(n447), .ZN(n566) );
  XNOR2_X1 U337 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U338 ( .A(n555), .B(n428), .ZN(n580) );
  NOR2_X1 U339 ( .A1(n531), .A2(n450), .ZN(n560) );
  XNOR2_X1 U340 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n451) );
  XNOR2_X1 U341 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT9), .B(KEYINPUT64), .Z(n293) );
  XNOR2_X1 U343 ( .A(G50GAT), .B(G106GAT), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n309) );
  XOR2_X1 U345 ( .A(G99GAT), .B(G85GAT), .Z(n389) );
  XOR2_X1 U346 ( .A(KEYINPUT10), .B(n389), .Z(n295) );
  XOR2_X1 U347 ( .A(G134GAT), .B(KEYINPUT79), .Z(n355) );
  XNOR2_X1 U348 ( .A(G36GAT), .B(n355), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n302) );
  XOR2_X1 U350 ( .A(G29GAT), .B(G43GAT), .Z(n297) );
  XNOR2_X1 U351 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n374) );
  NAND2_X1 U353 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XOR2_X1 U354 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U355 ( .A(G218GAT), .B(G162GAT), .Z(n333) );
  XOR2_X1 U356 ( .A(KEYINPUT78), .B(G92GAT), .Z(n304) );
  XNOR2_X1 U357 ( .A(KEYINPUT11), .B(KEYINPUT66), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n333), .B(n305), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n555) );
  XOR2_X1 U362 ( .A(KEYINPUT82), .B(KEYINPUT80), .Z(n311) );
  XNOR2_X1 U363 ( .A(G99GAT), .B(G134GAT), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U365 ( .A(n312), .B(KEYINPUT20), .Z(n314) );
  XOR2_X1 U366 ( .A(G120GAT), .B(G71GAT), .Z(n395) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(n395), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n319) );
  XNOR2_X1 U369 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n315), .B(G127GAT), .ZN(n359) );
  XOR2_X1 U371 ( .A(G15GAT), .B(n359), .Z(n317) );
  NAND2_X1 U372 ( .A1(G227GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U374 ( .A(n319), .B(n318), .Z(n328) );
  XNOR2_X1 U375 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n320), .B(KEYINPUT18), .ZN(n321) );
  XOR2_X1 U377 ( .A(n321), .B(KEYINPUT17), .Z(n323) );
  XNOR2_X1 U378 ( .A(G183GAT), .B(G190GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n435) );
  XOR2_X1 U380 ( .A(G176GAT), .B(KEYINPUT83), .Z(n325) );
  XNOR2_X1 U381 ( .A(G169GAT), .B(KEYINPUT65), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n435), .B(n326), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n531) );
  XNOR2_X1 U385 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n329), .B(KEYINPUT2), .ZN(n354) );
  XOR2_X1 U387 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n331) );
  XNOR2_X1 U388 ( .A(KEYINPUT23), .B(KEYINPUT85), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(n333), .B(n332), .Z(n335) );
  NAND2_X1 U391 ( .A1(G228GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U393 ( .A(G204GAT), .B(KEYINPUT24), .Z(n337) );
  XNOR2_X1 U394 ( .A(KEYINPUT88), .B(KEYINPUT84), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U396 ( .A(n339), .B(n338), .Z(n344) );
  XNOR2_X1 U397 ( .A(G50GAT), .B(G22GAT), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n340), .B(G141GAT), .ZN(n382) );
  XOR2_X1 U399 ( .A(G211GAT), .B(KEYINPUT21), .Z(n342) );
  XNOR2_X1 U400 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n436) );
  XNOR2_X1 U402 ( .A(n382), .B(n436), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n354), .B(n345), .ZN(n347) );
  XNOR2_X1 U405 ( .A(G106GAT), .B(G78GAT), .ZN(n346) );
  XOR2_X1 U406 ( .A(n346), .B(G148GAT), .Z(n402) );
  XNOR2_X1 U407 ( .A(n347), .B(n402), .ZN(n469) );
  XOR2_X1 U408 ( .A(G57GAT), .B(G148GAT), .Z(n349) );
  XNOR2_X1 U409 ( .A(G141GAT), .B(G1GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U411 ( .A(G85GAT), .B(G162GAT), .Z(n351) );
  XNOR2_X1 U412 ( .A(G29GAT), .B(G120GAT), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n371) );
  XOR2_X1 U415 ( .A(n355), .B(n354), .Z(n357) );
  NAND2_X1 U416 ( .A1(G225GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U418 ( .A(n358), .B(KEYINPUT93), .Z(n361) );
  XNOR2_X1 U419 ( .A(n359), .B(KEYINPUT89), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n369) );
  XOR2_X1 U421 ( .A(KEYINPUT94), .B(KEYINPUT6), .Z(n363) );
  XNOR2_X1 U422 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U424 ( .A(KEYINPUT90), .B(KEYINPUT4), .Z(n365) );
  XNOR2_X1 U425 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U427 ( .A(n367), .B(n366), .Z(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n371), .B(n370), .ZN(n516) );
  INV_X1 U430 ( .A(KEYINPUT54), .ZN(n446) );
  XOR2_X1 U431 ( .A(G197GAT), .B(G113GAT), .Z(n373) );
  XNOR2_X1 U432 ( .A(KEYINPUT72), .B(KEYINPUT29), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n386) );
  XOR2_X1 U434 ( .A(n374), .B(KEYINPUT67), .Z(n376) );
  NAND2_X1 U435 ( .A1(G229GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U437 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n378) );
  XNOR2_X1 U438 ( .A(KEYINPUT70), .B(KEYINPUT68), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U440 ( .A(n380), .B(n379), .Z(n384) );
  XNOR2_X1 U441 ( .A(G15GAT), .B(G1GAT), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n381), .B(KEYINPUT71), .ZN(n420) );
  XNOR2_X1 U443 ( .A(n382), .B(n420), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n388) );
  XOR2_X1 U446 ( .A(G169GAT), .B(G36GAT), .Z(n387) );
  XOR2_X1 U447 ( .A(G8GAT), .B(n387), .Z(n444) );
  XNOR2_X1 U448 ( .A(n388), .B(n444), .ZN(n567) );
  INV_X1 U449 ( .A(n567), .ZN(n405) );
  XNOR2_X1 U450 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n390), .B(KEYINPUT74), .ZN(n409) );
  XOR2_X1 U452 ( .A(n392), .B(KEYINPUT76), .Z(n399) );
  XOR2_X1 U453 ( .A(KEYINPUT75), .B(KEYINPUT77), .Z(n394) );
  XNOR2_X1 U454 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n393) );
  XOR2_X1 U455 ( .A(n394), .B(n393), .Z(n397) );
  XNOR2_X1 U456 ( .A(n395), .B(KEYINPUT32), .ZN(n396) );
  XOR2_X1 U457 ( .A(G64GAT), .B(G92GAT), .Z(n401) );
  XNOR2_X1 U458 ( .A(G176GAT), .B(G204GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n440) );
  XOR2_X1 U460 ( .A(n402), .B(n440), .Z(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n570) );
  XNOR2_X1 U462 ( .A(KEYINPUT41), .B(n570), .ZN(n547) );
  NAND2_X1 U463 ( .A1(n405), .A2(n547), .ZN(n406) );
  XOR2_X1 U464 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n412) );
  XOR2_X1 U465 ( .A(KEYINPUT15), .B(G64GAT), .Z(n408) );
  XNOR2_X1 U466 ( .A(G22GAT), .B(G8GAT), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U470 ( .A(G127GAT), .B(G183GAT), .Z(n414) );
  NAND2_X1 U471 ( .A1(G231GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U473 ( .A(n416), .B(n415), .Z(n422) );
  XOR2_X1 U474 ( .A(G211GAT), .B(G78GAT), .Z(n418) );
  XNOR2_X1 U475 ( .A(G71GAT), .B(G155GAT), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n574) );
  NAND2_X1 U479 ( .A1(n423), .A2(n574), .ZN(n424) );
  XNOR2_X1 U480 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n433) );
  XNOR2_X1 U482 ( .A(n567), .B(KEYINPUT73), .ZN(n558) );
  NOR2_X1 U483 ( .A1(n574), .A2(n580), .ZN(n429) );
  XNOR2_X1 U484 ( .A(KEYINPUT45), .B(n429), .ZN(n430) );
  NAND2_X1 U485 ( .A1(n430), .A2(n570), .ZN(n431) );
  NOR2_X1 U486 ( .A1(n558), .A2(n431), .ZN(n432) );
  NOR2_X1 U487 ( .A1(n433), .A2(n432), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n434), .B(KEYINPUT48), .ZN(n526) );
  INV_X1 U489 ( .A(n435), .ZN(n442) );
  XOR2_X1 U490 ( .A(G218GAT), .B(n436), .Z(n438) );
  NAND2_X1 U491 ( .A1(G226GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U493 ( .A(n440), .B(n439), .Z(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n464) );
  NOR2_X1 U496 ( .A1(n526), .A2(n464), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U498 ( .A1(n469), .A2(n566), .ZN(n449) );
  NAND2_X1 U499 ( .A1(n555), .A2(n560), .ZN(n452) );
  XOR2_X1 U500 ( .A(KEYINPUT107), .B(n547), .Z(n533) );
  NAND2_X1 U501 ( .A1(n560), .A2(n533), .ZN(n455) );
  XOR2_X1 U502 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n453) );
  XNOR2_X1 U503 ( .A(n453), .B(G176GAT), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  XOR2_X1 U505 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n476) );
  NAND2_X1 U506 ( .A1(n570), .A2(n558), .ZN(n488) );
  NOR2_X1 U507 ( .A1(n574), .A2(n555), .ZN(n456) );
  XNOR2_X1 U508 ( .A(n456), .B(KEYINPUT16), .ZN(n474) );
  INV_X1 U509 ( .A(n516), .ZN(n468) );
  INV_X1 U510 ( .A(n531), .ZN(n520) );
  INV_X1 U511 ( .A(n464), .ZN(n518) );
  NAND2_X1 U512 ( .A1(n520), .A2(n518), .ZN(n457) );
  NAND2_X1 U513 ( .A1(n457), .A2(n469), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n458), .B(KEYINPUT98), .ZN(n459) );
  XNOR2_X1 U515 ( .A(KEYINPUT25), .B(n459), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n460), .B(KEYINPUT97), .ZN(n466) );
  NOR2_X1 U517 ( .A1(n520), .A2(n469), .ZN(n462) );
  XNOR2_X1 U518 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U520 ( .A(KEYINPUT95), .B(n463), .Z(n565) );
  XOR2_X1 U521 ( .A(KEYINPUT27), .B(n464), .Z(n470) );
  NAND2_X1 U522 ( .A1(n565), .A2(n470), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U524 ( .A1(n468), .A2(n467), .ZN(n473) );
  XNOR2_X1 U525 ( .A(KEYINPUT28), .B(n469), .ZN(n529) );
  NAND2_X1 U526 ( .A1(n516), .A2(n470), .ZN(n527) );
  NOR2_X1 U527 ( .A1(n520), .A2(n527), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n529), .A2(n471), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n473), .A2(n472), .ZN(n485) );
  NAND2_X1 U530 ( .A1(n474), .A2(n485), .ZN(n502) );
  NOR2_X1 U531 ( .A1(n488), .A2(n502), .ZN(n482) );
  NAND2_X1 U532 ( .A1(n482), .A2(n516), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NAND2_X1 U535 ( .A1(n482), .A2(n518), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U538 ( .A1(n482), .A2(n520), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n481), .ZN(G1326GAT) );
  XOR2_X1 U541 ( .A(G22GAT), .B(KEYINPUT101), .Z(n484) );
  INV_X1 U542 ( .A(n529), .ZN(n523) );
  NAND2_X1 U543 ( .A1(n482), .A2(n523), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT104), .Z(n492) );
  NAND2_X1 U546 ( .A1(n574), .A2(n485), .ZN(n486) );
  NOR2_X1 U547 ( .A1(n580), .A2(n486), .ZN(n487) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n487), .ZN(n514) );
  NOR2_X1 U549 ( .A1(n514), .A2(n488), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT103), .B(KEYINPUT38), .Z(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(n498) );
  NAND2_X1 U552 ( .A1(n498), .A2(n516), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U554 ( .A(KEYINPUT39), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n498), .A2(n518), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n496) );
  NAND2_X1 U558 ( .A1(n498), .A2(n520), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  XNOR2_X1 U561 ( .A(G50GAT), .B(KEYINPUT106), .ZN(n500) );
  NAND2_X1 U562 ( .A1(n523), .A2(n498), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT42), .B(KEYINPUT110), .Z(n505) );
  NAND2_X1 U565 ( .A1(n533), .A2(n567), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n501), .B(KEYINPUT108), .ZN(n515) );
  NOR2_X1 U567 ( .A1(n515), .A2(n502), .ZN(n503) );
  XOR2_X1 U568 ( .A(KEYINPUT109), .B(n503), .Z(n509) );
  NAND2_X1 U569 ( .A1(n509), .A2(n516), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n506), .Z(G1332GAT) );
  NAND2_X1 U572 ( .A1(n509), .A2(n518), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n520), .A2(n509), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U577 ( .A1(n509), .A2(n523), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n513) );
  XOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT111), .Z(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n522) );
  NAND2_X1 U582 ( .A1(n522), .A2(n516), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n522), .A2(n518), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n520), .A2(n522), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(KEYINPUT114), .ZN(n544) );
  NAND2_X1 U593 ( .A1(n529), .A2(n544), .ZN(n530) );
  NOR2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n540), .A2(n558), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U598 ( .A1(n540), .A2(n533), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U600 ( .A(G120GAT), .B(n536), .Z(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n538) );
  INV_X1 U602 ( .A(n574), .ZN(n561) );
  NAND2_X1 U603 ( .A1(n540), .A2(n561), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U605 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U607 ( .A1(n540), .A2(n555), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U609 ( .A(G134GAT), .B(n543), .Z(G1343GAT) );
  NAND2_X1 U610 ( .A1(n565), .A2(n544), .ZN(n546) );
  NOR2_X1 U611 ( .A1(n567), .A2(n546), .ZN(n545) );
  XOR2_X1 U612 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  INV_X1 U614 ( .A(n546), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n554), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n552) );
  NAND2_X1 U619 ( .A1(n554), .A2(n561), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n553), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT120), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n560), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n564) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n579) );
  NOR2_X1 U633 ( .A1(n567), .A2(n579), .ZN(n568) );
  XOR2_X1 U634 ( .A(n569), .B(n568), .Z(G1352GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n579), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT123), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n579), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT124), .B(n575), .Z(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n578) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n582) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(n582), .B(n581), .Z(G1355GAT) );
endmodule

