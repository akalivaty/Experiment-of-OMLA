//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G134), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G137), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n189), .B1(KEYINPUT11), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G134), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  AOI211_X1 g010(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n188), .C2(G134), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n192), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G131), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n192), .B(new_n200), .C1(new_n196), .C2(new_n197), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(KEYINPUT65), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(new_n203), .A3(G131), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n205), .B(new_n207), .C1(new_n209), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(G146), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT0), .A4(G128), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n212), .A2(KEYINPUT67), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT67), .B1(new_n212), .B2(new_n215), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n202), .A2(new_n204), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n191), .A2(new_n189), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n201), .B1(new_n200), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n213), .A2(new_n214), .A3(new_n222), .A4(G128), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(G128), .B1(new_n213), .B2(new_n214), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n214), .A2(new_n222), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT66), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n229));
  XNOR2_X1  g043(.A(G143), .B(G146), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n228), .B(new_n229), .C1(new_n230), .C2(G128), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n224), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  OR2_X1    g046(.A1(new_n221), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n219), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g048(.A(G116), .B(G119), .Z(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT2), .B(G113), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n235), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n237), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n219), .A2(new_n233), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n187), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n241), .A2(new_n242), .B1(new_n187), .B2(new_n240), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT26), .B(G101), .Z(new_n246));
  XNOR2_X1  g060(.A(new_n246), .B(KEYINPUT69), .ZN(new_n247));
  NOR2_X1   g061(.A1(G237), .A2(G953), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G210), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n247), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT29), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n244), .A2(new_n245), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G902), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n240), .A2(new_n187), .ZN(new_n257));
  INV_X1    g071(.A(new_n205), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n230), .A2(new_n258), .A3(new_n206), .ZN(new_n259));
  INV_X1    g073(.A(new_n215), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n202), .A2(new_n261), .A3(new_n204), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n233), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n237), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n219), .A2(new_n233), .A3(KEYINPUT28), .A4(new_n239), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n257), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n253), .B1(new_n266), .B2(new_n252), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n250), .B(new_n251), .Z(new_n268));
  INV_X1    g082(.A(KEYINPUT30), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n219), .A2(new_n233), .A3(KEYINPUT30), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n237), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n268), .B1(new_n272), .B2(new_n240), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n256), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(G472), .B1(new_n255), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n268), .A3(new_n240), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT31), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT70), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n266), .A2(new_n252), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n272), .A2(new_n268), .A3(new_n240), .A4(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n279), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(G472), .A2(G902), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g100(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n284), .A2(KEYINPUT32), .A3(new_n285), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n275), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT15), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G478), .ZN(new_n293));
  XNOR2_X1  g107(.A(G128), .B(G143), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n294), .B(new_n190), .ZN(new_n295));
  INV_X1    g109(.A(G128), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G143), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT13), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(G134), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n294), .A2(new_n298), .A3(G134), .A4(new_n297), .ZN(new_n301));
  INV_X1    g115(.A(G107), .ZN(new_n302));
  INV_X1    g116(.A(G122), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT90), .B1(new_n303), .B2(G116), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT90), .ZN(new_n305));
  INV_X1    g119(.A(G116), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(G122), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n306), .A2(G122), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n302), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n308), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n312), .A2(G107), .A3(new_n309), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n300), .B(new_n301), .C1(new_n311), .C2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  INV_X1    g129(.A(G217), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n315), .A2(new_n316), .A3(G953), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT14), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(new_n304), .B2(new_n307), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(new_n309), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n320), .A2(KEYINPUT91), .B1(new_n318), .B2(new_n312), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT91), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n319), .B2(new_n309), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n302), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n294), .B(G134), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n313), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n314), .B(new_n317), .C1(new_n324), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT92), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n320), .A2(KEYINPUT91), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n312), .A2(new_n318), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n323), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G107), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n326), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT92), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n335), .A3(new_n314), .A4(new_n317), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n314), .B1(new_n324), .B2(new_n327), .ZN(new_n337));
  INV_X1    g151(.A(new_n317), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n329), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT94), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n256), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT93), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT93), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n344), .A3(new_n256), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n293), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT20), .ZN(new_n347));
  NOR2_X1   g161(.A1(G475), .A2(G902), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n248), .A2(G214), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n208), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n248), .A2(G143), .A3(G214), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G131), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT17), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n200), .A3(new_n351), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(KEYINPUT74), .A2(G125), .ZN(new_n357));
  INV_X1    g171(.A(G140), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(KEYINPUT74), .A2(G125), .A3(G140), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(KEYINPUT16), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT16), .ZN(new_n362));
  INV_X1    g176(.A(G125), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(G140), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n210), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n364), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G146), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n352), .A2(KEYINPUT17), .A3(G131), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n356), .A2(new_n365), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  AND2_X1   g183(.A1(KEYINPUT18), .A2(G131), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n352), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n359), .A2(new_n360), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G146), .ZN(new_n373));
  XNOR2_X1  g187(.A(G125), .B(G140), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT76), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n374), .A2(new_n375), .A3(new_n210), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n375), .B1(new_n374), .B2(new_n210), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n352), .A2(new_n370), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n371), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  XOR2_X1   g194(.A(G113), .B(G122), .Z(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT88), .B(G104), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n369), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n353), .A2(new_n355), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n367), .A2(KEYINPUT75), .ZN(new_n387));
  XOR2_X1   g201(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n388));
  AOI22_X1  g202(.A1(new_n372), .A2(KEYINPUT19), .B1(new_n388), .B2(new_n374), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n210), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT75), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n366), .A2(new_n391), .A3(G146), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n386), .A2(new_n387), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n383), .B1(new_n393), .B2(new_n380), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n347), .B(new_n348), .C1(new_n385), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT89), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n393), .A2(new_n380), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n384), .B1(new_n397), .B2(new_n383), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT89), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n398), .A2(new_n399), .A3(new_n347), .A4(new_n348), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n348), .B1(new_n385), .B2(new_n394), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT20), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n396), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n383), .B1(new_n369), .B2(new_n380), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n256), .B1(new_n385), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G475), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n342), .A2(KEYINPUT93), .B1(new_n292), .B2(G478), .ZN(new_n408));
  INV_X1    g222(.A(G953), .ZN(new_n409));
  INV_X1    g223(.A(G952), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n410), .A2(KEYINPUT95), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(KEYINPUT95), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(G234), .B2(G237), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT21), .B(G898), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n256), .B(new_n409), .C1(G234), .C2(G237), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR4_X1   g231(.A1(new_n346), .A2(new_n407), .A3(new_n408), .A4(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(KEYINPUT24), .B(G110), .Z(new_n419));
  XNOR2_X1  g233(.A(G119), .B(G128), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n421), .B(KEYINPUT73), .Z(new_n422));
  NAND2_X1  g236(.A1(new_n367), .A2(new_n365), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT23), .ZN(new_n424));
  INV_X1    g238(.A(G119), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n424), .B1(new_n425), .B2(G128), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n296), .A2(KEYINPUT23), .A3(G119), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n426), .B(new_n427), .C1(G119), .C2(new_n296), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G110), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n422), .A2(new_n423), .A3(new_n429), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n376), .A2(new_n377), .ZN(new_n431));
  OAI22_X1  g245(.A1(new_n428), .A2(G110), .B1(new_n420), .B2(new_n419), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n387), .A2(new_n431), .A3(new_n392), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT22), .B(G137), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n409), .A2(G221), .A3(G234), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n435), .B(new_n436), .Z(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n430), .B2(new_n433), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n316), .B1(G234), .B2(new_n256), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G902), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n256), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT25), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n444), .B1(new_n447), .B2(new_n442), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n291), .A2(new_n418), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G469), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G140), .ZN(new_n451));
  INV_X1    g265(.A(G227), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G953), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n451), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT79), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT67), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n259), .B2(new_n260), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n302), .A2(KEYINPUT78), .A3(G104), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT3), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n460), .A2(new_n302), .A3(KEYINPUT78), .A4(G104), .ZN(new_n461));
  INV_X1    g275(.A(G104), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G107), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT4), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n465), .A3(G101), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n212), .A2(KEYINPUT67), .A3(new_n215), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n457), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G101), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n459), .A2(new_n469), .A3(new_n461), .A4(new_n463), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT4), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n458), .A2(KEYINPUT3), .B1(new_n462), .B2(G107), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n469), .B1(new_n472), .B2(new_n461), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n455), .B1(new_n468), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n464), .A2(G101), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(KEYINPUT4), .A3(new_n470), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n218), .A2(KEYINPUT79), .A3(new_n477), .A4(new_n466), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n202), .A2(new_n204), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n223), .B(new_n228), .C1(G128), .C2(new_n230), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT80), .B1(new_n302), .B2(G104), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT80), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n462), .A3(G107), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n482), .B(new_n484), .C1(new_n462), .C2(G107), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G101), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n481), .A2(new_n470), .A3(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(KEYINPUT10), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n470), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT10), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n232), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n479), .A2(new_n480), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n480), .B1(new_n479), .B2(new_n492), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n454), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT82), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n202), .A2(new_n204), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT12), .ZN(new_n498));
  INV_X1    g312(.A(new_n487), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n232), .A2(new_n489), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n487), .B1(new_n232), .B2(new_n489), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT12), .B1(new_n503), .B2(new_n480), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n493), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n454), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n495), .A2(new_n496), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n479), .A2(new_n480), .A3(new_n492), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n504), .A3(new_n502), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n510), .A2(KEYINPUT82), .A3(new_n454), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n450), .B(new_n256), .C1(new_n508), .C2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n450), .A2(new_n256), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT81), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n493), .B2(new_n505), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n509), .A2(KEYINPUT81), .A3(new_n504), .A4(new_n502), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n454), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n493), .A2(new_n494), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n507), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n512), .B(new_n514), .C1(new_n450), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n232), .A2(new_n363), .ZN(new_n523));
  OAI21_X1  g337(.A(G125), .B1(new_n259), .B2(new_n260), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n409), .A2(G224), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n525), .B(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n237), .B(new_n466), .C1(new_n473), .C2(new_n471), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT5), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n425), .A3(G116), .ZN(new_n531));
  OAI211_X1 g345(.A(G113), .B(new_n531), .C1(new_n235), .C2(new_n530), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n235), .A2(new_n236), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n532), .A2(new_n533), .A3(new_n486), .A4(new_n470), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(G110), .B(G122), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n529), .A2(new_n534), .A3(new_n536), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(KEYINPUT6), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n536), .B1(new_n529), .B2(new_n534), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT6), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n541), .A2(KEYINPUT83), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT83), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n528), .B(new_n540), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(G210), .B1(G237), .B2(G902), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT86), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT84), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT7), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n527), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n549), .B2(new_n550), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n525), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT85), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT7), .B1(new_n526), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n554), .B2(new_n526), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n523), .A2(new_n524), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n536), .B(KEYINPUT8), .ZN(new_n558));
  INV_X1    g372(.A(new_n534), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n533), .A2(new_n532), .B1(new_n486), .B2(new_n470), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n553), .A2(new_n557), .A3(new_n561), .A4(new_n539), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n562), .A2(new_n256), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n545), .A2(new_n548), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n548), .B1(new_n545), .B2(new_n563), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G214), .B1(G237), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G221), .ZN(new_n570));
  INV_X1    g384(.A(new_n315), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n571), .B2(new_n256), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n572), .B(KEYINPUT77), .Z(new_n573));
  NAND3_X1  g387(.A1(new_n522), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n449), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT96), .B(G101), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(G3));
  AND2_X1   g391(.A1(new_n522), .A2(new_n573), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n284), .A2(new_n256), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n579), .A2(G472), .B1(new_n284), .B2(new_n285), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n580), .A2(new_n448), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n545), .A2(new_n563), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n547), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n545), .A2(new_n563), .A3(new_n548), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n545), .A2(new_n563), .A3(KEYINPUT97), .A4(new_n548), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n587), .A2(new_n567), .ZN(new_n588));
  INV_X1    g402(.A(new_n417), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n337), .B2(new_n338), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n340), .A2(new_n591), .B1(new_n328), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(G478), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(G902), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n340), .A2(new_n256), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n594), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n407), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n590), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n578), .A2(new_n581), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G104), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  AOI22_X1  g419(.A1(new_n402), .A2(new_n395), .B1(G475), .B2(new_n405), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n346), .B2(new_n408), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n590), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n578), .A2(new_n581), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G107), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  NAND4_X1  g425(.A1(new_n522), .A2(new_n580), .A3(new_n569), .A4(new_n573), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n445), .A2(new_n446), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT25), .B1(new_n441), .B2(new_n256), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n442), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n438), .A2(KEYINPUT36), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n434), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n443), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n418), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT37), .B(G110), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G12));
  NOR2_X1   g437(.A1(new_n346), .A2(new_n408), .ZN(new_n624));
  INV_X1    g438(.A(G900), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n414), .B1(new_n625), .B2(new_n416), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n606), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n619), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n586), .A2(new_n588), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n578), .A2(new_n291), .A3(new_n629), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G128), .ZN(G30));
  INV_X1    g448(.A(new_n408), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n340), .A2(new_n344), .A3(new_n256), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(KEYINPUT93), .B2(new_n342), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n635), .B1(new_n637), .B2(new_n293), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n630), .A2(new_n638), .A3(new_n567), .A4(new_n407), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n640), .A2(KEYINPUT100), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(KEYINPUT100), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n583), .A2(new_n585), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT38), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n272), .A2(new_n240), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n252), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n238), .A2(new_n240), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(KEYINPUT99), .A3(new_n252), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT99), .B1(new_n647), .B2(new_n252), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(G472), .B1(new_n651), .B2(G902), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n289), .A2(new_n652), .A3(new_n290), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n641), .A2(new_n642), .A3(new_n644), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n626), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n578), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT102), .Z(new_n658));
  AOI21_X1  g472(.A(new_n654), .B1(new_n658), .B2(KEYINPUT40), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n659), .B1(KEYINPUT40), .B2(new_n658), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G143), .ZN(G45));
  NAND3_X1  g475(.A1(new_n599), .A2(new_n407), .A3(new_n627), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n578), .A2(new_n291), .A3(new_n632), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G146), .ZN(G48));
  INV_X1    g479(.A(new_n572), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n508), .A2(new_n511), .ZN(new_n667));
  OAI21_X1  g481(.A(G469), .B1(new_n667), .B2(G902), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n601), .A2(new_n512), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n291), .A2(new_n448), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT41), .B(G113), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G15));
  NAND4_X1  g487(.A1(new_n608), .A2(new_n512), .A3(new_n666), .A4(new_n668), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n670), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n306), .ZN(G18));
  NAND2_X1  g490(.A1(new_n587), .A2(new_n567), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n566), .B2(new_n584), .ZN(new_n678));
  AND4_X1   g492(.A1(new_n512), .A2(new_n668), .A3(new_n666), .A4(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n418), .A2(new_n619), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n680), .A3(new_n291), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G119), .ZN(G21));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT104), .B(G472), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n579), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n285), .B(KEYINPUT103), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n268), .B1(new_n244), .B2(new_n245), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n279), .A2(new_n283), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n448), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT105), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n407), .B1(new_n346), .B2(new_n408), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n692), .B1(new_n693), .B2(new_n631), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n638), .A2(new_n678), .A3(KEYINPUT106), .A4(new_n407), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n668), .A2(new_n512), .A3(new_n666), .A4(new_n589), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n683), .B1(new_n691), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n690), .B(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n697), .B1(new_n694), .B2(new_n695), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(KEYINPUT107), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NAND2_X1  g520(.A1(new_n685), .A2(new_n689), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n707), .A2(new_n630), .A3(new_n662), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n679), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT108), .B(G125), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G27));
  INV_X1    g525(.A(new_n670), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n643), .A2(new_n568), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n518), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n507), .B1(new_n510), .B2(new_n515), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n717), .A2(new_n517), .B1(new_n519), .B2(new_n507), .ZN(new_n718));
  OAI211_X1 g532(.A(G469), .B(new_n716), .C1(new_n718), .C2(new_n715), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n512), .A4(new_n514), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n479), .A2(new_n492), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n497), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n507), .B1(new_n724), .B2(new_n509), .ZN(new_n725));
  OAI22_X1  g539(.A1(new_n725), .A2(KEYINPUT82), .B1(new_n454), .B2(new_n510), .ZN(new_n726));
  INV_X1    g540(.A(new_n511), .ZN(new_n727));
  AOI21_X1  g541(.A(G902), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n513), .B1(new_n728), .B2(new_n450), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n720), .B1(new_n729), .B2(new_n719), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n666), .B1(new_n722), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n714), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n512), .A2(new_n514), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n715), .B1(new_n518), .B2(new_n520), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT109), .B1(new_n717), .B2(new_n517), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n735), .A2(new_n450), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT110), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n572), .B1(new_n738), .B2(new_n721), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT111), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT112), .B1(new_n733), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n713), .B1(new_n739), .B2(KEYINPUT111), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n732), .B(new_n572), .C1(new_n738), .C2(new_n721), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n712), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n662), .A2(KEYINPUT42), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n275), .A2(new_n290), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT32), .B1(new_n284), .B2(new_n285), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n448), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n751), .A2(new_n662), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n731), .A2(new_n732), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(KEYINPUT112), .A3(new_n740), .A4(new_n713), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  OAI22_X1  g571(.A1(new_n746), .A2(new_n748), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n200), .ZN(G33));
  OAI211_X1 g573(.A(new_n712), .B(new_n629), .C1(new_n741), .C2(new_n745), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  AOI21_X1  g575(.A(new_n407), .B1(new_n598), .B2(new_n596), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT43), .ZN(new_n763));
  INV_X1    g577(.A(new_n580), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n619), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n763), .A2(KEYINPUT44), .A3(new_n764), .A4(new_n619), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n713), .A3(new_n768), .ZN(new_n769));
  OAI211_X1 g583(.A(KEYINPUT45), .B(new_n716), .C1(new_n718), .C2(new_n715), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n450), .B1(new_n521), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n513), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(KEYINPUT46), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n512), .B1(new_n773), .B2(KEYINPUT46), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n666), .B(new_n656), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n769), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n188), .ZN(G39));
  OR4_X1    g592(.A1(new_n291), .A2(new_n448), .A3(new_n662), .A4(new_n714), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n666), .B1(new_n774), .B2(new_n775), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n780), .A2(new_n782), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n779), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n358), .ZN(G42));
  AND2_X1   g600(.A1(new_n668), .A2(new_n512), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n790));
  INV_X1    g604(.A(new_n653), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n448), .A2(new_n762), .A3(new_n567), .A4(new_n573), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n644), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n789), .A2(new_n790), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n763), .A2(new_n414), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n691), .A2(new_n795), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n788), .A2(new_n567), .A3(new_n572), .A4(new_n644), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT50), .Z(new_n799));
  NAND3_X1  g613(.A1(new_n787), .A2(new_n666), .A3(new_n713), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n414), .A3(new_n448), .A4(new_n791), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n802), .A2(new_n407), .A3(new_n599), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n685), .A2(new_n619), .A3(new_n689), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n795), .A2(new_n800), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT114), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n799), .B(new_n803), .C1(new_n804), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT115), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n783), .B(new_n784), .C1(new_n573), .C2(new_n788), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(KEYINPUT116), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n691), .A2(new_n714), .A3(new_n795), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n809), .B2(KEYINPUT116), .ZN(new_n812));
  AND2_X1   g626(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n813));
  OAI221_X1 g627(.A(new_n808), .B1(new_n810), .B2(new_n812), .C1(new_n807), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n796), .A2(new_n679), .ZN(new_n815));
  INV_X1    g629(.A(new_n413), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n815), .B(new_n816), .C1(new_n600), .C2(new_n802), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n806), .A2(new_n751), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n818), .A2(KEYINPUT48), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(KEYINPUT48), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n807), .B1(new_n809), .B2(new_n811), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n814), .B(new_n821), .C1(KEYINPUT51), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n753), .A2(new_n755), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n708), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n346), .A2(new_n408), .A3(new_n407), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n407), .A2(new_n598), .A3(new_n596), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n643), .A2(new_n567), .A3(new_n589), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n578), .A2(new_n581), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n681), .A2(new_n830), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n449), .A2(new_n574), .B1(new_n612), .B2(new_n620), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n670), .B1(new_n674), .B2(new_n669), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n630), .A2(new_n714), .A3(new_n628), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n578), .A2(new_n835), .A3(new_n624), .A4(new_n291), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n834), .A2(new_n705), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n653), .A2(new_n630), .A3(new_n627), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n739), .A2(new_n839), .A3(new_n696), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n633), .A2(new_n664), .A3(new_n709), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n633), .A2(new_n709), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(KEYINPUT52), .A3(new_n664), .A4(new_n840), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n760), .A2(new_n825), .A3(new_n837), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n752), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n824), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n670), .B1(new_n753), .B2(new_n755), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n849), .A2(KEYINPUT42), .B1(new_n850), .B2(new_n747), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT53), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n760), .A2(new_n825), .A3(new_n837), .A4(new_n846), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n844), .A2(new_n838), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n853), .A2(new_n758), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT54), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n854), .A2(KEYINPUT53), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n847), .A2(new_n851), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n855), .B1(new_n853), .B2(new_n758), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n823), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(G952), .A2(G953), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n794), .B1(new_n866), .B2(new_n867), .ZN(G75));
  NOR2_X1   g682(.A1(new_n409), .A2(G952), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n256), .B1(new_n861), .B2(new_n862), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT56), .B1(new_n871), .B2(new_n547), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(new_n528), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT55), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n870), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n872), .A2(new_n875), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n872), .A2(KEYINPUT117), .A3(new_n875), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(G51));
  NOR3_X1   g695(.A1(new_n853), .A2(new_n758), .A3(new_n859), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT54), .B1(new_n852), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n864), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n861), .A2(new_n862), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n513), .B(KEYINPUT57), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n667), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n871), .A2(new_n770), .A3(new_n772), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n869), .B1(new_n891), .B2(new_n892), .ZN(G54));
  NAND2_X1  g707(.A1(KEYINPUT58), .A2(G475), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT119), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n871), .A2(new_n398), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n398), .B1(new_n871), .B2(new_n895), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n869), .ZN(G60));
  XNOR2_X1  g712(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n594), .A2(new_n256), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n899), .B(new_n900), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n858), .B2(new_n864), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n870), .B1(new_n903), .B2(new_n593), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n593), .A2(new_n901), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n885), .A2(new_n887), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n885), .A2(KEYINPUT121), .A3(new_n887), .A4(new_n905), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(G63));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT60), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n861), .B2(new_n862), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n617), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n441), .B(KEYINPUT122), .Z(new_n915));
  OAI211_X1 g729(.A(new_n914), .B(new_n870), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(G66));
  INV_X1    g732(.A(G224), .ZN(new_n919));
  OAI21_X1  g733(.A(G953), .B1(new_n415), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n834), .A2(new_n705), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n922), .B2(G953), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n873), .B1(G898), .B2(new_n409), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(G69));
  NAND2_X1  g739(.A1(new_n270), .A2(new_n271), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT124), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n389), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT125), .Z(new_n929));
  INV_X1    g743(.A(new_n842), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n660), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT62), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n660), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  OR4_X1    g748(.A1(new_n826), .A2(new_n670), .A3(new_n714), .A4(new_n827), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n658), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n936), .A2(new_n785), .A3(new_n777), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n932), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n929), .B1(new_n938), .B2(new_n409), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n625), .A2(G953), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT126), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n696), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n776), .A2(new_n943), .A3(new_n751), .ZN(new_n944));
  NOR4_X1   g758(.A1(new_n785), .A2(new_n777), .A3(new_n842), .A4(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n851), .A2(new_n945), .A3(new_n760), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n946), .B2(new_n409), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(KEYINPUT127), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n928), .B1(new_n947), .B2(KEYINPUT127), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n939), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(G953), .B1(new_n452), .B2(new_n625), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G72));
  NAND2_X1  g766(.A1(G472), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT63), .Z(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n938), .B2(new_n921), .ZN(new_n955));
  INV_X1    g769(.A(new_n645), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n252), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n852), .A2(new_n857), .ZN(new_n959));
  INV_X1    g773(.A(new_n957), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n956), .A2(new_n252), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n961), .A3(new_n954), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n946), .A2(new_n921), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n961), .B1(new_n964), .B2(new_n954), .ZN(new_n965));
  NOR4_X1   g779(.A1(new_n958), .A2(new_n869), .A3(new_n963), .A4(new_n965), .ZN(G57));
endmodule


