

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577;

  INV_X1 U317 ( .A(KEYINPUT26), .ZN(n393) );
  INV_X1 U318 ( .A(n421), .ZN(n296) );
  XNOR2_X1 U319 ( .A(n367), .B(n340), .ZN(n522) );
  XOR2_X1 U320 ( .A(n335), .B(n334), .Z(n285) );
  XNOR2_X1 U321 ( .A(n289), .B(n288), .ZN(n290) );
  XNOR2_X1 U322 ( .A(n343), .B(n290), .ZN(n292) );
  XNOR2_X1 U323 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n458) );
  XNOR2_X1 U324 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U325 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U326 ( .A(n299), .B(n298), .ZN(n304) );
  XNOR2_X1 U327 ( .A(n394), .B(n393), .ZN(n559) );
  XOR2_X1 U328 ( .A(KEYINPUT38), .B(n441), .Z(n491) );
  XNOR2_X1 U329 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U330 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n442) );
  XNOR2_X1 U331 ( .A(n471), .B(n470), .ZN(G1351GAT) );
  XNOR2_X1 U332 ( .A(n443), .B(n442), .ZN(G1330GAT) );
  XOR2_X1 U333 ( .A(G64GAT), .B(G92GAT), .Z(n287) );
  XNOR2_X1 U334 ( .A(G176GAT), .B(G204GAT), .ZN(n286) );
  XNOR2_X1 U335 ( .A(n287), .B(n286), .ZN(n343) );
  NAND2_X1 U336 ( .A1(G230GAT), .A2(G233GAT), .ZN(n289) );
  INV_X1 U337 ( .A(KEYINPUT33), .ZN(n288) );
  INV_X1 U338 ( .A(KEYINPUT32), .ZN(n291) );
  NAND2_X1 U339 ( .A1(n292), .A2(n291), .ZN(n295) );
  INV_X1 U340 ( .A(n292), .ZN(n293) );
  NAND2_X1 U341 ( .A1(n293), .A2(KEYINPUT32), .ZN(n294) );
  NAND2_X1 U342 ( .A1(n295), .A2(n294), .ZN(n299) );
  XOR2_X1 U343 ( .A(G57GAT), .B(KEYINPUT13), .Z(n406) );
  XNOR2_X1 U344 ( .A(n406), .B(KEYINPUT31), .ZN(n297) );
  XOR2_X1 U345 ( .A(G99GAT), .B(G85GAT), .Z(n421) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G71GAT), .Z(n335) );
  XOR2_X1 U347 ( .A(G148GAT), .B(G106GAT), .Z(n301) );
  XNOR2_X1 U348 ( .A(KEYINPUT70), .B(G78GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U350 ( .A(KEYINPUT69), .B(n302), .ZN(n388) );
  XOR2_X1 U351 ( .A(n335), .B(n388), .Z(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n566) );
  XNOR2_X1 U353 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n305), .B(G29GAT), .ZN(n306) );
  XOR2_X1 U355 ( .A(n306), .B(KEYINPUT7), .Z(n308) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G50GAT), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n435) );
  XOR2_X1 U358 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n310) );
  NAND2_X1 U359 ( .A1(G229GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U361 ( .A(n311), .B(KEYINPUT30), .Z(n315) );
  XNOR2_X1 U362 ( .A(G22GAT), .B(G197GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n312), .B(G141GAT), .ZN(n383) );
  XNOR2_X1 U364 ( .A(G15GAT), .B(G1GAT), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n313), .B(KEYINPUT67), .ZN(n407) );
  XNOR2_X1 U366 ( .A(n383), .B(n407), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U368 ( .A(n316), .B(KEYINPUT66), .Z(n318) );
  XOR2_X1 U369 ( .A(G169GAT), .B(G8GAT), .Z(n351) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(n351), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n435), .B(n319), .ZN(n561) );
  XOR2_X1 U373 ( .A(KEYINPUT68), .B(n561), .Z(n525) );
  OR2_X1 U374 ( .A1(n566), .A2(n525), .ZN(n478) );
  XOR2_X1 U375 ( .A(KEYINPUT37), .B(KEYINPUT97), .Z(n440) );
  XOR2_X1 U376 ( .A(KEYINPUT76), .B(G134GAT), .Z(n321) );
  XNOR2_X1 U377 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n320) );
  XNOR2_X1 U378 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U379 ( .A(G113GAT), .B(n322), .Z(n367) );
  XOR2_X1 U380 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n324) );
  XNOR2_X1 U381 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U383 ( .A(G176GAT), .B(KEYINPUT82), .Z(n326) );
  XNOR2_X1 U384 ( .A(G169GAT), .B(KEYINPUT78), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U386 ( .A(n328), .B(n327), .Z(n339) );
  XOR2_X1 U387 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n330) );
  XNOR2_X1 U388 ( .A(KEYINPUT80), .B(G183GAT), .ZN(n329) );
  XNOR2_X1 U389 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U390 ( .A(KEYINPUT18), .B(n331), .Z(n350) );
  XOR2_X1 U391 ( .A(KEYINPUT77), .B(G190GAT), .Z(n333) );
  XNOR2_X1 U392 ( .A(G43GAT), .B(G99GAT), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n334) );
  NAND2_X1 U394 ( .A1(G227GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n285), .B(n336), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n350), .B(n337), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U398 ( .A(G197GAT), .B(KEYINPUT90), .Z(n342) );
  NAND2_X1 U399 ( .A1(G226GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n344) );
  XOR2_X1 U401 ( .A(n344), .B(n343), .Z(n348) );
  XOR2_X1 U402 ( .A(G211GAT), .B(KEYINPUT86), .Z(n346) );
  XNOR2_X1 U403 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n382) );
  XNOR2_X1 U405 ( .A(G36GAT), .B(n382), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U407 ( .A(G190GAT), .B(KEYINPUT73), .Z(n422) );
  XOR2_X1 U408 ( .A(n349), .B(n422), .Z(n353) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n512) );
  XNOR2_X1 U411 ( .A(n512), .B(KEYINPUT27), .ZN(n395) );
  XOR2_X1 U412 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n355) );
  XNOR2_X1 U413 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n371) );
  XOR2_X1 U415 ( .A(G85GAT), .B(G120GAT), .Z(n357) );
  XNOR2_X1 U416 ( .A(G29GAT), .B(G141GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U418 ( .A(KEYINPUT6), .B(G57GAT), .Z(n359) );
  XNOR2_X1 U419 ( .A(G1GAT), .B(G148GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U421 ( .A(n361), .B(n360), .Z(n369) );
  XOR2_X1 U422 ( .A(G155GAT), .B(KEYINPUT3), .Z(n363) );
  XNOR2_X1 U423 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n373) );
  XOR2_X1 U425 ( .A(n373), .B(KEYINPUT5), .Z(n365) );
  NAND2_X1 U426 ( .A1(G225GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U430 ( .A(n371), .B(n370), .Z(n510) );
  NAND2_X1 U431 ( .A1(n395), .A2(n510), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n372), .B(KEYINPUT91), .ZN(n539) );
  XOR2_X1 U433 ( .A(n373), .B(G204GAT), .Z(n375) );
  NAND2_X1 U434 ( .A1(G228GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n387) );
  XOR2_X1 U436 ( .A(KEYINPUT85), .B(KEYINPUT23), .Z(n377) );
  XNOR2_X1 U437 ( .A(G50GAT), .B(KEYINPUT83), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U439 ( .A(KEYINPUT24), .B(KEYINPUT84), .Z(n379) );
  XNOR2_X1 U440 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U442 ( .A(n381), .B(n380), .Z(n385) );
  XNOR2_X1 U443 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n461) );
  XNOR2_X1 U447 ( .A(KEYINPUT28), .B(n461), .ZN(n485) );
  NAND2_X1 U448 ( .A1(n539), .A2(n485), .ZN(n524) );
  XNOR2_X1 U449 ( .A(KEYINPUT92), .B(n524), .ZN(n390) );
  NOR2_X1 U450 ( .A1(n522), .A2(n390), .ZN(n402) );
  NAND2_X1 U451 ( .A1(n512), .A2(n522), .ZN(n391) );
  NAND2_X1 U452 ( .A1(n461), .A2(n391), .ZN(n392) );
  XNOR2_X1 U453 ( .A(KEYINPUT25), .B(n392), .ZN(n399) );
  NOR2_X1 U454 ( .A1(n522), .A2(n461), .ZN(n394) );
  INV_X1 U455 ( .A(n395), .ZN(n396) );
  NOR2_X1 U456 ( .A1(n559), .A2(n396), .ZN(n397) );
  XOR2_X1 U457 ( .A(KEYINPUT93), .B(n397), .Z(n398) );
  NOR2_X1 U458 ( .A1(n399), .A2(n398), .ZN(n400) );
  NOR2_X1 U459 ( .A1(n510), .A2(n400), .ZN(n401) );
  NOR2_X1 U460 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n403), .B(KEYINPUT94), .ZN(n475) );
  XOR2_X1 U462 ( .A(G155GAT), .B(G211GAT), .Z(n405) );
  XNOR2_X1 U463 ( .A(G22GAT), .B(G71GAT), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n420) );
  XOR2_X1 U465 ( .A(n406), .B(G183GAT), .Z(n409) );
  XNOR2_X1 U466 ( .A(n407), .B(G127GAT), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U468 ( .A(KEYINPUT74), .B(KEYINPUT12), .Z(n411) );
  NAND2_X1 U469 ( .A1(G231GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U471 ( .A(n413), .B(n412), .Z(n418) );
  XOR2_X1 U472 ( .A(KEYINPUT14), .B(G64GAT), .Z(n415) );
  XNOR2_X1 U473 ( .A(G8GAT), .B(G78GAT), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n416), .B(KEYINPUT15), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n570) );
  NOR2_X1 U478 ( .A1(n475), .A2(n570), .ZN(n438) );
  XOR2_X1 U479 ( .A(KEYINPUT9), .B(KEYINPUT71), .Z(n424) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U482 ( .A(KEYINPUT64), .B(G92GAT), .Z(n426) );
  XNOR2_X1 U483 ( .A(G134GAT), .B(G106GAT), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U485 ( .A(n428), .B(n427), .Z(n430) );
  XNOR2_X1 U486 ( .A(G218GAT), .B(G162GAT), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U488 ( .A(KEYINPUT72), .B(KEYINPUT10), .Z(n432) );
  NAND2_X1 U489 ( .A1(G232GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n437) );
  XOR2_X1 U492 ( .A(n435), .B(KEYINPUT11), .Z(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n550) );
  XNOR2_X1 U494 ( .A(KEYINPUT36), .B(n550), .ZN(n573) );
  NAND2_X1 U495 ( .A1(n438), .A2(n573), .ZN(n439) );
  XOR2_X1 U496 ( .A(n440), .B(n439), .Z(n509) );
  OR2_X1 U497 ( .A1(n478), .A2(n509), .ZN(n441) );
  NAND2_X1 U498 ( .A1(n491), .A2(n522), .ZN(n443) );
  XOR2_X1 U499 ( .A(n566), .B(KEYINPUT41), .Z(n544) );
  NAND2_X1 U500 ( .A1(n544), .A2(n561), .ZN(n446) );
  XOR2_X1 U501 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n444) );
  XNOR2_X1 U502 ( .A(KEYINPUT108), .B(n444), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n448) );
  NOR2_X1 U504 ( .A1(n550), .A2(n570), .ZN(n447) );
  AND2_X1 U505 ( .A1(n448), .A2(n447), .ZN(n450) );
  XNOR2_X1 U506 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n456) );
  XNOR2_X1 U508 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n452) );
  NAND2_X1 U509 ( .A1(n570), .A2(n573), .ZN(n451) );
  XOR2_X1 U510 ( .A(n452), .B(n451), .Z(n453) );
  NOR2_X1 U511 ( .A1(n566), .A2(n453), .ZN(n454) );
  NAND2_X1 U512 ( .A1(n525), .A2(n454), .ZN(n455) );
  NAND2_X1 U513 ( .A1(n456), .A2(n455), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n457), .B(KEYINPUT48), .ZN(n540) );
  NAND2_X1 U515 ( .A1(n540), .A2(n512), .ZN(n459) );
  NOR2_X1 U516 ( .A1(n510), .A2(n460), .ZN(n558) );
  NAND2_X1 U517 ( .A1(n558), .A2(n461), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT55), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n463), .A2(n522), .ZN(n464) );
  XNOR2_X1 U520 ( .A(KEYINPUT119), .B(n464), .ZN(n556) );
  XNOR2_X1 U521 ( .A(n544), .B(KEYINPUT98), .ZN(n529) );
  NAND2_X1 U522 ( .A1(n556), .A2(n529), .ZN(n467) );
  XOR2_X1 U523 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(G176GAT), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n467), .B(n466), .ZN(G1349GAT) );
  NAND2_X1 U526 ( .A1(n556), .A2(n550), .ZN(n471) );
  XOR2_X1 U527 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n469) );
  XNOR2_X1 U528 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n468) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n480) );
  XNOR2_X1 U530 ( .A(KEYINPUT16), .B(KEYINPUT75), .ZN(n474) );
  INV_X1 U531 ( .A(n570), .ZN(n472) );
  NOR2_X1 U532 ( .A1(n550), .A2(n472), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n476) );
  NOR2_X1 U534 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U535 ( .A(KEYINPUT95), .B(n477), .ZN(n494) );
  NOR2_X1 U536 ( .A1(n478), .A2(n494), .ZN(n486) );
  NAND2_X1 U537 ( .A1(n510), .A2(n486), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(G1324GAT) );
  NAND2_X1 U539 ( .A1(n486), .A2(n512), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT96), .ZN(n482) );
  XNOR2_X1 U541 ( .A(G8GAT), .B(n482), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U543 ( .A1(n486), .A2(n522), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  INV_X1 U545 ( .A(n485), .ZN(n516) );
  NAND2_X1 U546 ( .A1(n516), .A2(n486), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n487), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .Z(n489) );
  NAND2_X1 U549 ( .A1(n510), .A2(n491), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  NAND2_X1 U551 ( .A1(n491), .A2(n512), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n490), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U553 ( .A1(n491), .A2(n516), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n492), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT99), .B(KEYINPUT42), .Z(n496) );
  INV_X1 U556 ( .A(n561), .ZN(n493) );
  NAND2_X1 U557 ( .A1(n493), .A2(n529), .ZN(n508) );
  NOR2_X1 U558 ( .A1(n494), .A2(n508), .ZN(n503) );
  NAND2_X1 U559 ( .A1(n503), .A2(n510), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(n497), .ZN(G1332GAT) );
  NAND2_X1 U562 ( .A1(n503), .A2(n512), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n498), .B(KEYINPUT100), .ZN(n499) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(n499), .ZN(G1333GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n501) );
  NAND2_X1 U566 ( .A1(n503), .A2(n522), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G71GAT), .B(n502), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT43), .B(KEYINPUT104), .Z(n505) );
  NAND2_X1 U570 ( .A1(n503), .A2(n516), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(n507) );
  XOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT103), .Z(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  NOR2_X1 U574 ( .A1(n509), .A2(n508), .ZN(n517) );
  NAND2_X1 U575 ( .A1(n510), .A2(n517), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U577 ( .A1(n517), .A2(n512), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U579 ( .A(G99GAT), .B(KEYINPUT105), .Z(n515) );
  NAND2_X1 U580 ( .A1(n517), .A2(n522), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(G1338GAT) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(KEYINPUT106), .ZN(n521) );
  XOR2_X1 U583 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n519) );
  NAND2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1339GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n527) );
  NAND2_X1 U588 ( .A1(n540), .A2(n522), .ZN(n523) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n536) );
  INV_X1 U590 ( .A(n525), .ZN(n553) );
  NAND2_X1 U591 ( .A1(n536), .A2(n553), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n531) );
  NAND2_X1 U595 ( .A1(n536), .A2(n529), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(n532), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n534) );
  NAND2_X1 U599 ( .A1(n536), .A2(n570), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U603 ( .A1(n536), .A2(n550), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U606 ( .A1(n559), .A2(n541), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n561), .A2(n551), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(KEYINPUT116), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n546) );
  NAND2_X1 U611 ( .A1(n551), .A2(n544), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT117), .Z(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n570), .A2(n551), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U619 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n556), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1348GAT) );
  NAND2_X1 U622 ( .A1(n570), .A2(n556), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U624 ( .A(n558), .ZN(n560) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n574) );
  AND2_X1 U626 ( .A1(n561), .A2(n574), .ZN(n563) );
  XNOR2_X1 U627 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U629 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1352GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n568) );
  NAND2_X1 U632 ( .A1(n574), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G204GAT), .B(n569), .ZN(G1353GAT) );
  XOR2_X1 U635 ( .A(G211GAT), .B(KEYINPUT125), .Z(n572) );
  NAND2_X1 U636 ( .A1(n574), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1354GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n576) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(G218GAT), .B(n577), .Z(G1355GAT) );
endmodule

