//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n574, new_n575, new_n576, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204, new_n1205, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n457), .B2(new_n458), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n463), .A2(new_n465), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n473), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n466), .A2(new_n473), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(G124), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT68), .ZN(G162));
  NAND4_X1  g060(.A1(new_n473), .A2(KEYINPUT70), .A3(KEYINPUT4), .A4(G138), .ZN(new_n486));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(new_n473), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(new_n479), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n473), .ZN(new_n490));
  XOR2_X1   g065(.A(KEYINPUT70), .B(KEYINPUT4), .Z(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(KEYINPUT69), .A2(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT69), .A2(G114), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n493), .A2(G2105), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n489), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  AND3_X1   g076(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n502));
  AOI21_X1  g077(.A(G543), .B1(KEYINPUT72), .B2(KEYINPUT5), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G62), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n502), .A2(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n506), .A2(G651), .B1(new_n510), .B2(G88), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT71), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR3_X1    g090(.A1(new_n513), .A2(KEYINPUT71), .A3(new_n514), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n511), .A2(new_n515), .A3(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(new_n512), .A2(G51), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  NAND3_X1  g098(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n523), .B1(new_n522), .B2(new_n524), .ZN(new_n527));
  OAI211_X1 g102(.A(G63), .B(G651), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n532), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n529), .B(new_n534), .C1(new_n509), .C2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n522), .A2(new_n524), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n538), .A2(G89), .A3(new_n512), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n529), .B1(new_n539), .B2(new_n534), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n519), .B(new_n528), .C1(new_n537), .C2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(KEYINPUT75), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n543));
  INV_X1    g118(.A(new_n519), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n534), .B1(new_n509), .B2(new_n535), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n544), .B1(new_n546), .B2(new_n536), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n543), .B1(new_n547), .B2(new_n528), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n542), .A2(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n513), .A2(new_n551), .B1(new_n509), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n538), .A2(KEYINPUT73), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(new_n525), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G64), .ZN(new_n556));
  NAND2_X1  g131(.A1(G77), .A2(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n553), .B1(new_n558), .B2(G651), .ZN(G171));
  INV_X1    g134(.A(G651), .ZN(new_n560));
  OAI21_X1  g135(.A(G56), .B1(new_n526), .B2(new_n527), .ZN(new_n561));
  INV_X1    g136(.A(G68), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(new_n521), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n560), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G43), .ZN(new_n566));
  INV_X1    g141(.A(G81), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n513), .A2(new_n566), .B1(new_n509), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT76), .Z(G153));
  AND3_X1   g146(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G36), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT77), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT8), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n572), .A2(new_n576), .ZN(G188));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n504), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n538), .A2(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G65), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n510), .A2(G91), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n512), .A2(G53), .A3(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT9), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(G299));
  INV_X1    g164(.A(G171), .ZN(G301));
  OAI21_X1  g165(.A(G651), .B1(new_n555), .B2(G74), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n512), .A2(G543), .ZN(new_n594));
  AOI22_X1  g169(.A1(G49), .A2(new_n594), .B1(new_n510), .B2(G87), .ZN(new_n595));
  OAI211_X1 g170(.A(KEYINPUT79), .B(G651), .C1(new_n555), .C2(G74), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(G288));
  NAND2_X1  g172(.A1(new_n594), .A2(G48), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n538), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n560), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(G86), .B2(new_n510), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n600), .A2(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(new_n555), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(new_n560), .ZN(new_n606));
  AOI22_X1  g181(.A1(G47), .A2(new_n594), .B1(new_n510), .B2(G85), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n510), .A2(G92), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT10), .Z(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n582), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(G54), .B2(new_n594), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n609), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(G868), .B2(new_n620), .ZN(G297));
  XNOR2_X1  g196(.A(G297), .B(KEYINPUT81), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g203(.A(new_n480), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G2104), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT82), .B(G2100), .Z(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT84), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n634), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT83), .Z(new_n638));
  AOI22_X1  g213(.A1(new_n629), .A2(G135), .B1(G123), .B2(new_n483), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(KEYINPUT85), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(KEYINPUT85), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n641), .B(new_n642), .C1(G111), .C2(new_n473), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT86), .B(G2096), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n636), .A2(new_n638), .A3(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2435), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2438), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(KEYINPUT87), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(KEYINPUT87), .ZN(new_n662));
  NAND4_X1  g237(.A1(new_n660), .A2(G14), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT88), .Z(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2067), .B(G2678), .Z(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2096), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT17), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n667), .B2(new_n668), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n670), .B1(new_n669), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n673), .B(new_n676), .Z(G227));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n679), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n681), .A2(new_n683), .A3(new_n685), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n688), .B(new_n689), .C1(new_n687), .C2(new_n686), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n690), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT90), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n600), .B2(new_n603), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(G6), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n703), .A2(new_n701), .A3(new_n704), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n700), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n707), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n709), .A2(new_n699), .A3(new_n705), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n702), .A2(G23), .ZN(new_n712));
  INV_X1    g287(.A(G288), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n702), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT92), .B(KEYINPUT33), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1976), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n717), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n702), .A2(G22), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G166), .B2(new_n702), .ZN(new_n722));
  INV_X1    g297(.A(G1971), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n711), .A2(KEYINPUT34), .A3(new_n720), .A4(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT34), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n708), .A2(new_n710), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n718), .A2(new_n724), .A3(new_n719), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n702), .A2(G24), .ZN(new_n731));
  INV_X1    g306(.A(G290), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n702), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(G1986), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(G1986), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n483), .A2(G119), .ZN(new_n736));
  INV_X1    g311(.A(G131), .ZN(new_n737));
  NOR2_X1   g312(.A1(G95), .A2(G2105), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(new_n473), .B2(G107), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n736), .B1(new_n480), .B2(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  MUX2_X1   g315(.A(G25), .B(new_n740), .S(G29), .Z(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT35), .B(G1991), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n741), .B(new_n742), .Z(new_n743));
  NAND3_X1  g318(.A1(new_n734), .A2(new_n735), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n730), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT94), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(KEYINPUT93), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT94), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n730), .A2(new_n750), .A3(new_n745), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n747), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G2090), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n754));
  NAND2_X1  g329(.A1(G162), .A2(G29), .ZN(new_n755));
  NOR2_X1   g330(.A1(G29), .A2(G35), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n754), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  AOI211_X1 g333(.A(KEYINPUT29), .B(new_n756), .C1(G162), .C2(G29), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n753), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT98), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  NAND2_X1  g337(.A1(G164), .A2(G29), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G27), .B2(G29), .ZN(new_n764));
  INV_X1    g339(.A(G2078), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(G28), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(G28), .ZN(new_n769));
  INV_X1    g344(.A(G29), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n766), .B(new_n771), .C1(new_n765), .C2(new_n764), .ZN(new_n772));
  OR2_X1    g347(.A1(G29), .A2(G33), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n629), .A2(G139), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT25), .Z(new_n776));
  AOI22_X1  g351(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT97), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n774), .B(new_n776), .C1(new_n778), .C2(new_n473), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n773), .B1(new_n779), .B2(new_n770), .ZN(new_n780));
  INV_X1    g355(.A(G2072), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n644), .A2(new_n770), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n772), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n483), .A2(G128), .ZN(new_n785));
  INV_X1    g360(.A(G140), .ZN(new_n786));
  NOR2_X1   g361(.A1(G104), .A2(G2105), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(new_n473), .B2(G116), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n785), .B1(new_n480), .B2(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G29), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n770), .A2(G26), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT96), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT28), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G2067), .ZN(new_n795));
  NOR2_X1   g370(.A1(G29), .A2(G32), .ZN(new_n796));
  NAND2_X1  g371(.A1(G105), .A2(G2104), .ZN(new_n797));
  INV_X1    g372(.A(G141), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n466), .B2(new_n798), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n799), .A2(new_n473), .B1(new_n483), .B2(G129), .ZN(new_n800));
  NAND3_X1  g375(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT26), .Z(new_n802));
  AND2_X1   g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT27), .B(G1996), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n795), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G19), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT95), .B1(new_n808), .B2(G16), .ZN(new_n809));
  OR3_X1    g384(.A1(new_n808), .A2(KEYINPUT95), .A3(G16), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n809), .B(new_n810), .C1(new_n569), .C2(new_n702), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1341), .Z(new_n812));
  NAND4_X1  g387(.A1(new_n761), .A2(new_n784), .A3(new_n807), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n702), .A2(G5), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G171), .B2(new_n702), .ZN(new_n815));
  INV_X1    g390(.A(G1961), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(G4), .A2(G16), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n616), .B2(G16), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n817), .B1(G1348), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n819), .A2(G1348), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n780), .A2(new_n781), .ZN(new_n822));
  AND2_X1   g397(.A1(KEYINPUT24), .A2(G34), .ZN(new_n823));
  NOR2_X1   g398(.A1(KEYINPUT24), .A2(G34), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n770), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n475), .B2(new_n770), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G2084), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  NOR4_X1   g403(.A1(new_n813), .A2(new_n820), .A3(new_n821), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n750), .B1(new_n730), .B2(new_n745), .ZN(new_n830));
  AOI211_X1 g405(.A(KEYINPUT94), .B(new_n744), .C1(new_n725), .C2(new_n729), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n830), .A2(new_n831), .B1(KEYINPUT93), .B2(new_n748), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n702), .A2(KEYINPUT23), .A3(G20), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT23), .ZN(new_n834));
  INV_X1    g409(.A(G20), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(G16), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n836), .C1(new_n620), .C2(new_n702), .ZN(new_n837));
  INV_X1    g412(.A(G1956), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n752), .A2(new_n829), .A3(new_n832), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n758), .A2(new_n759), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G2090), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(G168), .A2(G16), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(G16), .B2(G21), .ZN(new_n845));
  INV_X1    g420(.A(G1966), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n840), .A2(new_n843), .A3(new_n847), .ZN(G311));
  AND3_X1   g423(.A1(new_n829), .A2(new_n752), .A3(new_n832), .ZN(new_n849));
  INV_X1    g424(.A(new_n847), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n849), .A2(new_n842), .A3(new_n850), .A4(new_n839), .ZN(G150));
  OAI21_X1  g426(.A(G67), .B1(new_n526), .B2(new_n527), .ZN(new_n852));
  INV_X1    g427(.A(G80), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(new_n521), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n560), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(G55), .ZN(new_n857));
  INV_X1    g432(.A(G93), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n513), .A2(new_n857), .B1(new_n509), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(G860), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  INV_X1    g436(.A(G56), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n554), .B2(new_n525), .ZN(new_n863));
  OAI21_X1  g438(.A(G651), .B1(new_n863), .B2(new_n563), .ZN(new_n864));
  INV_X1    g439(.A(new_n568), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n864), .B(new_n865), .C1(new_n856), .C2(new_n859), .ZN(new_n866));
  INV_X1    g441(.A(G67), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n554), .B2(new_n525), .ZN(new_n868));
  OAI21_X1  g443(.A(G651), .B1(new_n868), .B2(new_n854), .ZN(new_n869));
  INV_X1    g444(.A(new_n859), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n869), .B(new_n870), .C1(new_n565), .C2(new_n568), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n611), .A2(new_n615), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(new_n623), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n874), .B(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n861), .B1(new_n877), .B2(G860), .ZN(G145));
  XNOR2_X1  g453(.A(new_n779), .B(new_n499), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n631), .B(new_n789), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n483), .A2(G130), .ZN(new_n882));
  INV_X1    g457(.A(G142), .ZN(new_n883));
  NOR2_X1   g458(.A1(G106), .A2(G2105), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n885));
  OAI221_X1 g460(.A(new_n882), .B1(new_n480), .B2(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n740), .B(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n881), .A2(new_n887), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n644), .B(new_n475), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(G162), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n803), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n890), .B(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g472(.A(new_n872), .B(KEYINPUT99), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n625), .ZN(new_n899));
  XOR2_X1   g474(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n900));
  NOR2_X1   g475(.A1(new_n875), .A2(G299), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n584), .A2(G651), .B1(G91), .B2(new_n510), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n615), .A2(new_n611), .B1(new_n902), .B2(new_n588), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n900), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n875), .B(G299), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n904), .B1(new_n905), .B2(KEYINPUT41), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n899), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n901), .A2(new_n903), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n908), .B1(new_n909), .B2(new_n899), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n911));
  NAND2_X1  g486(.A1(G290), .A2(G166), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n606), .A2(G303), .A3(new_n607), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(G288), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(G288), .B1(new_n912), .B2(new_n913), .ZN(new_n916));
  OAI21_X1  g491(.A(G305), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  INV_X1    g493(.A(G305), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n911), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n911), .B2(new_n923), .ZN(new_n925));
  OAI21_X1  g500(.A(G868), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n856), .A2(new_n859), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n926), .B1(G868), .B2(new_n927), .ZN(G295));
  OAI21_X1  g503(.A(new_n926), .B1(G868), .B2(new_n927), .ZN(G331));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n541), .A2(KEYINPUT75), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n546), .A2(new_n536), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(new_n543), .A3(new_n519), .A4(new_n528), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n932), .A2(new_n934), .A3(G171), .ZN(new_n935));
  AOI21_X1  g510(.A(G171), .B1(new_n932), .B2(new_n934), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n935), .A2(new_n936), .A3(new_n872), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n866), .A2(new_n871), .ZN(new_n938));
  OAI21_X1  g513(.A(G301), .B1(new_n542), .B2(new_n548), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n932), .A2(G171), .A3(new_n934), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n931), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n872), .B1(new_n935), .B2(new_n936), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT101), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n909), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n906), .B1(new_n937), .B2(new_n941), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n921), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n895), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n921), .B1(new_n945), .B2(new_n946), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n930), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n905), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n909), .A2(new_n900), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n939), .A2(new_n938), .A3(new_n940), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT101), .B1(new_n943), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n939), .A2(new_n940), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n931), .B1(new_n956), .B2(new_n872), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n952), .B(new_n953), .C1(new_n955), .C2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n943), .A2(new_n954), .A3(new_n909), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n922), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n961), .A2(KEYINPUT43), .A3(new_n895), .A4(new_n947), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n950), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT44), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n909), .A2(new_n951), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n966), .A2(new_n904), .B1(new_n954), .B2(new_n943), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n955), .A2(new_n957), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(new_n909), .ZN(new_n969));
  AOI21_X1  g544(.A(G37), .B1(new_n969), .B2(new_n921), .ZN(new_n970));
  INV_X1    g545(.A(new_n949), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n930), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n921), .B1(new_n958), .B2(new_n959), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n948), .A2(KEYINPUT43), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n965), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT102), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n964), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n965), .B1(new_n950), .B2(new_n962), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT43), .B1(new_n948), .B2(new_n949), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n961), .A2(new_n930), .A3(new_n895), .A4(new_n947), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT44), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT102), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n977), .A2(new_n982), .ZN(G397));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n499), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT103), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n488), .A2(new_n479), .B1(new_n495), .B2(new_n497), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n988), .B2(new_n492), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT103), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT104), .B(G40), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n469), .A2(new_n474), .A3(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  OR3_X1    g570(.A1(new_n995), .A2(G1986), .A3(G290), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n996), .B(KEYINPUT127), .Z(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT48), .ZN(new_n998));
  INV_X1    g573(.A(G2067), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n789), .B(new_n999), .ZN(new_n1000));
  OR3_X1    g575(.A1(new_n995), .A2(KEYINPUT106), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT106), .B1(new_n995), .B2(new_n1000), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n803), .B(G1996), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1001), .B(new_n1002), .C1(new_n995), .C2(new_n1003), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n740), .A2(new_n742), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n740), .A2(new_n742), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n995), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n998), .A2(new_n1008), .ZN(new_n1009));
  OAI22_X1  g584(.A1(new_n1004), .A2(new_n1005), .B1(G2067), .B2(new_n789), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n992), .A2(new_n994), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n995), .B1(new_n803), .B2(new_n1000), .ZN(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1011), .A2(KEYINPUT46), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT46), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT126), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT47), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1009), .A2(new_n1012), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n985), .A2(new_n994), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT49), .ZN(new_n1026));
  INV_X1    g601(.A(G1981), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n600), .A2(new_n1027), .A3(new_n603), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n600), .B2(new_n603), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1025), .A2(KEYINPUT49), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1024), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1034));
  AOI211_X1 g609(.A(G1976), .B(G288), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1035), .A2(new_n1028), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n994), .B1(new_n985), .B2(new_n991), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n723), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n989), .A2(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n469), .A2(new_n474), .A3(new_n993), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1040), .B1(G2090), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT109), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G303), .A2(G8), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT55), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT109), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1040), .B(new_n1052), .C1(G2090), .C2(new_n1046), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1048), .A2(G8), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1976), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1023), .B1(G288), .B2(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  OR3_X1    g634(.A1(new_n713), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1059), .A2(new_n1060), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1036), .A2(new_n1023), .B1(new_n1055), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1048), .A2(G8), .A3(new_n1053), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1050), .A2(KEYINPUT116), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1064), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(new_n994), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1045), .B(KEYINPUT113), .C1(KEYINPUT45), .C2(new_n989), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1038), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n846), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT114), .B(G2084), .Z(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1046), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n994), .B1(new_n989), .B2(new_n1043), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1076), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(KEYINPUT115), .A3(new_n1041), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1074), .A2(new_n1081), .A3(G168), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G8), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G286), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1068), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1048), .A2(G8), .A3(new_n1066), .A4(new_n1053), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1061), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1063), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1061), .A2(new_n1086), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(KEYINPUT117), .A3(new_n1084), .A4(new_n1068), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1045), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n989), .A2(new_n1043), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1040), .B1(new_n1094), .B2(G2090), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1095), .A2(KEYINPUT112), .ZN(new_n1096));
  OAI21_X1  g671(.A(G8), .B1(new_n1095), .B2(KEYINPUT112), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1050), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(new_n1061), .A3(new_n1054), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT63), .B1(new_n1100), .B2(new_n1084), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1062), .B1(new_n1091), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n902), .B2(new_n588), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n838), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1037), .A2(new_n1038), .A3(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1112));
  NAND2_X1  g687(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n902), .A2(new_n1104), .A3(new_n588), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT119), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT61), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1111), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT120), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1111), .A2(new_n1116), .A3(new_n1118), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G1348), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1046), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1021), .A2(new_n999), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(KEYINPUT60), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n616), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT122), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1130), .A3(new_n616), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT121), .B1(new_n1127), .B2(new_n616), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1046), .A2(new_n1124), .B1(new_n999), .B2(new_n1021), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1134), .A2(new_n1135), .A3(KEYINPUT60), .A4(new_n875), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1132), .A2(new_n1137), .B1(KEYINPUT60), .B2(new_n1134), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1117), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1037), .A2(new_n1014), .A3(new_n1038), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1045), .A2(new_n989), .ZN(new_n1144));
  XOR2_X1   g719(.A(KEYINPUT58), .B(G1341), .Z(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1142), .B1(new_n1147), .B2(new_n569), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n569), .ZN(new_n1150));
  AOI211_X1 g725(.A(KEYINPUT118), .B(new_n1150), .C1(new_n1143), .C2(new_n1146), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT59), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1148), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1123), .A2(new_n1138), .A3(new_n1141), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1139), .ZN(new_n1158));
  OR3_X1    g733(.A1(new_n1140), .A2(new_n875), .A3(new_n1134), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  XOR2_X1   g735(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1161));
  NAND3_X1  g736(.A1(new_n1037), .A2(new_n765), .A3(new_n1038), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1162), .A2(new_n1163), .B1(new_n816), .B2(new_n1046), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n765), .A2(KEYINPUT53), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1073), .B2(new_n1165), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1166), .A2(G171), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n474), .A2(KEYINPUT125), .B1(G2105), .B2(new_n468), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n474), .A2(KEYINPUT125), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1169), .A2(G40), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n992), .A2(new_n1038), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1164), .B(G301), .C1(new_n1165), .C2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1161), .B1(new_n1167), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1164), .B1(new_n1171), .B2(new_n1165), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(G171), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1176), .B(KEYINPUT54), .C1(G171), .C2(new_n1166), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1179));
  AOI21_X1  g754(.A(G168), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT51), .ZN(new_n1181));
  OAI211_X1 g756(.A(G8), .B(new_n1082), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(KEYINPUT123), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1179), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1178), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1160), .A2(new_n1187), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1179), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1185), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1190));
  OAI21_X1  g765(.A(KEYINPUT62), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1184), .A2(new_n1192), .A3(new_n1186), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1191), .A2(new_n1193), .A3(new_n1167), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1188), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1102), .B1(new_n1195), .B2(new_n1100), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1011), .A2(G1986), .A3(G290), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n996), .A2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT105), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1199), .A2(new_n1008), .ZN(new_n1200));
  XOR2_X1   g775(.A(new_n1200), .B(KEYINPUT107), .Z(new_n1201));
  OAI21_X1  g776(.A(new_n1020), .B1(new_n1196), .B2(new_n1201), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g777(.A(G227), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n663), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g779(.A(new_n1205), .B1(new_n894), .B2(new_n895), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n980), .ZN(new_n1207));
  NAND4_X1  g781(.A1(new_n1206), .A2(G319), .A3(new_n697), .A4(new_n1207), .ZN(G225));
  INV_X1    g782(.A(G225), .ZN(G308));
endmodule


