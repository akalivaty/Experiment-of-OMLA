

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751;

  XNOR2_X1 U385 ( .A(n578), .B(KEYINPUT1), .ZN(n500) );
  INV_X2 U386 ( .A(G953), .ZN(n744) );
  NOR2_X2 U387 ( .A1(n598), .A2(n597), .ZN(n599) );
  AND2_X2 U388 ( .A1(n602), .A2(n629), .ZN(n441) );
  XNOR2_X2 U389 ( .A(n439), .B(n723), .ZN(n629) );
  XNOR2_X2 U390 ( .A(n399), .B(G104), .ZN(n432) );
  XNOR2_X2 U391 ( .A(G143), .B(G128), .ZN(n425) );
  AND2_X1 U392 ( .A1(n612), .A2(n697), .ZN(n704) );
  INV_X1 U393 ( .A(n501), .ZN(n670) );
  AND2_X1 U394 ( .A1(n618), .A2(n617), .ZN(n620) );
  NOR2_X1 U395 ( .A1(n699), .A2(n610), .ZN(n611) );
  BUF_X1 U396 ( .A(n699), .Z(n700) );
  AND2_X1 U397 ( .A1(n527), .A2(n526), .ZN(n538) );
  AND2_X1 U398 ( .A1(n550), .A2(n510), .ZN(n503) );
  XNOR2_X1 U399 ( .A(n377), .B(n376), .ZN(n667) );
  XNOR2_X1 U400 ( .A(n433), .B(KEYINPUT73), .ZN(n434) );
  XNOR2_X1 U401 ( .A(G122), .B(KEYINPUT16), .ZN(n433) );
  NOR2_X2 U402 ( .A1(n748), .A2(KEYINPUT44), .ZN(n507) );
  XNOR2_X1 U403 ( .A(n364), .B(n607), .ZN(n613) );
  INV_X1 U404 ( .A(KEYINPUT64), .ZN(n364) );
  XNOR2_X2 U405 ( .A(n539), .B(KEYINPUT45), .ZN(n727) );
  INV_X1 U406 ( .A(n454), .ZN(n372) );
  NOR2_X1 U407 ( .A1(n670), .A2(n543), .ZN(n545) );
  INV_X1 U408 ( .A(n667), .ZN(n550) );
  AND2_X1 U409 ( .A1(n667), .A2(n666), .ZN(n664) );
  XNOR2_X1 U410 ( .A(n367), .B(G125), .ZN(n428) );
  INV_X1 U411 ( .A(G146), .ZN(n367) );
  AND2_X1 U412 ( .A1(n371), .A2(n574), .ZN(n370) );
  NAND2_X1 U413 ( .A1(n373), .A2(n372), .ZN(n371) );
  XNOR2_X1 U414 ( .A(n464), .B(n397), .ZN(n409) );
  NAND2_X1 U415 ( .A1(n664), .A2(n663), .ZN(n517) );
  NOR2_X1 U416 ( .A1(n552), .A2(n551), .ZN(n566) );
  XNOR2_X1 U417 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U418 ( .A(n428), .B(n366), .ZN(n737) );
  XNOR2_X1 U419 ( .A(KEYINPUT10), .B(G140), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n425), .B(G134), .ZN(n464) );
  XNOR2_X1 U421 ( .A(n409), .B(n398), .ZN(n738) );
  NOR2_X1 U422 ( .A1(n552), .A2(n546), .ZN(n548) );
  XNOR2_X1 U423 ( .A(n545), .B(n544), .ZN(n546) );
  INV_X1 U424 ( .A(KEYINPUT30), .ZN(n544) );
  XNOR2_X1 U425 ( .A(n392), .B(n393), .ZN(n376) );
  OR2_X1 U426 ( .A1(n720), .A2(G902), .ZN(n377) );
  XNOR2_X1 U427 ( .A(n431), .B(n430), .ZN(n439) );
  AND2_X1 U428 ( .A1(n616), .A2(G953), .ZN(n722) );
  OR2_X1 U429 ( .A1(n580), .A2(n578), .ZN(n569) );
  XNOR2_X1 U430 ( .A(n563), .B(n562), .ZN(n750) );
  NAND2_X1 U431 ( .A1(n365), .A2(n368), .ZN(n488) );
  XOR2_X1 U432 ( .A(n581), .B(KEYINPUT78), .Z(n650) );
  OR2_X1 U433 ( .A1(n580), .A2(n380), .ZN(n581) );
  AND2_X1 U434 ( .A1(n374), .A2(n370), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n549), .B(KEYINPUT39), .ZN(n561) );
  NAND2_X1 U436 ( .A1(n369), .A2(n372), .ZN(n368) );
  INV_X1 U437 ( .A(n709), .ZN(n369) );
  INV_X1 U438 ( .A(n493), .ZN(n373) );
  NAND2_X1 U439 ( .A1(n709), .A2(n375), .ZN(n374) );
  AND2_X1 U440 ( .A1(n493), .A2(n454), .ZN(n375) );
  XNOR2_X2 U441 ( .A(n421), .B(n420), .ZN(n709) );
  XNOR2_X1 U442 ( .A(KEYINPUT62), .B(n614), .ZN(n378) );
  XOR2_X1 U443 ( .A(n412), .B(n436), .Z(n379) );
  OR2_X1 U444 ( .A1(n579), .A2(n578), .ZN(n380) );
  AND2_X1 U445 ( .A1(n577), .A2(n590), .ZN(n582) );
  INV_X1 U446 ( .A(KEYINPUT75), .ZN(n406) );
  XNOR2_X1 U447 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U448 ( .A(n409), .B(n408), .ZN(n415) );
  INV_X1 U449 ( .A(n436), .ZN(n437) );
  BUF_X1 U450 ( .A(n727), .Z(n697) );
  XNOR2_X1 U451 ( .A(KEYINPUT38), .B(n557), .ZN(n680) );
  XNOR2_X1 U452 ( .A(n496), .B(n495), .ZN(n510) );
  XNOR2_X1 U453 ( .A(n737), .B(n385), .ZN(n390) );
  BUF_X1 U454 ( .A(n714), .Z(n718) );
  AND2_X1 U455 ( .A1(n548), .A2(n547), .ZN(n573) );
  INV_X1 U456 ( .A(n722), .ZN(n617) );
  XNOR2_X1 U457 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n570) );
  XNOR2_X1 U458 ( .A(n571), .B(n570), .ZN(n751) );
  XOR2_X1 U459 ( .A(KEYINPUT23), .B(G110), .Z(n382) );
  XNOR2_X1 U460 ( .A(G128), .B(G119), .ZN(n381) );
  XNOR2_X1 U461 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U462 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n383) );
  XNOR2_X1 U463 ( .A(KEYINPUT68), .B(G137), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n398), .B(KEYINPUT76), .ZN(n388) );
  NAND2_X1 U465 ( .A1(G234), .A2(n744), .ZN(n386) );
  XOR2_X1 U466 ( .A(KEYINPUT8), .B(n386), .Z(n461) );
  NAND2_X1 U467 ( .A1(G221), .A2(n461), .ZN(n387) );
  XNOR2_X1 U468 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U469 ( .A(n390), .B(n389), .ZN(n720) );
  XNOR2_X1 U470 ( .A(G902), .B(KEYINPUT15), .ZN(n602) );
  NAND2_X1 U471 ( .A1(G234), .A2(n602), .ZN(n391) );
  XNOR2_X1 U472 ( .A(KEYINPUT20), .B(n391), .ZN(n394) );
  NAND2_X1 U473 ( .A1(G217), .A2(n394), .ZN(n392) );
  INV_X1 U474 ( .A(KEYINPUT25), .ZN(n393) );
  NAND2_X1 U475 ( .A1(n394), .A2(G221), .ZN(n396) );
  INV_X1 U476 ( .A(KEYINPUT21), .ZN(n395) );
  XNOR2_X1 U477 ( .A(n396), .B(n395), .ZN(n666) );
  XNOR2_X1 U478 ( .A(KEYINPUT4), .B(G131), .ZN(n397) );
  XNOR2_X2 U479 ( .A(G110), .B(G107), .ZN(n399) );
  NAND2_X1 U480 ( .A1(n744), .A2(G227), .ZN(n400) );
  XNOR2_X1 U481 ( .A(n400), .B(G140), .ZN(n401) );
  XNOR2_X1 U482 ( .A(n432), .B(n401), .ZN(n402) );
  XNOR2_X2 U483 ( .A(KEYINPUT67), .B(G101), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n429), .B(G146), .ZN(n412) );
  XNOR2_X1 U485 ( .A(n402), .B(n412), .ZN(n403) );
  XNOR2_X1 U486 ( .A(n738), .B(n403), .ZN(n635) );
  OR2_X2 U487 ( .A1(n635), .A2(G902), .ZN(n405) );
  XNOR2_X1 U488 ( .A(KEYINPUT69), .B(G469), .ZN(n404) );
  XNOR2_X2 U489 ( .A(n405), .B(n404), .ZN(n578) );
  INV_X1 U490 ( .A(n500), .ZN(n663) );
  XNOR2_X1 U491 ( .A(n517), .B(KEYINPUT105), .ZN(n418) );
  XNOR2_X1 U492 ( .A(G137), .B(KEYINPUT5), .ZN(n407) );
  XOR2_X1 U493 ( .A(G113), .B(G116), .Z(n411) );
  XNOR2_X1 U494 ( .A(KEYINPUT3), .B(G119), .ZN(n410) );
  XNOR2_X1 U495 ( .A(n411), .B(n410), .ZN(n436) );
  NOR2_X1 U496 ( .A1(G953), .A2(G237), .ZN(n473) );
  NAND2_X1 U497 ( .A1(n473), .A2(G210), .ZN(n413) );
  XNOR2_X1 U498 ( .A(n379), .B(n413), .ZN(n414) );
  XNOR2_X1 U499 ( .A(n415), .B(n414), .ZN(n614) );
  INV_X1 U500 ( .A(G902), .ZN(n482) );
  NAND2_X1 U501 ( .A1(n614), .A2(n482), .ZN(n416) );
  XNOR2_X2 U502 ( .A(n416), .B(G472), .ZN(n501) );
  XNOR2_X1 U503 ( .A(n501), .B(KEYINPUT6), .ZN(n553) );
  INV_X1 U504 ( .A(n553), .ZN(n417) );
  NAND2_X1 U505 ( .A1(n418), .A2(n417), .ZN(n421) );
  INV_X1 U506 ( .A(KEYINPUT87), .ZN(n419) );
  XNOR2_X1 U507 ( .A(n419), .B(KEYINPUT33), .ZN(n420) );
  XOR2_X1 U508 ( .A(KEYINPUT88), .B(KEYINPUT17), .Z(n423) );
  XNOR2_X1 U509 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n422) );
  XNOR2_X1 U510 ( .A(n423), .B(n422), .ZN(n427) );
  NAND2_X1 U511 ( .A1(G224), .A2(n744), .ZN(n424) );
  XNOR2_X1 U512 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U513 ( .A(n427), .B(n426), .ZN(n431) );
  XNOR2_X1 U514 ( .A(n429), .B(n428), .ZN(n430) );
  INV_X1 U515 ( .A(n432), .ZN(n435) );
  XNOR2_X2 U516 ( .A(n435), .B(n434), .ZN(n438) );
  XNOR2_X2 U517 ( .A(n438), .B(n437), .ZN(n723) );
  OR2_X1 U518 ( .A1(G237), .A2(G902), .ZN(n442) );
  NAND2_X1 U519 ( .A1(n442), .A2(G210), .ZN(n440) );
  XNOR2_X2 U520 ( .A(n441), .B(n440), .ZN(n576) );
  NAND2_X1 U521 ( .A1(G214), .A2(n442), .ZN(n443) );
  XOR2_X1 U522 ( .A(KEYINPUT89), .B(n443), .Z(n679) );
  AND2_X2 U523 ( .A1(n576), .A2(n679), .ZN(n584) );
  XNOR2_X1 U524 ( .A(n584), .B(KEYINPUT19), .ZN(n579) );
  NAND2_X1 U525 ( .A1(G234), .A2(G237), .ZN(n444) );
  XNOR2_X1 U526 ( .A(n444), .B(KEYINPUT14), .ZN(n445) );
  XNOR2_X1 U527 ( .A(KEYINPUT74), .B(n445), .ZN(n446) );
  NAND2_X1 U528 ( .A1(G952), .A2(n446), .ZN(n695) );
  NOR2_X1 U529 ( .A1(G953), .A2(n695), .ZN(n542) );
  NAND2_X1 U530 ( .A1(G902), .A2(n446), .ZN(n447) );
  XOR2_X1 U531 ( .A(KEYINPUT90), .B(n447), .Z(n448) );
  NAND2_X1 U532 ( .A1(G953), .A2(n448), .ZN(n540) );
  NOR2_X1 U533 ( .A1(G898), .A2(n540), .ZN(n449) );
  NOR2_X1 U534 ( .A1(n542), .A2(n449), .ZN(n450) );
  NOR2_X1 U535 ( .A1(n579), .A2(n450), .ZN(n452) );
  XNOR2_X1 U536 ( .A(KEYINPUT86), .B(KEYINPUT0), .ZN(n451) );
  XNOR2_X2 U537 ( .A(n452), .B(n451), .ZN(n493) );
  XNOR2_X1 U538 ( .A(KEYINPUT77), .B(KEYINPUT34), .ZN(n453) );
  XNOR2_X1 U539 ( .A(n453), .B(KEYINPUT70), .ZN(n454) );
  XOR2_X1 U540 ( .A(KEYINPUT100), .B(G107), .Z(n456) );
  XNOR2_X1 U541 ( .A(G116), .B(G122), .ZN(n455) );
  XNOR2_X1 U542 ( .A(n456), .B(n455), .ZN(n460) );
  XOR2_X1 U543 ( .A(KEYINPUT7), .B(KEYINPUT99), .Z(n458) );
  XNOR2_X1 U544 ( .A(KEYINPUT98), .B(KEYINPUT9), .ZN(n457) );
  XNOR2_X1 U545 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U546 ( .A(n460), .B(n459), .Z(n463) );
  NAND2_X1 U547 ( .A1(G217), .A2(n461), .ZN(n462) );
  XNOR2_X1 U548 ( .A(n463), .B(n462), .ZN(n466) );
  INV_X1 U549 ( .A(n464), .ZN(n465) );
  XNOR2_X1 U550 ( .A(n466), .B(n465), .ZN(n716) );
  NAND2_X1 U551 ( .A1(n716), .A2(n482), .ZN(n469) );
  INV_X1 U552 ( .A(KEYINPUT101), .ZN(n467) );
  XNOR2_X1 U553 ( .A(n467), .B(G478), .ZN(n468) );
  XNOR2_X1 U554 ( .A(n469), .B(n468), .ZN(n519) );
  INV_X1 U555 ( .A(n519), .ZN(n490) );
  XOR2_X1 U556 ( .A(G104), .B(G122), .Z(n471) );
  XNOR2_X1 U557 ( .A(G143), .B(G113), .ZN(n470) );
  XNOR2_X1 U558 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U559 ( .A(n737), .B(n472), .ZN(n481) );
  XOR2_X1 U560 ( .A(KEYINPUT11), .B(KEYINPUT93), .Z(n475) );
  NAND2_X1 U561 ( .A1(G214), .A2(n473), .ZN(n474) );
  XNOR2_X1 U562 ( .A(n475), .B(n474), .ZN(n479) );
  XOR2_X1 U563 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n477) );
  XNOR2_X1 U564 ( .A(G131), .B(KEYINPUT12), .ZN(n476) );
  XNOR2_X1 U565 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U566 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U567 ( .A(n481), .B(n480), .ZN(n621) );
  NAND2_X1 U568 ( .A1(n621), .A2(n482), .ZN(n486) );
  XOR2_X1 U569 ( .A(KEYINPUT97), .B(KEYINPUT13), .Z(n484) );
  XNOR2_X1 U570 ( .A(KEYINPUT96), .B(G475), .ZN(n483) );
  XNOR2_X1 U571 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U572 ( .A(n486), .B(n485), .ZN(n520) );
  NOR2_X1 U573 ( .A1(n490), .A2(n520), .ZN(n574) );
  INV_X1 U574 ( .A(KEYINPUT35), .ZN(n487) );
  XNOR2_X2 U575 ( .A(n488), .B(n487), .ZN(n531) );
  XOR2_X1 U576 ( .A(G122), .B(KEYINPUT127), .Z(n489) );
  XNOR2_X1 U577 ( .A(n531), .B(n489), .ZN(G24) );
  NAND2_X1 U578 ( .A1(n520), .A2(n490), .ZN(n682) );
  INV_X1 U579 ( .A(n666), .ZN(n491) );
  NOR2_X1 U580 ( .A1(n682), .A2(n491), .ZN(n492) );
  NAND2_X1 U581 ( .A1(n493), .A2(n492), .ZN(n496) );
  XNOR2_X1 U582 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n494) );
  XNOR2_X1 U583 ( .A(n494), .B(KEYINPUT71), .ZN(n495) );
  AND2_X1 U584 ( .A1(n553), .A2(n663), .ZN(n497) );
  NAND2_X1 U585 ( .A1(n503), .A2(n497), .ZN(n499) );
  INV_X1 U586 ( .A(KEYINPUT32), .ZN(n498) );
  XNOR2_X2 U587 ( .A(n499), .B(n498), .ZN(n748) );
  AND2_X1 U588 ( .A1(n500), .A2(n670), .ZN(n502) );
  NAND2_X1 U589 ( .A1(n503), .A2(n502), .ZN(n505) );
  INV_X1 U590 ( .A(KEYINPUT104), .ZN(n504) );
  XNOR2_X2 U591 ( .A(n505), .B(n504), .ZN(n749) );
  INV_X1 U592 ( .A(n749), .ZN(n506) );
  NAND2_X1 U593 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U594 ( .A1(n508), .A2(KEYINPUT84), .ZN(n509) );
  NAND2_X1 U595 ( .A1(n509), .A2(n531), .ZN(n527) );
  NAND2_X1 U596 ( .A1(n510), .A2(n553), .ZN(n511) );
  XNOR2_X1 U597 ( .A(KEYINPUT83), .B(n511), .ZN(n513) );
  AND2_X1 U598 ( .A1(n500), .A2(n667), .ZN(n512) );
  AND2_X1 U599 ( .A1(n513), .A2(n512), .ZN(n639) );
  INV_X1 U600 ( .A(n664), .ZN(n514) );
  NOR2_X1 U601 ( .A1(n514), .A2(n578), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n493), .A2(n547), .ZN(n515) );
  NOR2_X1 U603 ( .A1(n515), .A2(n501), .ZN(n516) );
  XNOR2_X1 U604 ( .A(n516), .B(KEYINPUT92), .ZN(n642) );
  NOR2_X1 U605 ( .A1(n517), .A2(n670), .ZN(n673) );
  NAND2_X1 U606 ( .A1(n493), .A2(n673), .ZN(n518) );
  XNOR2_X1 U607 ( .A(n518), .B(KEYINPUT31), .ZN(n657) );
  NOR2_X1 U608 ( .A1(n642), .A2(n657), .ZN(n524) );
  AND2_X1 U609 ( .A1(n519), .A2(n520), .ZN(n656) );
  NOR2_X1 U610 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U611 ( .A(n521), .B(KEYINPUT102), .ZN(n653) );
  NOR2_X1 U612 ( .A1(n656), .A2(n653), .ZN(n522) );
  XOR2_X1 U613 ( .A(KEYINPUT103), .B(n522), .Z(n685) );
  XOR2_X1 U614 ( .A(KEYINPUT79), .B(n685), .Z(n523) );
  NOR2_X1 U615 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U616 ( .A1(n639), .A2(n525), .ZN(n526) );
  INV_X1 U617 ( .A(n748), .ZN(n528) );
  NAND2_X1 U618 ( .A1(n528), .A2(KEYINPUT44), .ZN(n529) );
  NOR2_X1 U619 ( .A1(n529), .A2(n749), .ZN(n533) );
  INV_X1 U620 ( .A(KEYINPUT84), .ZN(n530) );
  OR2_X2 U621 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U622 ( .A1(n533), .A2(n532), .ZN(n536) );
  INV_X1 U623 ( .A(KEYINPUT44), .ZN(n534) );
  NAND2_X1 U624 ( .A1(n534), .A2(KEYINPUT84), .ZN(n535) );
  NAND2_X1 U625 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U626 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U627 ( .A1(G900), .A2(n540), .ZN(n541) );
  NOR2_X1 U628 ( .A1(n542), .A2(n541), .ZN(n552) );
  INV_X1 U629 ( .A(n679), .ZN(n543) );
  INV_X1 U630 ( .A(n576), .ZN(n557) );
  NAND2_X1 U631 ( .A1(n573), .A2(n680), .ZN(n549) );
  NAND2_X1 U632 ( .A1(n656), .A2(n561), .ZN(n661) );
  NAND2_X1 U633 ( .A1(n550), .A2(n666), .ZN(n551) );
  NAND2_X1 U634 ( .A1(n566), .A2(n653), .ZN(n554) );
  NOR2_X1 U635 ( .A1(n554), .A2(n553), .ZN(n585) );
  AND2_X1 U636 ( .A1(n500), .A2(n679), .ZN(n555) );
  NAND2_X1 U637 ( .A1(n585), .A2(n555), .ZN(n556) );
  XNOR2_X1 U638 ( .A(n556), .B(KEYINPUT43), .ZN(n558) );
  AND2_X1 U639 ( .A1(n558), .A2(n557), .ZN(n662) );
  INV_X1 U640 ( .A(n662), .ZN(n559) );
  AND2_X1 U641 ( .A1(n661), .A2(n559), .ZN(n608) );
  INV_X1 U642 ( .A(n608), .ZN(n560) );
  NOR2_X1 U643 ( .A1(n602), .A2(n560), .ZN(n600) );
  XOR2_X1 U644 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n563) );
  NAND2_X1 U645 ( .A1(n561), .A2(n653), .ZN(n562) );
  NAND2_X1 U646 ( .A1(n680), .A2(n679), .ZN(n684) );
  NOR2_X1 U647 ( .A1(n682), .A2(n684), .ZN(n565) );
  XNOR2_X1 U648 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n564) );
  XNOR2_X1 U649 ( .A(n565), .B(n564), .ZN(n710) );
  XOR2_X1 U650 ( .A(KEYINPUT106), .B(KEYINPUT28), .Z(n568) );
  AND2_X1 U651 ( .A1(n501), .A2(n566), .ZN(n567) );
  XNOR2_X1 U652 ( .A(n568), .B(n567), .ZN(n580) );
  NOR2_X1 U653 ( .A1(n710), .A2(n569), .ZN(n571) );
  NAND2_X1 U654 ( .A1(n750), .A2(n751), .ZN(n572) );
  XNOR2_X1 U655 ( .A(n572), .B(KEYINPUT46), .ZN(n598) );
  AND2_X1 U656 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U657 ( .A1(n576), .A2(n575), .ZN(n649) );
  NOR2_X1 U658 ( .A1(KEYINPUT79), .A2(n685), .ZN(n577) );
  INV_X1 U659 ( .A(KEYINPUT47), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n582), .A2(n650), .ZN(n583) );
  NAND2_X1 U661 ( .A1(n649), .A2(n583), .ZN(n589) );
  XOR2_X1 U662 ( .A(KEYINPUT110), .B(KEYINPUT36), .Z(n587) );
  NAND2_X1 U663 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U664 ( .A(n587), .B(n586), .Z(n588) );
  NOR2_X1 U665 ( .A1(n588), .A2(n500), .ZN(n659) );
  NOR2_X1 U666 ( .A1(n589), .A2(n659), .ZN(n596) );
  NAND2_X1 U667 ( .A1(KEYINPUT79), .A2(n650), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n594) );
  INV_X1 U669 ( .A(n685), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n592), .A2(n650), .ZN(n593) );
  NAND2_X1 U671 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n599), .B(KEYINPUT48), .ZN(n609) );
  AND2_X1 U674 ( .A1(n600), .A2(n609), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n727), .A2(n601), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n602), .B(KEYINPUT81), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n603), .A2(KEYINPUT2), .ZN(n604) );
  XOR2_X1 U678 ( .A(KEYINPUT65), .B(n604), .Z(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n699) );
  INV_X1 U681 ( .A(KEYINPUT2), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT82), .ZN(n612) );
  NOR2_X2 U683 ( .A1(n613), .A2(n704), .ZN(n714) );
  NAND2_X1 U684 ( .A1(n714), .A2(G472), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n615), .B(n378), .ZN(n618) );
  INV_X1 U686 ( .A(G952), .ZN(n616) );
  XNOR2_X1 U687 ( .A(KEYINPUT85), .B(KEYINPUT63), .ZN(n619) );
  XNOR2_X1 U688 ( .A(n620), .B(n619), .ZN(G57) );
  NAND2_X1 U689 ( .A1(n714), .A2(G475), .ZN(n623) );
  XNOR2_X1 U690 ( .A(n621), .B(KEYINPUT59), .ZN(n622) );
  XNOR2_X1 U691 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X2 U692 ( .A1(n624), .A2(n722), .ZN(n626) );
  XNOR2_X1 U693 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n625) );
  XNOR2_X1 U694 ( .A(n626), .B(n625), .ZN(G60) );
  NAND2_X1 U695 ( .A1(n714), .A2(G210), .ZN(n631) );
  XNOR2_X1 U696 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n627), .B(KEYINPUT55), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n631), .B(n630), .ZN(n632) );
  NOR2_X2 U700 ( .A1(n632), .A2(n722), .ZN(n633) );
  XNOR2_X1 U701 ( .A(n633), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U702 ( .A1(n718), .A2(G469), .ZN(n637) );
  XOR2_X1 U703 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n634) );
  XNOR2_X1 U704 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X1 U706 ( .A1(n638), .A2(n722), .ZN(G54) );
  XOR2_X1 U707 ( .A(G101), .B(n639), .Z(G3) );
  XOR2_X1 U708 ( .A(G104), .B(KEYINPUT111), .Z(n641) );
  NAND2_X1 U709 ( .A1(n642), .A2(n653), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n641), .B(n640), .ZN(G6) );
  XNOR2_X1 U711 ( .A(G107), .B(KEYINPUT27), .ZN(n646) );
  XOR2_X1 U712 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n644) );
  NAND2_X1 U713 ( .A1(n656), .A2(n642), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U715 ( .A(n646), .B(n645), .ZN(G9) );
  XOR2_X1 U716 ( .A(G128), .B(KEYINPUT29), .Z(n648) );
  NAND2_X1 U717 ( .A1(n656), .A2(n650), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(G30) );
  XNOR2_X1 U719 ( .A(G143), .B(n649), .ZN(G45) );
  XOR2_X1 U720 ( .A(G146), .B(KEYINPUT113), .Z(n652) );
  NAND2_X1 U721 ( .A1(n650), .A2(n653), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(G48) );
  NAND2_X1 U723 ( .A1(n653), .A2(n657), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n654), .B(KEYINPUT114), .ZN(n655) );
  XNOR2_X1 U725 ( .A(G113), .B(n655), .ZN(G15) );
  NAND2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n658), .B(G116), .ZN(G18) );
  XNOR2_X1 U728 ( .A(n659), .B(G125), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n660), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U730 ( .A(G134), .B(n661), .ZN(G36) );
  XOR2_X1 U731 ( .A(G140), .B(n662), .Z(G42) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(KEYINPUT50), .ZN(n672) );
  NOR2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n668), .B(KEYINPUT49), .ZN(n669) );
  NAND2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  OR2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n675) );
  INV_X1 U738 ( .A(n673), .ZN(n674) );
  AND2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U740 ( .A(KEYINPUT51), .B(n676), .Z(n677) );
  XOR2_X1 U741 ( .A(KEYINPUT115), .B(n677), .Z(n678) );
  NOR2_X1 U742 ( .A1(n710), .A2(n678), .ZN(n692) );
  NOR2_X1 U743 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U744 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U745 ( .A(KEYINPUT116), .B(n683), .Z(n688) );
  NOR2_X1 U746 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U747 ( .A(KEYINPUT117), .B(n686), .ZN(n687) );
  NAND2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U749 ( .A1(n689), .A2(n709), .ZN(n690) );
  XOR2_X1 U750 ( .A(KEYINPUT118), .B(n690), .Z(n691) );
  NOR2_X1 U751 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U752 ( .A(n693), .B(KEYINPUT52), .ZN(n694) );
  NOR2_X1 U753 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U754 ( .A(KEYINPUT119), .B(n696), .ZN(n708) );
  INV_X1 U755 ( .A(n697), .ZN(n698) );
  NAND2_X1 U756 ( .A1(n698), .A2(n610), .ZN(n703) );
  NAND2_X1 U757 ( .A1(n700), .A2(n610), .ZN(n701) );
  XNOR2_X1 U758 ( .A(n701), .B(KEYINPUT80), .ZN(n702) );
  NAND2_X1 U759 ( .A1(n703), .A2(n702), .ZN(n705) );
  NOR2_X1 U760 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U761 ( .A1(G953), .A2(n706), .ZN(n707) );
  NAND2_X1 U762 ( .A1(n708), .A2(n707), .ZN(n712) );
  NOR2_X1 U763 ( .A1(n710), .A2(n369), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U765 ( .A(n713), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U766 ( .A1(n714), .A2(G478), .ZN(n715) );
  XOR2_X1 U767 ( .A(n716), .B(n715), .Z(n717) );
  NOR2_X1 U768 ( .A1(n722), .A2(n717), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n718), .A2(G217), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U771 ( .A1(n722), .A2(n721), .ZN(G66) );
  XNOR2_X1 U772 ( .A(G101), .B(n723), .ZN(n724) );
  XNOR2_X1 U773 ( .A(n724), .B(KEYINPUT122), .ZN(n726) );
  NOR2_X1 U774 ( .A1(G898), .A2(n744), .ZN(n725) );
  NOR2_X1 U775 ( .A1(n726), .A2(n725), .ZN(n736) );
  NAND2_X1 U776 ( .A1(n727), .A2(n744), .ZN(n728) );
  XOR2_X1 U777 ( .A(KEYINPUT121), .B(n728), .Z(n732) );
  NAND2_X1 U778 ( .A1(G953), .A2(G224), .ZN(n729) );
  XNOR2_X1 U779 ( .A(KEYINPUT61), .B(n729), .ZN(n730) );
  NAND2_X1 U780 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U781 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U782 ( .A(n733), .B(KEYINPUT124), .ZN(n734) );
  XOR2_X1 U783 ( .A(KEYINPUT123), .B(n734), .Z(n735) );
  XNOR2_X1 U784 ( .A(n736), .B(n735), .ZN(G69) );
  XNOR2_X1 U785 ( .A(n737), .B(KEYINPUT125), .ZN(n739) );
  XNOR2_X1 U786 ( .A(n739), .B(n738), .ZN(n743) );
  XOR2_X1 U787 ( .A(G227), .B(n743), .Z(n740) );
  NAND2_X1 U788 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U789 ( .A1(G953), .A2(n741), .ZN(n742) );
  XNOR2_X1 U790 ( .A(n742), .B(KEYINPUT126), .ZN(n747) );
  XOR2_X1 U791 ( .A(n743), .B(n700), .Z(n745) );
  NAND2_X1 U792 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U793 ( .A1(n747), .A2(n746), .ZN(G72) );
  XOR2_X1 U794 ( .A(G119), .B(n748), .Z(G21) );
  XOR2_X1 U795 ( .A(n749), .B(G110), .Z(G12) );
  XNOR2_X1 U796 ( .A(n750), .B(G131), .ZN(G33) );
  XNOR2_X1 U797 ( .A(n751), .B(G137), .ZN(G39) );
endmodule

