

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U549 ( .A1(n806), .A2(n805), .ZN(n836) );
  NOR2_X2 U550 ( .A1(n688), .A2(G164), .ZN(n690) );
  XNOR2_X1 U551 ( .A(KEYINPUT89), .B(n686), .ZN(n769) );
  NOR2_X1 U552 ( .A1(n693), .A2(n980), .ZN(n695) );
  NOR2_X1 U553 ( .A1(n710), .A2(n975), .ZN(n696) );
  INV_X1 U554 ( .A(KEYINPUT29), .ZN(n719) );
  INV_X1 U555 ( .A(G1384), .ZN(n687) );
  AND2_X1 U556 ( .A1(n744), .A2(n743), .ZN(n745) );
  INV_X1 U557 ( .A(KEYINPUT64), .ZN(n689) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  NOR2_X1 U559 ( .A1(G651), .A2(G543), .ZN(n653) );
  NOR2_X1 U560 ( .A1(G651), .A2(n630), .ZN(n649) );
  NOR2_X1 U561 ( .A1(n523), .A2(n522), .ZN(G160) );
  NAND2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n513) );
  XNOR2_X2 U563 ( .A(n513), .B(KEYINPUT65), .ZN(n892) );
  NAND2_X1 U564 ( .A1(n892), .A2(G113), .ZN(n516) );
  INV_X1 U565 ( .A(G2104), .ZN(n519) );
  NOR2_X4 U566 ( .A1(G2105), .A2(n519), .ZN(n886) );
  NAND2_X1 U567 ( .A1(G101), .A2(n886), .ZN(n514) );
  XOR2_X1 U568 ( .A(KEYINPUT23), .B(n514), .Z(n515) );
  NAND2_X1 U569 ( .A1(n516), .A2(n515), .ZN(n523) );
  XNOR2_X1 U570 ( .A(KEYINPUT17), .B(n517), .ZN(n518) );
  INV_X1 U571 ( .A(n518), .ZN(n888) );
  NAND2_X1 U572 ( .A1(G137), .A2(n888), .ZN(n521) );
  AND2_X1 U573 ( .A1(n519), .A2(G2105), .ZN(n893) );
  NAND2_X1 U574 ( .A1(G125), .A2(n893), .ZN(n520) );
  NAND2_X1 U575 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n888), .A2(G138), .ZN(n526) );
  NAND2_X1 U577 ( .A1(n886), .A2(G102), .ZN(n524) );
  XNOR2_X1 U578 ( .A(n524), .B(KEYINPUT86), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U580 ( .A(n527), .B(KEYINPUT87), .ZN(n532) );
  NAND2_X1 U581 ( .A1(G114), .A2(n892), .ZN(n529) );
  NAND2_X1 U582 ( .A1(G126), .A2(n893), .ZN(n528) );
  NAND2_X1 U583 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U584 ( .A(n530), .B(KEYINPUT85), .ZN(n531) );
  AND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U586 ( .A(n533), .B(KEYINPUT88), .ZN(G164) );
  XNOR2_X1 U587 ( .A(G2451), .B(G2427), .ZN(n543) );
  XOR2_X1 U588 ( .A(G2430), .B(G2443), .Z(n535) );
  XNOR2_X1 U589 ( .A(G2435), .B(KEYINPUT106), .ZN(n534) );
  XNOR2_X1 U590 ( .A(n535), .B(n534), .ZN(n539) );
  XOR2_X1 U591 ( .A(G2438), .B(G2454), .Z(n537) );
  XNOR2_X1 U592 ( .A(G1341), .B(G1348), .ZN(n536) );
  XNOR2_X1 U593 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U594 ( .A(n539), .B(n538), .Z(n541) );
  XNOR2_X1 U595 ( .A(G2446), .B(KEYINPUT107), .ZN(n540) );
  XNOR2_X1 U596 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n543), .B(n542), .ZN(n544) );
  AND2_X1 U598 ( .A1(n544), .A2(G14), .ZN(G401) );
  INV_X1 U599 ( .A(G651), .ZN(n549) );
  NOR2_X1 U600 ( .A1(G543), .A2(n549), .ZN(n545) );
  XOR2_X1 U601 ( .A(KEYINPUT1), .B(n545), .Z(n648) );
  NAND2_X1 U602 ( .A1(G64), .A2(n648), .ZN(n547) );
  XOR2_X1 U603 ( .A(KEYINPUT0), .B(G543), .Z(n630) );
  NAND2_X1 U604 ( .A1(G52), .A2(n649), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U606 ( .A(KEYINPUT67), .B(n548), .Z(n555) );
  NOR2_X1 U607 ( .A1(n630), .A2(n549), .ZN(n654) );
  NAND2_X1 U608 ( .A1(n654), .A2(G77), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n550), .B(KEYINPUT68), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G90), .A2(n653), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U613 ( .A1(n555), .A2(n554), .ZN(G171) );
  AND2_X1 U614 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  NAND2_X1 U617 ( .A1(G63), .A2(n648), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G51), .A2(n649), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n558), .B(KEYINPUT75), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n559), .B(KEYINPUT6), .ZN(n566) );
  XNOR2_X1 U622 ( .A(KEYINPUT74), .B(KEYINPUT5), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n653), .A2(G89), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G76), .A2(n654), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U629 ( .A(KEYINPUT7), .B(n567), .ZN(G168) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U632 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U633 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n570) );
  INV_X1 U634 ( .A(G223), .ZN(n838) );
  NAND2_X1 U635 ( .A1(G567), .A2(n838), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G234) );
  NAND2_X1 U637 ( .A1(G56), .A2(n648), .ZN(n571) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n571), .Z(n577) );
  NAND2_X1 U639 ( .A1(n653), .A2(G81), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G68), .A2(n654), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT13), .B(n575), .Z(n576) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n649), .A2(G43), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n980) );
  INV_X1 U647 ( .A(G860), .ZN(n600) );
  OR2_X1 U648 ( .A1(n980), .A2(n600), .ZN(G153) );
  INV_X1 U649 ( .A(G171), .ZN(G301) );
  NAND2_X1 U650 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n649), .A2(G54), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G92), .A2(n653), .ZN(n581) );
  NAND2_X1 U653 ( .A1(G79), .A2(n654), .ZN(n580) );
  NAND2_X1 U654 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U655 ( .A1(G66), .A2(n648), .ZN(n582) );
  XNOR2_X1 U656 ( .A(KEYINPUT73), .B(n582), .ZN(n583) );
  NOR2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U659 ( .A(KEYINPUT15), .B(n587), .Z(n975) );
  INV_X1 U660 ( .A(G868), .ZN(n668) );
  NAND2_X1 U661 ( .A1(n975), .A2(n668), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U663 ( .A1(G65), .A2(n648), .ZN(n590) );
  XNOR2_X1 U664 ( .A(n590), .B(KEYINPUT70), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G53), .A2(n649), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G91), .A2(n653), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G78), .A2(n654), .ZN(n593) );
  XNOR2_X1 U669 ( .A(KEYINPUT69), .B(n593), .ZN(n594) );
  NOR2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(G299) );
  NOR2_X1 U672 ( .A1(G286), .A2(n668), .ZN(n599) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U674 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U675 ( .A1(n600), .A2(G559), .ZN(n601) );
  INV_X1 U676 ( .A(n975), .ZN(n708) );
  NAND2_X1 U677 ( .A1(n601), .A2(n708), .ZN(n602) );
  XNOR2_X1 U678 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U679 ( .A1(G868), .A2(n980), .ZN(n605) );
  NAND2_X1 U680 ( .A1(G868), .A2(n708), .ZN(n603) );
  NOR2_X1 U681 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n605), .A2(n604), .ZN(G282) );
  XOR2_X1 U683 ( .A(G2100), .B(KEYINPUT78), .Z(n616) );
  NAND2_X1 U684 ( .A1(G111), .A2(n892), .ZN(n607) );
  NAND2_X1 U685 ( .A1(G99), .A2(n886), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n614) );
  NAND2_X1 U687 ( .A1(G123), .A2(n893), .ZN(n608) );
  XNOR2_X1 U688 ( .A(n608), .B(KEYINPUT18), .ZN(n609) );
  XNOR2_X1 U689 ( .A(n609), .B(KEYINPUT76), .ZN(n611) );
  NAND2_X1 U690 ( .A1(G135), .A2(n888), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U692 ( .A(KEYINPUT77), .B(n612), .Z(n613) );
  NOR2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n928) );
  XNOR2_X1 U694 ( .A(G2096), .B(n928), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(G156) );
  NAND2_X1 U696 ( .A1(n708), .A2(G559), .ZN(n666) );
  XNOR2_X1 U697 ( .A(n980), .B(n666), .ZN(n617) );
  NOR2_X1 U698 ( .A1(n617), .A2(G860), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G67), .A2(n648), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G93), .A2(n653), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G55), .A2(n649), .ZN(n621) );
  NAND2_X1 U703 ( .A1(G80), .A2(n654), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n622) );
  OR2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n669) );
  XOR2_X1 U706 ( .A(n624), .B(n669), .Z(G145) );
  NAND2_X1 U707 ( .A1(n649), .A2(G49), .ZN(n625) );
  XOR2_X1 U708 ( .A(KEYINPUT79), .B(n625), .Z(n627) );
  NAND2_X1 U709 ( .A1(G651), .A2(G74), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U711 ( .A1(n648), .A2(n628), .ZN(n629) );
  XNOR2_X1 U712 ( .A(n629), .B(KEYINPUT80), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G87), .A2(n630), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G73), .A2(n654), .ZN(n633) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n633), .Z(n638) );
  NAND2_X1 U717 ( .A1(G61), .A2(n648), .ZN(n635) );
  NAND2_X1 U718 ( .A1(G86), .A2(n653), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U720 ( .A(KEYINPUT81), .B(n636), .Z(n637) );
  NOR2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n649), .A2(G48), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U724 ( .A1(G62), .A2(n648), .ZN(n642) );
  NAND2_X1 U725 ( .A1(G75), .A2(n654), .ZN(n641) );
  NAND2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n653), .A2(G88), .ZN(n643) );
  XOR2_X1 U728 ( .A(KEYINPUT82), .B(n643), .Z(n644) );
  NOR2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n649), .A2(G50), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(G303) );
  INV_X1 U732 ( .A(G303), .ZN(G166) );
  NAND2_X1 U733 ( .A1(G60), .A2(n648), .ZN(n651) );
  NAND2_X1 U734 ( .A1(G47), .A2(n649), .ZN(n650) );
  NAND2_X1 U735 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U736 ( .A(KEYINPUT66), .B(n652), .Z(n658) );
  NAND2_X1 U737 ( .A1(G85), .A2(n653), .ZN(n656) );
  NAND2_X1 U738 ( .A1(G72), .A2(n654), .ZN(n655) );
  AND2_X1 U739 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U740 ( .A1(n658), .A2(n657), .ZN(G290) );
  XOR2_X1 U741 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n659) );
  XNOR2_X1 U742 ( .A(G305), .B(n659), .ZN(n660) );
  XNOR2_X1 U743 ( .A(n660), .B(n669), .ZN(n662) );
  INV_X1 U744 ( .A(G299), .ZN(n711) );
  XNOR2_X1 U745 ( .A(n711), .B(G166), .ZN(n661) );
  XNOR2_X1 U746 ( .A(n662), .B(n661), .ZN(n663) );
  XOR2_X1 U747 ( .A(n663), .B(G290), .Z(n664) );
  XNOR2_X1 U748 ( .A(n980), .B(n664), .ZN(n665) );
  XNOR2_X1 U749 ( .A(G288), .B(n665), .ZN(n909) );
  XNOR2_X1 U750 ( .A(n666), .B(n909), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n667), .A2(G868), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U753 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U758 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U760 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U761 ( .A1(G219), .A2(G220), .ZN(n676) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U763 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U764 ( .A1(G96), .A2(n678), .ZN(n843) );
  AND2_X1 U765 ( .A1(G2106), .A2(n843), .ZN(n683) );
  NAND2_X1 U766 ( .A1(G69), .A2(G120), .ZN(n679) );
  NOR2_X1 U767 ( .A1(G237), .A2(n679), .ZN(n680) );
  NAND2_X1 U768 ( .A1(G108), .A2(n680), .ZN(n842) );
  NAND2_X1 U769 ( .A1(G567), .A2(n842), .ZN(n681) );
  XOR2_X1 U770 ( .A(KEYINPUT84), .B(n681), .Z(n682) );
  NOR2_X1 U771 ( .A1(n683), .A2(n682), .ZN(G319) );
  INV_X1 U772 ( .A(G319), .ZN(n685) );
  NAND2_X1 U773 ( .A1(G483), .A2(G661), .ZN(n684) );
  NOR2_X1 U774 ( .A1(n685), .A2(n684), .ZN(n841) );
  NAND2_X1 U775 ( .A1(n841), .A2(G36), .ZN(G176) );
  NAND2_X1 U776 ( .A1(G40), .A2(G160), .ZN(n686) );
  NAND2_X1 U777 ( .A1(n769), .A2(n687), .ZN(n688) );
  XNOR2_X2 U778 ( .A(n690), .B(n689), .ZN(n736) );
  INV_X1 U779 ( .A(n736), .ZN(n699) );
  NAND2_X1 U780 ( .A1(n699), .A2(G1996), .ZN(n692) );
  INV_X1 U781 ( .A(KEYINPUT26), .ZN(n691) );
  XNOR2_X1 U782 ( .A(n692), .B(n691), .ZN(n693) );
  NAND2_X1 U783 ( .A1(n736), .A2(G1341), .ZN(n694) );
  NAND2_X1 U784 ( .A1(n695), .A2(n694), .ZN(n710) );
  XOR2_X1 U785 ( .A(n696), .B(KEYINPUT96), .Z(n705) );
  INV_X1 U786 ( .A(n736), .ZN(n721) );
  NOR2_X1 U787 ( .A1(G1348), .A2(n721), .ZN(n698) );
  NOR2_X1 U788 ( .A1(G2067), .A2(n736), .ZN(n697) );
  NOR2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n703) );
  NAND2_X1 U790 ( .A1(G2072), .A2(n699), .ZN(n700) );
  XNOR2_X1 U791 ( .A(n700), .B(KEYINPUT27), .ZN(n702) );
  INV_X1 U792 ( .A(G1956), .ZN(n997) );
  NOR2_X1 U793 ( .A1(n721), .A2(n997), .ZN(n701) );
  NOR2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n712) );
  NAND2_X1 U795 ( .A1(n711), .A2(n712), .ZN(n706) );
  AND2_X1 U796 ( .A1(n703), .A2(n706), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n718) );
  INV_X1 U798 ( .A(n706), .ZN(n707) );
  NOR2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n716) );
  NOR2_X1 U801 ( .A1(n712), .A2(n711), .ZN(n714) );
  INV_X1 U802 ( .A(KEYINPUT28), .ZN(n713) );
  XNOR2_X1 U803 ( .A(n714), .B(n713), .ZN(n715) );
  AND2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U805 ( .A1(n718), .A2(n717), .ZN(n720) );
  XNOR2_X1 U806 ( .A(n720), .B(n719), .ZN(n725) );
  XOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .Z(n945) );
  NAND2_X1 U808 ( .A1(n945), .A2(n721), .ZN(n723) );
  NAND2_X1 U809 ( .A1(n736), .A2(G1961), .ZN(n722) );
  NAND2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n726) );
  OR2_X1 U811 ( .A1(G301), .A2(n726), .ZN(n724) );
  NAND2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n735) );
  NAND2_X1 U813 ( .A1(G301), .A2(n726), .ZN(n727) );
  XNOR2_X1 U814 ( .A(n727), .B(KEYINPUT97), .ZN(n732) );
  NAND2_X1 U815 ( .A1(n736), .A2(G8), .ZN(n813) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n813), .ZN(n749) );
  NOR2_X1 U817 ( .A1(n736), .A2(G2084), .ZN(n746) );
  NOR2_X1 U818 ( .A1(n749), .A2(n746), .ZN(n728) );
  NAND2_X1 U819 ( .A1(G8), .A2(n728), .ZN(n729) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n729), .ZN(n730) );
  NOR2_X1 U821 ( .A1(n730), .A2(G168), .ZN(n731) );
  NOR2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U823 ( .A(KEYINPUT31), .B(n733), .Z(n734) );
  NAND2_X1 U824 ( .A1(n735), .A2(n734), .ZN(n747) );
  NAND2_X1 U825 ( .A1(n747), .A2(G286), .ZN(n744) );
  INV_X1 U826 ( .A(G8), .ZN(n742) );
  NOR2_X1 U827 ( .A1(n736), .A2(G2090), .ZN(n737) );
  XNOR2_X1 U828 ( .A(n737), .B(KEYINPUT98), .ZN(n739) );
  NOR2_X1 U829 ( .A1(n813), .A2(G1971), .ZN(n738) );
  NOR2_X1 U830 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U831 ( .A1(n740), .A2(G303), .ZN(n741) );
  OR2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U833 ( .A(n745), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U834 ( .A1(G8), .A2(n746), .ZN(n751) );
  INV_X1 U835 ( .A(n747), .ZN(n748) );
  NOR2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n753), .A2(n752), .ZN(n807) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n968) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n754) );
  NOR2_X1 U841 ( .A1(n968), .A2(n754), .ZN(n755) );
  XOR2_X1 U842 ( .A(KEYINPUT99), .B(n755), .Z(n757) );
  INV_X1 U843 ( .A(KEYINPUT33), .ZN(n756) );
  AND2_X1 U844 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U845 ( .A1(n807), .A2(n758), .ZN(n762) );
  NAND2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n969) );
  INV_X1 U847 ( .A(n969), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n759), .A2(n813), .ZN(n760) );
  OR2_X1 U849 ( .A1(KEYINPUT33), .A2(n760), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U851 ( .A(n763), .B(KEYINPUT100), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n968), .A2(KEYINPUT33), .ZN(n764) );
  NOR2_X1 U853 ( .A1(n813), .A2(n764), .ZN(n765) );
  NOR2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U855 ( .A(n767), .B(KEYINPUT101), .ZN(n806) );
  XNOR2_X1 U856 ( .A(G1981), .B(KEYINPUT102), .ZN(n768) );
  XNOR2_X1 U857 ( .A(n768), .B(G305), .ZN(n972) );
  XNOR2_X1 U858 ( .A(G1986), .B(G290), .ZN(n982) );
  OR2_X1 U859 ( .A1(G1384), .A2(G164), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n800) );
  INV_X1 U861 ( .A(n800), .ZN(n831) );
  NAND2_X1 U862 ( .A1(n982), .A2(n831), .ZN(n803) );
  NAND2_X1 U863 ( .A1(G116), .A2(n892), .ZN(n772) );
  NAND2_X1 U864 ( .A1(G128), .A2(n893), .ZN(n771) );
  NAND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U866 ( .A(KEYINPUT35), .B(n773), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n888), .A2(G140), .ZN(n774) );
  XNOR2_X1 U868 ( .A(n774), .B(KEYINPUT90), .ZN(n776) );
  NAND2_X1 U869 ( .A1(G104), .A2(n886), .ZN(n775) );
  NAND2_X1 U870 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U871 ( .A(KEYINPUT34), .B(n777), .Z(n778) );
  NAND2_X1 U872 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U873 ( .A(KEYINPUT36), .B(n780), .Z(n904) );
  XNOR2_X1 U874 ( .A(G2067), .B(KEYINPUT37), .ZN(n829) );
  OR2_X1 U875 ( .A1(n904), .A2(n829), .ZN(n781) );
  XNOR2_X1 U876 ( .A(KEYINPUT91), .B(n781), .ZN(n940) );
  NAND2_X1 U877 ( .A1(n831), .A2(n940), .ZN(n826) );
  NAND2_X1 U878 ( .A1(G119), .A2(n893), .ZN(n783) );
  NAND2_X1 U879 ( .A1(G95), .A2(n886), .ZN(n782) );
  NAND2_X1 U880 ( .A1(n783), .A2(n782), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n892), .A2(G107), .ZN(n784) );
  XNOR2_X1 U882 ( .A(n784), .B(KEYINPUT92), .ZN(n786) );
  NAND2_X1 U883 ( .A1(G131), .A2(n888), .ZN(n785) );
  NAND2_X1 U884 ( .A1(n786), .A2(n785), .ZN(n787) );
  OR2_X1 U885 ( .A1(n788), .A2(n787), .ZN(n899) );
  XOR2_X1 U886 ( .A(KEYINPUT93), .B(G1991), .Z(n949) );
  AND2_X1 U887 ( .A1(n899), .A2(n949), .ZN(n799) );
  NAND2_X1 U888 ( .A1(G105), .A2(n886), .ZN(n789) );
  XNOR2_X1 U889 ( .A(n789), .B(KEYINPUT38), .ZN(n796) );
  NAND2_X1 U890 ( .A1(G117), .A2(n892), .ZN(n791) );
  NAND2_X1 U891 ( .A1(G141), .A2(n888), .ZN(n790) );
  NAND2_X1 U892 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U893 ( .A1(n893), .A2(G129), .ZN(n792) );
  XOR2_X1 U894 ( .A(KEYINPUT94), .B(n792), .Z(n793) );
  NOR2_X1 U895 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U896 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U897 ( .A(KEYINPUT95), .B(n797), .ZN(n903) );
  INV_X1 U898 ( .A(G1996), .ZN(n818) );
  NOR2_X1 U899 ( .A1(n903), .A2(n818), .ZN(n798) );
  NOR2_X1 U900 ( .A1(n799), .A2(n798), .ZN(n926) );
  NOR2_X1 U901 ( .A1(n926), .A2(n800), .ZN(n823) );
  INV_X1 U902 ( .A(n823), .ZN(n801) );
  AND2_X1 U903 ( .A1(n826), .A2(n801), .ZN(n802) );
  AND2_X1 U904 ( .A1(n803), .A2(n802), .ZN(n817) );
  INV_X1 U905 ( .A(n817), .ZN(n804) );
  OR2_X1 U906 ( .A1(n972), .A2(n804), .ZN(n805) );
  NOR2_X1 U907 ( .A1(G2090), .A2(G303), .ZN(n808) );
  NAND2_X1 U908 ( .A1(G8), .A2(n808), .ZN(n809) );
  NAND2_X1 U909 ( .A1(n807), .A2(n809), .ZN(n810) );
  AND2_X1 U910 ( .A1(n810), .A2(n813), .ZN(n815) );
  NOR2_X1 U911 ( .A1(G1981), .A2(G305), .ZN(n811) );
  XOR2_X1 U912 ( .A(n811), .B(KEYINPUT24), .Z(n812) );
  NOR2_X1 U913 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U914 ( .A1(n815), .A2(n814), .ZN(n816) );
  AND2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n834) );
  AND2_X1 U916 ( .A1(n818), .A2(n903), .ZN(n921) );
  NOR2_X1 U917 ( .A1(n949), .A2(n899), .ZN(n924) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n819) );
  XOR2_X1 U919 ( .A(n819), .B(KEYINPUT103), .Z(n820) );
  NOR2_X1 U920 ( .A1(n924), .A2(n820), .ZN(n821) );
  XNOR2_X1 U921 ( .A(n821), .B(KEYINPUT104), .ZN(n822) );
  NOR2_X1 U922 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U923 ( .A1(n921), .A2(n824), .ZN(n825) );
  XNOR2_X1 U924 ( .A(n825), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U925 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U926 ( .A(KEYINPUT105), .B(n828), .Z(n830) );
  NAND2_X1 U927 ( .A1(n904), .A2(n829), .ZN(n929) );
  NAND2_X1 U928 ( .A1(n830), .A2(n929), .ZN(n832) );
  AND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U930 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U932 ( .A(n837), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n838), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U935 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(G188) );
  XOR2_X1 U938 ( .A(G96), .B(KEYINPUT108), .Z(G221) );
  NOR2_X1 U939 ( .A1(n843), .A2(n842), .ZN(G325) );
  XNOR2_X1 U940 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  INV_X1 U943 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U944 ( .A(G1996), .B(KEYINPUT41), .ZN(n853) );
  XOR2_X1 U945 ( .A(G1971), .B(G1956), .Z(n845) );
  XNOR2_X1 U946 ( .A(G1991), .B(G1986), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U948 ( .A(G1976), .B(G1981), .Z(n847) );
  XNOR2_X1 U949 ( .A(G1966), .B(G1961), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U951 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U952 ( .A(KEYINPUT112), .B(G2474), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U955 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U956 ( .A(KEYINPUT110), .B(G2678), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U958 ( .A(KEYINPUT42), .B(G2090), .Z(n857) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U961 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U962 ( .A(G2100), .B(G2096), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n863) );
  XOR2_X1 U964 ( .A(G2078), .B(G2084), .Z(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(G227) );
  NAND2_X1 U966 ( .A1(G124), .A2(n893), .ZN(n864) );
  XOR2_X1 U967 ( .A(KEYINPUT44), .B(n864), .Z(n865) );
  XNOR2_X1 U968 ( .A(n865), .B(KEYINPUT113), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G136), .A2(n888), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U971 ( .A(KEYINPUT114), .B(n868), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G112), .A2(n892), .ZN(n870) );
  NAND2_X1 U973 ( .A1(G100), .A2(n886), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U975 ( .A1(n872), .A2(n871), .ZN(G162) );
  XOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n874) );
  XNOR2_X1 U977 ( .A(G160), .B(KEYINPUT117), .ZN(n873) );
  XNOR2_X1 U978 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U979 ( .A(n875), .B(n928), .Z(n885) );
  NAND2_X1 U980 ( .A1(G115), .A2(n892), .ZN(n877) );
  NAND2_X1 U981 ( .A1(G127), .A2(n893), .ZN(n876) );
  NAND2_X1 U982 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U983 ( .A(n878), .B(KEYINPUT47), .ZN(n880) );
  NAND2_X1 U984 ( .A1(G103), .A2(n886), .ZN(n879) );
  NAND2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n888), .A2(G139), .ZN(n881) );
  XOR2_X1 U987 ( .A(KEYINPUT118), .B(n881), .Z(n882) );
  NOR2_X1 U988 ( .A1(n883), .A2(n882), .ZN(n931) );
  XNOR2_X1 U989 ( .A(n931), .B(G162), .ZN(n884) );
  XNOR2_X1 U990 ( .A(n885), .B(n884), .ZN(n902) );
  NAND2_X1 U991 ( .A1(n886), .A2(G106), .ZN(n887) );
  XNOR2_X1 U992 ( .A(n887), .B(KEYINPUT116), .ZN(n890) );
  NAND2_X1 U993 ( .A1(G142), .A2(n888), .ZN(n889) );
  NAND2_X1 U994 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U995 ( .A(n891), .B(KEYINPUT45), .ZN(n898) );
  NAND2_X1 U996 ( .A1(G118), .A2(n892), .ZN(n895) );
  NAND2_X1 U997 ( .A1(G130), .A2(n893), .ZN(n894) );
  NAND2_X1 U998 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U999 ( .A(KEYINPUT115), .B(n896), .ZN(n897) );
  NAND2_X1 U1000 ( .A1(n898), .A2(n897), .ZN(n900) );
  XOR2_X1 U1001 ( .A(n900), .B(n899), .Z(n901) );
  XOR2_X1 U1002 ( .A(n902), .B(n901), .Z(n906) );
  XOR2_X1 U1003 ( .A(n904), .B(n903), .Z(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n907), .B(G164), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n908), .ZN(G395) );
  XNOR2_X1 U1007 ( .A(G286), .B(n975), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(G171), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n912), .ZN(G397) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(KEYINPUT119), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(n915), .A2(G319), .ZN(n916) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n916), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(KEYINPUT120), .B(n917), .ZN(n919) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n920) );
  NOR2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1023 ( .A(KEYINPUT51), .B(n922), .Z(n938) );
  XOR2_X1 U1024 ( .A(G160), .B(G2084), .Z(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n936) );
  XOR2_X1 U1029 ( .A(G2072), .B(n931), .Z(n933) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1032 ( .A(KEYINPUT50), .B(n934), .Z(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT52), .B(n941), .Z(n942) );
  NOR2_X1 U1037 ( .A1(KEYINPUT55), .A2(n942), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(KEYINPUT121), .B(n943), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(G29), .ZN(n996) );
  XOR2_X1 U1040 ( .A(G2090), .B(G35), .Z(n960) );
  XNOR2_X1 U1041 ( .A(G1996), .B(G32), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(n945), .B(G27), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(KEYINPUT122), .B(n948), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(G25), .B(n949), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1049 ( .A(G2072), .B(G33), .Z(n954) );
  NAND2_X1 U1050 ( .A1(G28), .A2(n954), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(n957), .B(KEYINPUT53), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(n958), .B(KEYINPUT123), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(G34), .B(G2084), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(KEYINPUT55), .B(n964), .ZN(n966) );
  INV_X1 U1059 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n967), .A2(G11), .ZN(n994) );
  XOR2_X1 U1062 ( .A(KEYINPUT56), .B(G16), .Z(n992) );
  INV_X1 U1063 ( .A(n968), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n990) );
  XOR2_X1 U1065 ( .A(G168), .B(G1966), .Z(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1067 ( .A(KEYINPUT57), .B(n973), .Z(n988) );
  XNOR2_X1 U1068 ( .A(G1971), .B(G166), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n974), .B(KEYINPUT124), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(n975), .B(G1348), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(G299), .B(G1956), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(G171), .B(G1961), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G1341), .B(n980), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n1023) );
  XOR2_X1 U1084 ( .A(G1961), .B(G5), .Z(n1011) );
  XOR2_X1 U1085 ( .A(G1341), .B(G19), .Z(n999) );
  XNOR2_X1 U1086 ( .A(n997), .B(G20), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1005) );
  XOR2_X1 U1088 ( .A(G1981), .B(G6), .Z(n1003) );
  XOR2_X1 U1089 ( .A(G1348), .B(G4), .Z(n1000) );
  XNOR2_X1 U1090 ( .A(KEYINPUT125), .B(n1000), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(n1001), .B(KEYINPUT59), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1006), .Z(n1008) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G21), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(KEYINPUT126), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1018) );
  XNOR2_X1 U1099 ( .A(G1971), .B(G22), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G23), .B(G1976), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(G1986), .B(G24), .Z(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(KEYINPUT58), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1019), .Z(n1020) );
  NOR2_X1 U1107 ( .A1(G16), .A2(n1020), .ZN(n1021) );
  XOR2_X1 U1108 ( .A(KEYINPUT127), .B(n1021), .Z(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(n1024), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

