//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n202));
  XOR2_X1   g001(.A(G127gat), .B(G134gat), .Z(new_n203));
  INV_X1    g002(.A(G120gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G113gat), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G120gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT71), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n208), .B1(new_n205), .B2(new_n207), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n203), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n205), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n204), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n207), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G162gat), .ZN(new_n229));
  OR2_X1    g028(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n225), .B(new_n228), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT78), .B1(new_n226), .B2(new_n227), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n227), .A2(KEYINPUT78), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n223), .A2(new_n233), .A3(new_n224), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n202), .B1(new_n220), .B2(new_n239), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n223), .B(new_n224), .C1(new_n226), .C2(new_n227), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT79), .B(G155gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G162gat), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n241), .B1(new_n243), .B2(KEYINPUT2), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT3), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n234), .A2(new_n247), .A3(new_n238), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n220), .A3(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n244), .A2(new_n245), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n250), .A2(KEYINPUT4), .A3(new_n213), .A4(new_n219), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n240), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT5), .ZN(new_n253));
  NAND2_X1  g052(.A1(G225gat), .A2(G233gat), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n252), .A2(KEYINPUT80), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT80), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n240), .A2(new_n249), .A3(new_n251), .A4(new_n254), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(KEYINPUT5), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n220), .B(new_n239), .ZN(new_n260));
  INV_X1    g059(.A(new_n254), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n253), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n257), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G1gat), .B(G29gat), .Z(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT0), .ZN(new_n266));
  XNOR2_X1  g065(.A(G57gat), .B(G85gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(KEYINPUT6), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT89), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n255), .A2(new_n258), .B1(new_n257), .B2(new_n262), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(new_n268), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT89), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT6), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n268), .A3(new_n263), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n268), .B(KEYINPUT86), .Z(new_n278));
  OAI211_X1 g077(.A(new_n276), .B(new_n277), .C1(new_n272), .C2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n271), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(G197gat), .B(G204gat), .Z(new_n281));
  AOI21_X1  g080(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(G211gat), .B(G218gat), .Z(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n281), .B2(new_n282), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n247), .B1(new_n288), .B2(KEYINPUT29), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n239), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(G228gat), .A3(G233gat), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n286), .A2(KEYINPUT76), .A3(new_n287), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT76), .B1(new_n286), .B2(new_n287), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n248), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(KEYINPUT83), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT83), .B1(new_n294), .B2(new_n296), .ZN(new_n299));
  OR3_X1    g098(.A1(new_n291), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n296), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n288), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n302), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(KEYINPUT29), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT3), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n301), .B1(new_n306), .B2(new_n250), .ZN(new_n307));
  NAND2_X1  g106(.A1(G228gat), .A2(G233gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G78gat), .B(G106gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(G50gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G22gat), .ZN(new_n314));
  INV_X1    g113(.A(G22gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(KEYINPUT84), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n316), .B2(new_n313), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n309), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n317), .ZN(new_n319));
  INV_X1    g118(.A(new_n309), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n291), .A2(new_n298), .A3(new_n299), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT35), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n318), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G8gat), .B(G36gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G64gat), .B(G92gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n325), .B(new_n326), .Z(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT66), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT64), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n334), .A2(G183gat), .A3(G190gat), .ZN(new_n335));
  INV_X1    g134(.A(G183gat), .ZN(new_n336));
  INV_X1    g135(.A(G190gat), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT65), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n333), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n329), .B1(new_n332), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n330), .B(KEYINPUT64), .ZN(new_n341));
  INV_X1    g140(.A(new_n333), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT65), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n334), .B1(G183gat), .B2(G190gat), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n341), .A2(KEYINPUT66), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT23), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(G169gat), .B2(G176gat), .ZN(new_n350));
  INV_X1    g149(.A(G169gat), .ZN(new_n351));
  INV_X1    g150(.A(G176gat), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n348), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n346), .A3(new_n355), .ZN(new_n356));
  AOI211_X1 g155(.A(new_n330), .B(new_n342), .C1(new_n336), .C2(new_n337), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n354), .B1(new_n357), .B2(new_n353), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT27), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT67), .B1(new_n361), .B2(G183gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT67), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(new_n336), .A3(KEYINPUT27), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n364), .A3(new_n337), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(KEYINPUT68), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT68), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT27), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n336), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n360), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n336), .A2(KEYINPUT27), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n361), .A2(G183gat), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT28), .A4(new_n337), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n351), .A2(new_n352), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT26), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n347), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT69), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n347), .B2(new_n376), .ZN(new_n379));
  OAI211_X1 g178(.A(KEYINPUT69), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n377), .A2(new_n381), .B1(G183gat), .B2(G190gat), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n374), .A2(KEYINPUT70), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT70), .B1(new_n374), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n359), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G226gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n356), .A2(new_n358), .B1(new_n374), .B2(new_n382), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n386), .B1(new_n389), .B2(KEYINPUT29), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n390), .A3(KEYINPUT77), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n385), .A2(new_n392), .A3(new_n387), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n294), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(new_n387), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT70), .ZN(new_n396));
  INV_X1    g195(.A(new_n373), .ZN(new_n397));
  AOI21_X1  g196(.A(G190gat), .B1(new_n371), .B2(KEYINPUT67), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n398), .B(new_n364), .C1(new_n336), .C2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n400), .B2(new_n360), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n377), .A2(new_n381), .ZN(new_n402));
  NAND2_X1  g201(.A1(G183gat), .A2(G190gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n396), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n374), .A2(KEYINPUT70), .A3(new_n382), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n405), .A2(new_n406), .B1(new_n358), .B2(new_n356), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n387), .A2(KEYINPUT29), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n395), .B(new_n294), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n328), .B1(new_n394), .B2(new_n411), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n407), .A2(KEYINPUT77), .A3(new_n386), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n392), .B1(new_n385), .B2(new_n387), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n390), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n410), .B(new_n327), .C1(new_n415), .C2(new_n294), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n412), .A2(new_n416), .A3(KEYINPUT30), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n391), .A2(new_n393), .ZN(new_n418));
  INV_X1    g217(.A(new_n294), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n411), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n327), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n324), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT75), .ZN(new_n424));
  INV_X1    g223(.A(new_n220), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n385), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G227gat), .A2(G233gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n405), .A2(new_n406), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(new_n220), .A3(new_n359), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G15gat), .B(G43gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(G71gat), .B(G99gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(KEYINPUT32), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT73), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT73), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n431), .A2(new_n439), .A3(KEYINPUT32), .A4(new_n436), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n431), .A2(new_n435), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n434), .B1(new_n431), .B2(KEYINPUT32), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n438), .A2(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n430), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n220), .B1(new_n429), .B2(new_n359), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n427), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT34), .B1(new_n446), .B2(KEYINPUT74), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n428), .B1(new_n426), .B2(new_n430), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT74), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT34), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n424), .B1(new_n443), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n440), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n442), .A2(new_n441), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n443), .A2(KEYINPUT75), .A3(new_n452), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n280), .B(new_n423), .C1(new_n457), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n318), .A2(new_n322), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n443), .B2(new_n452), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n454), .A2(new_n455), .ZN(new_n463));
  OR2_X1    g262(.A1(new_n447), .A2(new_n451), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n417), .A2(new_n422), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n276), .A2(new_n277), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n270), .B1(new_n468), .B2(new_n273), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT35), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n460), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n443), .A2(new_n452), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n465), .A2(new_n424), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n458), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(KEYINPUT36), .A3(new_n473), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n461), .B(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n410), .B1(new_n415), .B2(new_n294), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n328), .B1(new_n482), .B2(KEYINPUT37), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n418), .A2(new_n294), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT37), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n385), .A2(new_n408), .B1(new_n387), .B2(new_n389), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n486), .B2(new_n419), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT88), .B(KEYINPUT38), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n416), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n327), .B1(new_n420), .B2(new_n485), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n482), .A2(KEYINPUT37), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n491), .A2(new_n494), .A3(new_n280), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n272), .A2(new_n278), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n240), .A2(new_n249), .A3(new_n251), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(new_n261), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n497), .A3(new_n261), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n260), .A2(new_n261), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n500), .A2(KEYINPUT39), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT39), .ZN(new_n504));
  INV_X1    g303(.A(new_n501), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(new_n499), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n506), .A3(new_n278), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n496), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n503), .A2(new_n506), .A3(KEYINPUT40), .A4(new_n278), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n509), .A2(new_n417), .A3(new_n422), .A4(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n461), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n481), .B1(new_n495), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n472), .B1(new_n478), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT90), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n476), .A2(new_n477), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n511), .A2(new_n512), .ZN(new_n519));
  INV_X1    g318(.A(new_n494), .ZN(new_n520));
  INV_X1    g319(.A(new_n280), .ZN(new_n521));
  INV_X1    g320(.A(new_n489), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n484), .B2(new_n487), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n492), .A2(new_n523), .B1(new_n420), .B2(new_n327), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n518), .A2(new_n526), .A3(new_n481), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(KEYINPUT90), .A3(new_n472), .ZN(new_n528));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529));
  INV_X1    g328(.A(G1gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(KEYINPUT93), .A3(KEYINPUT16), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT16), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(G1gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n529), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  OAI221_X1 g334(.A(new_n535), .B1(KEYINPUT94), .B2(G8gat), .C1(new_n530), .C2(new_n529), .ZN(new_n536));
  NAND2_X1  g335(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n536), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G43gat), .B(G50gat), .ZN(new_n540));
  INV_X1    g339(.A(G29gat), .ZN(new_n541));
  INV_X1    g340(.A(G36gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT14), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT14), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(G29gat), .B2(G36gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n546), .A2(new_n547), .B1(new_n541), .B2(new_n542), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT92), .B1(new_n543), .B2(new_n545), .ZN(new_n549));
  OAI211_X1 g348(.A(KEYINPUT15), .B(new_n540), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n540), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n551));
  INV_X1    g350(.A(new_n546), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n551), .B(new_n552), .C1(KEYINPUT15), .C2(new_n540), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(KEYINPUT17), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(new_n550), .B2(new_n553), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n539), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT95), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT95), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n560), .B(new_n539), .C1(new_n555), .C2(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n536), .B(new_n537), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT96), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n539), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n554), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT18), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(G229gat), .B2(G233gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n562), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT97), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n559), .A2(new_n561), .B1(new_n567), .B2(new_n554), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n574), .A3(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G229gat), .A2(G233gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n577), .A3(new_n568), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n564), .A2(new_n566), .A3(new_n550), .A4(new_n553), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n568), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n577), .B(KEYINPUT13), .Z(new_n581));
  AOI22_X1  g380(.A1(new_n578), .A2(new_n569), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n578), .B2(new_n569), .ZN(new_n585));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(G169gat), .B(G197gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT12), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n583), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n576), .B(new_n582), .C1(new_n585), .C2(new_n592), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT99), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT99), .B1(new_n594), .B2(new_n595), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT100), .ZN(new_n600));
  XNOR2_X1  g399(.A(G57gat), .B(G64gat), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G71gat), .B(G78gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n607));
  AND2_X1   g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G127gat), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n567), .B1(KEYINPUT21), .B2(new_n606), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G155gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n612), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  INV_X1    g419(.A(G92gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT7), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n622), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G99gat), .B(G106gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(G99gat), .A2(G106gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(KEYINPUT8), .A2(new_n627), .B1(new_n620), .B2(new_n621), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n626), .B1(new_n625), .B2(new_n628), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n631), .A2(new_n554), .B1(KEYINPUT41), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n555), .A2(new_n557), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n631), .ZN(new_n635));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n638));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n637), .B(new_n640), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n631), .A2(new_n606), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n605), .B1(new_n629), .B2(new_n630), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n631), .A2(new_n606), .A3(KEYINPUT10), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n643), .A2(new_n645), .ZN(new_n655));
  INV_X1    g454(.A(new_n649), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n650), .A2(new_n659), .ZN(new_n662));
  AOI22_X1  g461(.A1(new_n661), .A2(new_n662), .B1(new_n655), .B2(new_n656), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n658), .B1(new_n663), .B2(new_n653), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n619), .A2(new_n642), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n517), .A2(new_n528), .A3(new_n599), .A4(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT103), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(KEYINPUT103), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n469), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n469), .A2(new_n672), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  INV_X1    g476(.A(new_n467), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT105), .B(KEYINPUT16), .ZN(new_n679));
  INV_X1    g478(.A(G8gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n671), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n680), .B1(new_n671), .B2(new_n678), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(KEYINPUT42), .B2(new_n682), .ZN(G1325gat));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n474), .A2(new_n458), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n518), .B1(new_n669), .B2(new_n670), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n689), .B2(new_n686), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n671), .A2(new_n480), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(new_n619), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n641), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n664), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n517), .A2(new_n528), .A3(new_n599), .A4(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n675), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n697), .A2(G29gat), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT45), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n619), .B(KEYINPUT106), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n594), .A2(new_n595), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n703), .A3(new_n665), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n517), .A2(new_n528), .A3(new_n641), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT44), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n460), .A2(new_n707), .A3(new_n471), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n460), .B2(new_n471), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n527), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n527), .B(KEYINPUT108), .C1(new_n708), .C2(new_n709), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n642), .A2(KEYINPUT44), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n704), .B1(new_n706), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n698), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n718), .ZN(G1328gat));
  NAND2_X1  g518(.A1(new_n678), .A2(new_n542), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n697), .A2(KEYINPUT46), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT110), .Z(new_n722));
  OAI21_X1  g521(.A(KEYINPUT46), .B1(new_n697), .B2(new_n720), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT109), .ZN(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n717), .B2(new_n467), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(G1329gat));
  NAND3_X1  g525(.A1(new_n716), .A2(G43gat), .A3(new_n478), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n697), .B1(new_n458), .B2(new_n474), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(G43gat), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n706), .A2(new_n715), .ZN(new_n732));
  INV_X1    g531(.A(new_n704), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n461), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G50gat), .ZN(new_n735));
  INV_X1    g534(.A(G50gat), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n736), .B(new_n480), .C1(new_n697), .C2(KEYINPUT111), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n697), .A2(KEYINPUT111), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n731), .B1(new_n735), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n736), .B1(new_n716), .B2(new_n480), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n731), .B1(new_n737), .B2(new_n738), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT112), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n742), .A2(new_n743), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n736), .B1(new_n716), .B2(new_n461), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT48), .B1(new_n747), .B2(new_n739), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n745), .A2(new_n750), .ZN(G1331gat));
  AND2_X1   g550(.A1(new_n712), .A2(new_n713), .ZN(new_n752));
  INV_X1    g551(.A(new_n703), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n664), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n754), .A2(new_n694), .A3(new_n641), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n675), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g558(.A(new_n467), .B(KEYINPUT113), .Z(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n763), .B(new_n764), .Z(G1333gat));
  OAI21_X1  g564(.A(G71gat), .B1(new_n756), .B2(new_n518), .ZN(new_n766));
  INV_X1    g565(.A(G71gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n687), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n756), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g569(.A1(new_n757), .A2(new_n480), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n754), .A2(new_n619), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n732), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774), .B2(new_n698), .ZN(new_n775));
  INV_X1    g574(.A(new_n695), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n710), .A2(new_n753), .A3(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(KEYINPUT51), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(KEYINPUT51), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n778), .A2(new_n779), .A3(new_n665), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n620), .A3(new_n675), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n775), .A2(new_n781), .ZN(G1336gat));
  NOR2_X1   g581(.A1(new_n761), .A2(G92gat), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT52), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G92gat), .B1(new_n774), .B2(new_n761), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n774), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n678), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n788), .A2(G92gat), .B1(new_n780), .B2(new_n783), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(G1337gat));
  AND3_X1   g590(.A1(new_n787), .A2(G99gat), .A3(new_n478), .ZN(new_n792));
  AOI21_X1  g591(.A(G99gat), .B1(new_n780), .B2(new_n687), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(G1338gat));
  NOR2_X1   g593(.A1(new_n512), .A2(G106gat), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT53), .B1(new_n780), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G106gat), .B1(new_n774), .B2(new_n512), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n787), .A2(new_n480), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n799), .A2(G106gat), .B1(new_n780), .B2(new_n795), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(G1339gat));
  NOR2_X1   g601(.A1(new_n666), .A2(new_n703), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n577), .A2(new_n573), .B1(new_n580), .B2(new_n581), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n590), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT115), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n576), .A2(new_n592), .A3(new_n582), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n664), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n662), .ZN(new_n809));
  XNOR2_X1  g608(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n809), .A2(new_n660), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n646), .A2(new_n656), .A3(new_n647), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n654), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n811), .A2(new_n815), .A3(KEYINPUT55), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n809), .A2(new_n660), .A3(new_n810), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n814), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n658), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n808), .B1(new_n753), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n642), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n806), .B2(new_n807), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n806), .A2(new_n823), .A3(new_n807), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n820), .A2(new_n642), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n803), .B1(new_n829), .B2(new_n702), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n480), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n698), .A2(new_n760), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n687), .A3(new_n832), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n833), .A2(new_n206), .A3(new_n598), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n830), .A2(new_n698), .ZN(new_n835));
  INV_X1    g634(.A(new_n466), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n760), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n703), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n834), .B1(new_n839), .B2(new_n206), .ZN(G1340gat));
  NOR3_X1   g639(.A1(new_n833), .A2(new_n204), .A3(new_n665), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n664), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n204), .ZN(G1341gat));
  INV_X1    g642(.A(G127gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n838), .A2(new_n844), .A3(new_n619), .ZN(new_n845));
  OAI21_X1  g644(.A(G127gat), .B1(new_n833), .B2(new_n702), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT117), .ZN(G1342gat));
  OR4_X1    g647(.A1(G134gat), .A2(new_n837), .A3(new_n678), .A4(new_n642), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n850));
  OAI21_X1  g649(.A(G134gat), .B1(new_n833), .B2(new_n642), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(G1343gat));
  NAND2_X1  g652(.A1(new_n832), .A2(new_n518), .ZN(new_n854));
  INV_X1    g653(.A(new_n820), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n596), .B2(new_n597), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n641), .B1(new_n856), .B2(new_n808), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n827), .A2(new_n826), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n824), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n694), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n703), .B2(new_n666), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(KEYINPUT57), .A3(new_n480), .ZN(new_n862));
  XNOR2_X1  g661(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n830), .B2(new_n512), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n854), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n221), .B1(new_n865), .B2(new_n703), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n478), .A2(new_n512), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n835), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n760), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n598), .A2(G141gat), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n870), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n872), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n221), .B1(new_n865), .B2(new_n599), .ZN(new_n875));
  OAI22_X1  g674(.A1(new_n871), .A2(new_n872), .B1(new_n874), .B2(new_n875), .ZN(G1344gat));
  NAND3_X1  g675(.A1(new_n869), .A2(new_n222), .A3(new_n664), .ZN(new_n877));
  AOI211_X1 g676(.A(KEYINPUT59), .B(new_n222), .C1(new_n865), .C2(new_n664), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  INV_X1    g678(.A(new_n863), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n701), .B1(new_n822), .B2(new_n828), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n461), .B(new_n880), .C1(new_n881), .C2(new_n803), .ZN(new_n882));
  INV_X1    g681(.A(new_n480), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n667), .A2(new_n598), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n860), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n885), .B2(KEYINPUT57), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n886), .A2(new_n518), .A3(new_n664), .A4(new_n832), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n879), .B1(new_n887), .B2(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n877), .B1(new_n878), .B2(new_n888), .ZN(G1345gat));
  INV_X1    g688(.A(new_n865), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n242), .B1(new_n890), .B2(new_n702), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n869), .A2(new_n230), .A3(new_n231), .A4(new_n619), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1346gat));
  OAI21_X1  g692(.A(G162gat), .B1(new_n890), .B2(new_n642), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n641), .A2(new_n467), .A3(new_n229), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n868), .B2(new_n895), .ZN(G1347gat));
  NAND2_X1  g695(.A1(new_n760), .A2(new_n836), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT120), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT119), .B1(new_n830), .B2(new_n675), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(new_n698), .C1(new_n881), .C2(new_n803), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n898), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n703), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n675), .A2(new_n467), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n831), .A2(new_n687), .A3(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(new_n351), .A3(new_n598), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n903), .A2(new_n906), .ZN(G1348gat));
  NAND3_X1  g706(.A1(new_n902), .A2(new_n352), .A3(new_n664), .ZN(new_n908));
  OAI21_X1  g707(.A(G176gat), .B1(new_n905), .B2(new_n665), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1349gat));
  OAI21_X1  g709(.A(G183gat), .B1(new_n905), .B2(new_n702), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n619), .A2(new_n371), .A3(new_n372), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n902), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n902), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT60), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n918), .B(new_n911), .C1(new_n914), .C2(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n905), .B2(new_n642), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n921), .A2(KEYINPUT122), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(KEYINPUT122), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(KEYINPUT61), .A3(new_n923), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n923), .A2(KEYINPUT61), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n902), .A2(new_n337), .A3(new_n641), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(G1351gat));
  NAND2_X1  g726(.A1(new_n899), .A2(new_n901), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n867), .A2(new_n760), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  OR3_X1    g730(.A1(new_n931), .A2(G197gat), .A3(new_n753), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n904), .A2(new_n518), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT123), .Z(new_n934));
  AND2_X1   g733(.A1(new_n886), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n599), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT124), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G197gat), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n936), .A2(KEYINPUT124), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n932), .B1(new_n938), .B2(new_n939), .ZN(G1352gat));
  NAND2_X1  g739(.A1(new_n935), .A2(new_n664), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G204gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n665), .A2(G204gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n930), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT62), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n928), .A2(new_n947), .A3(new_n930), .A4(new_n944), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n942), .A2(new_n943), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n946), .A2(new_n948), .ZN(new_n950));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n951), .B1(new_n935), .B2(new_n664), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT125), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n949), .A2(new_n953), .ZN(G1353gat));
  OR3_X1    g753(.A1(new_n931), .A2(G211gat), .A3(new_n694), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n886), .A2(KEYINPUT126), .A3(new_n619), .A4(new_n934), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n956), .A2(G211gat), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n886), .A2(new_n619), .A3(new_n934), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  AND4_X1   g760(.A1(KEYINPUT63), .A2(new_n960), .A3(G211gat), .A4(new_n956), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n955), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  INV_X1    g762(.A(G218gat), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n928), .A2(new_n964), .A3(new_n641), .A4(new_n930), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n935), .A2(new_n641), .ZN(new_n966));
  OAI211_X1 g765(.A(KEYINPUT127), .B(new_n965), .C1(new_n966), .C2(new_n964), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n964), .B1(new_n935), .B2(new_n641), .ZN(new_n969));
  INV_X1    g768(.A(new_n965), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n967), .A2(new_n971), .ZN(G1355gat));
endmodule


