//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND3_X1  g0009(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n203), .A2(G50), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT66), .B(G244), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G77), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G97), .A2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT65), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n209), .B1(new_n210), .B2(new_n212), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT2), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XOR2_X1   g0028(.A(G250), .B(G257), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT67), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n228), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XNOR2_X1  g0034(.A(G50), .B(G58), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(KEYINPUT74), .ZN(new_n241));
  INV_X1    g0041(.A(G41), .ZN(new_n242));
  INV_X1    g0042(.A(G45), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT68), .ZN(new_n245));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  NAND4_X1  g0046(.A1(new_n244), .A2(new_n245), .A3(new_n246), .A4(G274), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(G274), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G41), .A2(G45), .ZN(new_n249));
  OAI21_X1  g0049(.A(KEYINPUT68), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  OAI211_X1 g0053(.A(G1), .B(G13), .C1(new_n253), .C2(new_n242), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT69), .B(G1), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n244), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n252), .B1(new_n257), .B2(G226), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  OAI21_X1  g0061(.A(KEYINPUT70), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n253), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT70), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT71), .B(G1698), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G222), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G77), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G223), .ZN(new_n273));
  OAI221_X1 g0073(.A(new_n270), .B1(new_n271), .B2(new_n268), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n259), .B1(new_n274), .B2(new_n255), .ZN(new_n275));
  INV_X1    g0075(.A(G200), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n241), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(G190), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G1), .A2(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n282));
  INV_X1    g0082(.A(G150), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(G20), .A3(new_n253), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n281), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n246), .A2(KEYINPUT69), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT69), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G1), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n290), .A2(new_n292), .A3(G13), .A4(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G50), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n256), .A2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n281), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n297), .A2(G50), .A3(new_n298), .A4(new_n293), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n289), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n300), .A2(KEYINPUT9), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(KEYINPUT9), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT10), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n277), .A2(new_n278), .A3(new_n303), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n275), .A2(new_n241), .A3(new_n276), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT75), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n278), .A2(new_n303), .ZN(new_n307));
  INV_X1    g0107(.A(new_n305), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT75), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .A4(new_n277), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n301), .A2(new_n302), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n278), .B(new_n311), .C1(new_n276), .C2(new_n275), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n306), .A2(new_n310), .B1(KEYINPUT10), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n275), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(G179), .B2(new_n275), .ZN(new_n316));
  INV_X1    g0116(.A(new_n300), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n262), .A2(new_n267), .A3(G226), .A4(new_n269), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n262), .A2(new_n267), .A3(G232), .A4(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n255), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n290), .A2(new_n292), .ZN(new_n326));
  OAI211_X1 g0126(.A(G238), .B(new_n254), .C1(new_n326), .C2(new_n249), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n251), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n320), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  AOI211_X1 g0130(.A(KEYINPUT13), .B(new_n328), .C1(new_n324), .C2(new_n255), .ZN(new_n331));
  OAI21_X1  g0131(.A(G169), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT14), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n334), .B(G169), .C1(new_n330), .C2(new_n331), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n330), .A2(new_n331), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G179), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G20), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n285), .A2(new_n295), .B1(new_n339), .B2(G68), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n253), .A2(new_n271), .A3(G20), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n281), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT11), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n293), .A2(new_n298), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(G68), .A3(new_n297), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n342), .A2(new_n343), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n344), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n293), .A2(G68), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT12), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n338), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT18), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G58), .A2(G68), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n339), .B1(new_n203), .B2(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n284), .A2(KEYINPUT76), .A3(G159), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT76), .B1(new_n284), .B2(G159), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n262), .A2(new_n267), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT7), .B1(new_n361), .B2(new_n339), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n260), .A2(new_n261), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n363), .A2(KEYINPUT7), .A3(new_n339), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n360), .B1(new_n365), .B2(new_n202), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT16), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT7), .B1(new_n363), .B2(new_n339), .ZN(new_n369));
  OAI21_X1  g0169(.A(G68), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(KEYINPUT16), .A3(new_n360), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n371), .A2(new_n281), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n287), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n297), .A2(new_n374), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n375), .A2(KEYINPUT77), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n345), .B1(new_n375), .B2(KEYINPUT77), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n376), .A2(new_n377), .B1(new_n287), .B2(new_n294), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n269), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n380));
  INV_X1    g0180(.A(G87), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n380), .A2(new_n363), .B1(new_n253), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n255), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n252), .B1(new_n257), .B2(G232), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n314), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(G179), .B2(new_n385), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n355), .B1(new_n379), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n378), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n368), .B2(new_n372), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n391), .A2(KEYINPUT18), .A3(new_n387), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n385), .A2(KEYINPUT78), .A3(G190), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n385), .A2(G190), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT78), .B1(new_n385), .B2(new_n276), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT17), .B1(new_n398), .B2(new_n391), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n397), .ZN(new_n401));
  INV_X1    g0201(.A(new_n396), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n394), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n379), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT17), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n393), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n268), .A2(G232), .A3(new_n269), .ZN(new_n408));
  INV_X1    g0208(.A(G107), .ZN(new_n409));
  INV_X1    g0209(.A(G238), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n408), .B1(new_n409), .B2(new_n268), .C1(new_n272), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n255), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n252), .B1(new_n257), .B2(new_n214), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(G179), .A3(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n314), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT15), .B(G87), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT72), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(new_n339), .A3(G33), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n374), .A2(new_n284), .B1(G20), .B2(G77), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n298), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n346), .A2(G77), .A3(new_n297), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT73), .B1(new_n293), .B2(G77), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n293), .A2(KEYINPUT73), .A3(G77), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n416), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n336), .A2(G200), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n330), .A2(new_n331), .A3(G190), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n352), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G190), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n412), .A2(new_n435), .A3(new_n413), .ZN(new_n436));
  AOI21_X1  g0236(.A(G200), .B1(new_n412), .B2(new_n413), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n428), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n431), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  AND4_X1   g0239(.A1(new_n319), .A2(new_n354), .A3(new_n407), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT88), .ZN(new_n442));
  INV_X1    g0242(.A(G1698), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT71), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT71), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G1698), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n446), .A3(G250), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G257), .A2(G1698), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n363), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G294), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n253), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n255), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  AND2_X1   g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n256), .B(G45), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(G264), .A3(new_n254), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n290), .A2(new_n292), .A3(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n454), .A2(new_n453), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(G274), .A3(new_n254), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n452), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G179), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(G169), .B2(new_n461), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT87), .ZN(new_n466));
  OR3_X1    g0266(.A1(new_n339), .A2(KEYINPUT23), .A3(G107), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n339), .A2(G33), .A3(G116), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT23), .B1(new_n339), .B2(G107), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n381), .A2(KEYINPUT22), .A3(G20), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n262), .A2(new_n267), .A3(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n339), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT22), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n473), .A2(new_n475), .A3(KEYINPUT86), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT86), .B1(new_n473), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n466), .B1(new_n478), .B2(KEYINPUT24), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT24), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(new_n471), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(new_n466), .A3(KEYINPUT24), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n298), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n345), .B1(G33), .B2(new_n256), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G107), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT25), .B1(new_n293), .B2(G107), .ZN(new_n488));
  OR3_X1    g0288(.A1(new_n293), .A2(KEYINPUT25), .A3(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n442), .B(new_n465), .C1(new_n485), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n473), .A2(new_n475), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT86), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n473), .A2(new_n475), .A3(KEYINPUT86), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n470), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT87), .B1(new_n496), .B2(new_n480), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(new_n484), .A3(new_n481), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n490), .B1(new_n498), .B2(new_n281), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT88), .B1(new_n499), .B2(new_n464), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n461), .A2(new_n276), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(G190), .B2(new_n461), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n491), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n290), .A2(new_n292), .A3(G33), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n293), .A2(new_n298), .A3(new_n505), .A4(G116), .ZN(new_n506));
  INV_X1    g0306(.A(G116), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n256), .A2(G13), .A3(G20), .A4(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT20), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n339), .A2(new_n507), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  INV_X1    g0312(.A(G97), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(G33), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n511), .B1(new_n514), .B2(new_n339), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n510), .B1(new_n515), .B2(new_n298), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n253), .A2(G97), .ZN(new_n517));
  AOI21_X1  g0317(.A(G20), .B1(new_n517), .B2(new_n512), .ZN(new_n518));
  OAI211_X1 g0318(.A(KEYINPUT20), .B(new_n281), .C1(new_n518), .C2(new_n511), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n509), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G303), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n262), .B2(new_n267), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n444), .A2(new_n446), .A3(G257), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G264), .A2(G1698), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n363), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n255), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(G270), .B(new_n254), .C1(new_n457), .C2(new_n458), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n455), .A2(KEYINPUT83), .A3(G270), .A4(new_n254), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n527), .A2(new_n460), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n532), .A2(new_n276), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(G190), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n521), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT85), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n314), .B1(new_n509), .B2(new_n520), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(KEYINPUT21), .A3(new_n532), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT84), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n538), .A2(new_n532), .A3(KEYINPUT84), .A4(KEYINPUT21), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n521), .A2(new_n532), .A3(new_n462), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT21), .B1(new_n538), .B2(new_n532), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(KEYINPUT85), .B(new_n521), .C1(new_n533), .C2(new_n534), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n537), .A2(new_n543), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n460), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n459), .A2(new_n255), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(G257), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(KEYINPUT4), .A2(G244), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n262), .A2(new_n267), .A3(new_n269), .A4(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT4), .ZN(new_n554));
  OAI21_X1  g0354(.A(G244), .B1(new_n260), .B2(new_n261), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n444), .A2(new_n446), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n557), .A3(new_n512), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n262), .A2(new_n267), .A3(G250), .A4(G1698), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n559), .A2(KEYINPUT79), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(KEYINPUT79), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n551), .B(G179), .C1(new_n562), .C2(new_n254), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n550), .A2(G257), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n460), .ZN(new_n565));
  INV_X1    g0365(.A(new_n558), .ZN(new_n566));
  INV_X1    g0366(.A(new_n561), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n559), .A2(KEYINPUT79), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n565), .B1(new_n569), .B2(new_n255), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n563), .B1(new_n570), .B2(new_n314), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT6), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n513), .A2(new_n409), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n409), .A2(KEYINPUT6), .A3(G97), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n365), .B2(new_n409), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n281), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n486), .A2(G97), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n294), .A2(new_n513), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n571), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n264), .A2(new_n266), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(new_n339), .A3(G68), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n339), .B1(new_n323), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n381), .A2(new_n513), .A3(new_n409), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n588), .B1(new_n323), .B2(G20), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n587), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n593), .A2(new_n281), .B1(new_n418), .B2(new_n294), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n486), .A2(new_n419), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n556), .A2(new_n363), .A3(new_n410), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n555), .A2(new_n443), .B1(new_n253), .B2(new_n507), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n255), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT81), .ZN(new_n600));
  AOI21_X1  g0400(.A(G274), .B1(new_n600), .B2(G250), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n457), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(KEYINPUT81), .A2(G250), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n256), .B2(G45), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n254), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G169), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n599), .A2(G179), .A3(new_n605), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n276), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n599), .A2(new_n435), .A3(new_n605), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n486), .A2(G87), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n594), .A2(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n596), .A2(new_n609), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n551), .B1(new_n562), .B2(new_n254), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT80), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n551), .B(KEYINPUT80), .C1(new_n562), .C2(new_n254), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n276), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n580), .B(new_n583), .C1(new_n616), .C2(new_n435), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n585), .B(new_n615), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n548), .B1(new_n622), .B2(KEYINPUT82), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n609), .A2(new_n596), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n612), .A2(new_n614), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n584), .B2(new_n571), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT82), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n627), .B(new_n628), .C1(new_n620), .C2(new_n621), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n441), .A2(new_n504), .A3(new_n630), .ZN(G372));
  AND3_X1   g0431(.A1(new_n398), .A2(KEYINPUT17), .A3(new_n391), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(new_n399), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n332), .A2(KEYINPUT14), .B1(new_n336), .B2(G179), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n352), .B1(new_n635), .B2(new_n335), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n430), .B2(new_n434), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n393), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n306), .A2(new_n310), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n318), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n498), .A2(new_n281), .ZN(new_n643));
  INV_X1    g0443(.A(new_n490), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n643), .A2(new_n644), .A3(new_n502), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n622), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT89), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n543), .A2(new_n647), .A3(new_n546), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(new_n543), .B2(new_n546), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n648), .A2(new_n649), .B1(new_n499), .B2(new_n464), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n646), .A2(KEYINPUT90), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n585), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(KEYINPUT26), .A3(new_n615), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n615), .A2(new_n584), .A3(new_n571), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n654), .A2(KEYINPUT91), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT91), .B1(new_n654), .B2(new_n655), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n651), .A2(new_n658), .A3(new_n624), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT90), .B1(new_n646), .B2(new_n650), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n642), .B1(new_n441), .B2(new_n661), .ZN(G369));
  OAI21_X1  g0462(.A(new_n465), .B1(new_n485), .B2(new_n490), .ZN(new_n663));
  INV_X1    g0463(.A(G13), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G20), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n256), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n663), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n671), .B1(new_n485), .B2(new_n490), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT92), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n504), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n543), .A2(new_n546), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n671), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n672), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n671), .ZN(new_n679));
  OAI22_X1  g0479(.A1(new_n674), .A2(new_n504), .B1(new_n663), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n548), .B1(new_n521), .B2(new_n679), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n679), .A2(new_n521), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n648), .B2(new_n649), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n678), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n207), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G1), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n381), .A2(new_n513), .A3(new_n409), .A4(new_n507), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n692), .A2(new_n693), .B1(new_n211), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n491), .A2(new_n500), .A3(new_n503), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(new_n629), .A3(new_n623), .A4(new_n679), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT30), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n532), .A2(new_n462), .ZN(new_n699));
  AND4_X1   g0499(.A1(new_n456), .A2(new_n599), .A3(new_n452), .A4(new_n605), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n698), .B1(new_n701), .B2(new_n616), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n570), .A2(KEYINPUT30), .A3(new_n699), .A4(new_n700), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n606), .A2(new_n461), .A3(new_n462), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n616), .A2(new_n704), .A3(new_n532), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT31), .B1(new_n706), .B2(new_n671), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n671), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n685), .B1(new_n697), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n679), .B1(new_n659), .B2(new_n660), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n654), .A2(new_n655), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n653), .A2(new_n715), .B1(new_n596), .B2(new_n609), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n491), .A2(new_n500), .A3(new_n676), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n717), .A2(new_n646), .A3(KEYINPUT93), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT93), .B1(new_n717), .B2(new_n646), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(KEYINPUT29), .A3(new_n679), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n711), .B1(new_n714), .B2(new_n721), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n722), .A2(KEYINPUT94), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(KEYINPUT94), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n695), .B1(new_n725), .B2(G1), .ZN(G364));
  AOI21_X1  g0526(.A(new_n692), .B1(G45), .B2(new_n665), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n268), .A2(G355), .A3(new_n207), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G116), .B2(new_n207), .ZN(new_n729));
  MUX2_X1   g0529(.A(new_n212), .B(new_n236), .S(G45), .Z(new_n730));
  NOR2_X1   g0530(.A1(new_n689), .A2(new_n586), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n280), .B1(G20), .B2(new_n314), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n727), .B1(new_n732), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT95), .ZN(new_n740));
  INV_X1    g0540(.A(new_n736), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n339), .A2(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n743), .A2(new_n462), .A3(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n462), .A2(new_n276), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n742), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT33), .B(G317), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n744), .A2(G311), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n339), .A2(new_n435), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(G179), .A3(new_n276), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n276), .A2(G179), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n752), .A2(G322), .B1(new_n755), .B2(G303), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n749), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n339), .B1(new_n758), .B2(G190), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n268), .B(new_n757), .C1(G294), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n742), .A2(new_n753), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n742), .A2(new_n758), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(G283), .A2(new_n763), .B1(new_n765), .B2(G329), .ZN(new_n766));
  INV_X1    g0566(.A(G326), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n745), .A2(new_n750), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n761), .B(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n752), .A2(G58), .B1(new_n763), .B2(G107), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n295), .B2(new_n768), .ZN(new_n771));
  INV_X1    g0571(.A(new_n744), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n772), .A2(KEYINPUT96), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(KEYINPUT96), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n771), .B1(new_n776), .B2(G77), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n760), .A2(G97), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n202), .A2(new_n746), .B1(new_n754), .B2(new_n381), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n361), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n764), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n777), .A2(new_n778), .A3(new_n780), .A4(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n769), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n740), .B1(new_n741), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT97), .Z(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n684), .B2(new_n735), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n686), .A2(new_n727), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n684), .A2(new_n685), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  NAND2_X1  g0592(.A1(new_n429), .A2(new_n671), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n438), .A2(new_n793), .B1(new_n416), .B2(new_n429), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n416), .A2(new_n429), .A3(new_n679), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(KEYINPUT101), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT101), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n438), .A2(new_n793), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n795), .C1(new_n799), .C2(new_n430), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n712), .B(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n727), .B1(new_n802), .B2(new_n711), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n711), .B2(new_n802), .ZN(new_n804));
  INV_X1    g0604(.A(new_n727), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n736), .A2(new_n733), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(new_n271), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT98), .ZN(new_n808));
  INV_X1    g0608(.A(new_n768), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G137), .A2(new_n809), .B1(new_n747), .B2(G150), .ZN(new_n810));
  INV_X1    g0610(.A(G143), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n810), .B1(new_n811), .B2(new_n751), .C1(new_n775), .C2(new_n781), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n760), .A2(G58), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n363), .B1(new_n765), .B2(G132), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n762), .A2(new_n202), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G50), .B2(new_n755), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n768), .A2(new_n522), .B1(new_n762), .B2(new_n381), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n778), .B1(new_n820), .B2(new_n746), .C1(new_n450), .C2(new_n751), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n819), .B(new_n821), .C1(G311), .C2(new_n765), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n361), .B1(new_n409), .B2(new_n754), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT99), .Z(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(new_n507), .C2(new_n775), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT100), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n741), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n808), .B1(new_n801), .B2(new_n734), .C1(new_n828), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n804), .A2(new_n831), .ZN(G384));
  NAND2_X1  g0632(.A1(new_n356), .A2(G77), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n211), .A2(new_n833), .B1(G50), .B2(new_n202), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n834), .A2(new_n664), .A3(new_n326), .ZN(new_n835));
  INV_X1    g0635(.A(new_n577), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT35), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n507), .B(new_n210), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT36), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT109), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n709), .B1(new_n707), .B2(KEYINPUT108), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT108), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n845), .B(KEYINPUT31), .C1(new_n706), .C2(new_n671), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n843), .B1(new_n697), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n697), .A2(new_n847), .A3(new_n843), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n440), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT110), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT104), .B1(new_n354), .B2(new_n679), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT104), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n636), .A2(new_n855), .A3(new_n671), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT103), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n354), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n636), .A2(KEYINPUT103), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n353), .A2(new_n671), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n434), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n857), .A2(new_n864), .A3(KEYINPUT105), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT105), .B1(new_n857), .B2(new_n864), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n801), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n850), .B2(new_n849), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT40), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n391), .A2(new_n387), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n391), .B2(new_n398), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  INV_X1    g0672(.A(new_n669), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n379), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n871), .A2(KEYINPUT107), .A3(new_n872), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n398), .A2(new_n391), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n379), .A2(new_n388), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n874), .A4(new_n872), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT107), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n876), .A2(new_n877), .A3(new_n874), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n875), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n874), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n406), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n370), .A2(new_n360), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n372), .B1(KEYINPUT16), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n378), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n873), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n406), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n387), .A2(new_n669), .B1(new_n890), .B2(new_n378), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n404), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n878), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n869), .B1(new_n888), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n797), .A2(new_n800), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT105), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n855), .B1(new_n636), .B2(new_n671), .ZN(new_n902));
  AND4_X1   g0702(.A1(new_n855), .A2(new_n338), .A3(new_n353), .A4(new_n671), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n338), .A2(KEYINPUT103), .A3(new_n353), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT103), .B1(new_n338), .B2(new_n353), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n905), .A2(new_n906), .A3(new_n862), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n901), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n857), .A2(new_n864), .A3(KEYINPUT105), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n900), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n892), .B1(new_n633), .B2(new_n393), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n896), .A2(new_n878), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n898), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n697), .A2(new_n847), .A3(new_n843), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n910), .B(new_n915), .C1(new_n916), .C2(new_n848), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n868), .A2(new_n899), .B1(new_n917), .B2(new_n869), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n853), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n853), .A2(new_n919), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(G330), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n393), .A2(new_n873), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n888), .A2(new_n924), .A3(new_n898), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n915), .A2(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n671), .B1(new_n859), .B2(new_n860), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n865), .A2(new_n866), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n801), .B(new_n679), .C1(new_n659), .C2(new_n660), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n795), .B(KEYINPUT102), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n915), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n714), .A2(new_n440), .A3(new_n721), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n642), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n935), .B(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n922), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT111), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n940), .B1(new_n256), .B2(new_n665), .C1(new_n922), .C2(new_n938), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n939), .A2(KEYINPUT111), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n842), .B1(new_n941), .B2(new_n942), .ZN(G367));
  INV_X1    g0743(.A(new_n731), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n232), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n737), .B1(new_n418), .B2(new_n207), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n776), .A2(G50), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n760), .A2(G68), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n746), .A2(new_n781), .B1(new_n762), .B2(new_n271), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n361), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n768), .A2(new_n811), .B1(new_n754), .B2(new_n201), .ZN(new_n951));
  INV_X1    g0751(.A(G137), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n751), .A2(new_n283), .B1(new_n764), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n947), .A2(new_n948), .A3(new_n950), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n755), .A2(G116), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT46), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n363), .B1(new_n450), .B2(new_n746), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n752), .A2(G303), .B1(new_n809), .B2(G311), .ZN(new_n959));
  INV_X1    g0759(.A(G317), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n959), .B1(new_n513), .B2(new_n762), .C1(new_n960), .C2(new_n764), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n958), .B(new_n961), .C1(new_n957), .C2(new_n956), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT113), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n776), .A2(G283), .B1(G107), .B2(new_n760), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n964), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(KEYINPUT113), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n955), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT47), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n736), .B1(new_n968), .B2(new_n969), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n727), .B1(new_n945), .B2(new_n946), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n626), .B1(new_n614), .B2(new_n679), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n614), .A2(new_n679), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n624), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n972), .B1(new_n735), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT114), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n246), .B1(new_n665), .B2(G45), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n687), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n584), .B1(new_n571), .B2(new_n671), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n620), .B2(new_n621), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n652), .A2(new_n671), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND3_X1   g0785(.A1(new_n678), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT45), .B1(new_n678), .B2(new_n985), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n675), .A2(new_n677), .ZN(new_n989));
  INV_X1    g0789(.A(new_n672), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT44), .ZN(new_n992));
  INV_X1    g0792(.A(new_n985), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(KEYINPUT44), .B1(new_n678), .B2(new_n985), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n981), .B1(new_n988), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n991), .B2(new_n993), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n678), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n1001), .A2(new_n687), .A3(new_n995), .A4(new_n994), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n680), .B(new_n686), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(new_n677), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n725), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n690), .B(KEYINPUT41), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n980), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n985), .B(KEYINPUT112), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n500), .B2(new_n491), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n679), .B1(new_n1013), .B2(new_n652), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n680), .A2(new_n677), .A3(new_n985), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT42), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(KEYINPUT42), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n976), .ZN(new_n1019));
  OR3_X1    g0819(.A1(new_n1018), .A2(KEYINPUT43), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n981), .A2(new_n1011), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1018), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1020), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  AND3_X1   g0827(.A1(new_n1018), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1024), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1021), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n978), .B1(new_n1010), .B2(new_n1031), .ZN(G387));
  AOI21_X1  g0832(.A(new_n1006), .B1(new_n723), .B2(new_n724), .ZN(new_n1033));
  OAI21_X1  g0833(.A(KEYINPUT116), .B1(new_n1033), .B2(new_n691), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n725), .A2(new_n1005), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT116), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n1036), .A3(new_n690), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1034), .B(new_n1037), .C1(new_n725), .C2(new_n1005), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n768), .A2(new_n781), .B1(new_n754), .B2(new_n271), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n363), .B(new_n1039), .C1(G97), .C2(new_n763), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n419), .A2(new_n760), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n752), .A2(G50), .B1(new_n765), .B2(G150), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n744), .A2(G68), .B1(new_n747), .B2(new_n374), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n586), .B1(new_n763), .B2(G116), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n754), .A2(new_n450), .B1(new_n759), .B2(new_n820), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n752), .A2(G317), .B1(new_n809), .B2(G322), .ZN(new_n1047));
  INV_X1    g0847(.A(G311), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1047), .B1(new_n1048), .B2(new_n746), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n776), .B2(G303), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1046), .B1(new_n1050), .B2(KEYINPUT48), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(KEYINPUT48), .B2(new_n1050), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1045), .B1(new_n767), .B2(new_n764), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1044), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n805), .B1(new_n1056), .B2(new_n736), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n374), .A2(new_n295), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT50), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n243), .B1(new_n202), .B2(new_n271), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1059), .A2(new_n693), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n731), .B1(new_n228), .B2(new_n243), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n268), .A2(new_n207), .A3(new_n693), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n207), .A2(G107), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n737), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n735), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1057), .B(new_n1066), .C1(new_n680), .C2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT115), .Z(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1005), .B2(new_n980), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1038), .A2(new_n1070), .ZN(G393));
  INV_X1    g0871(.A(new_n1003), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n691), .B1(new_n1033), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1035), .A2(new_n1003), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1012), .A2(new_n735), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n737), .B1(new_n513), .B2(new_n207), .C1(new_n239), .C2(new_n944), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n727), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n744), .A2(G294), .B1(G322), .B2(new_n765), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n522), .B2(new_n746), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n752), .A2(G311), .B1(new_n809), .B2(G317), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT118), .B(KEYINPUT52), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n754), .A2(new_n820), .B1(new_n762), .B2(new_n409), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n268), .B(new_n1084), .C1(G116), .C2(new_n760), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1083), .B(new_n1085), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n775), .A2(new_n287), .B1(new_n295), .B2(new_n746), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT117), .Z(new_n1088));
  OAI22_X1  g0888(.A1(new_n754), .A2(new_n202), .B1(new_n764), .B2(new_n811), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n363), .B(new_n1089), .C1(G87), .C2(new_n763), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n751), .A2(new_n781), .B1(new_n768), .B2(new_n283), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n759), .A2(new_n271), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1090), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1086), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1078), .B1(new_n1096), .B2(new_n736), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1076), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n1003), .B2(new_n979), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1075), .A2(new_n1100), .ZN(G390));
  OAI22_X1  g0901(.A1(new_n746), .A2(new_n952), .B1(new_n759), .B2(new_n781), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT54), .B(G143), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1102), .B1(new_n776), .B2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT119), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n752), .A2(G132), .B1(new_n765), .B2(G125), .ZN(new_n1107));
  INV_X1    g0907(.A(G128), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1107), .B1(new_n295), .B2(new_n762), .C1(new_n1108), .C2(new_n768), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n754), .A2(KEYINPUT53), .A3(new_n283), .ZN(new_n1110));
  OAI21_X1  g0910(.A(KEYINPUT53), .B1(new_n754), .B2(new_n283), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n268), .A2(new_n1111), .ZN(new_n1112));
  OR4_X1    g0912(.A1(new_n1106), .A2(new_n1109), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n776), .A2(G97), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n816), .B(new_n268), .C1(G87), .C2(new_n755), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n751), .A2(new_n507), .B1(new_n768), .B2(new_n820), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n746), .A2(new_n409), .B1(new_n764), .B2(new_n450), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1114), .A2(new_n1094), .A3(new_n1115), .A4(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n741), .B1(new_n1113), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n805), .B(new_n1120), .C1(new_n287), .C2(new_n806), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n927), .B2(new_n734), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n900), .A2(new_n685), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n908), .A2(new_n909), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(new_n916), .C2(new_n848), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n931), .A2(new_n932), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1124), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n928), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n927), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n720), .A2(new_n679), .A3(new_n801), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n930), .B1(new_n1131), .B2(new_n932), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n888), .A2(new_n898), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1129), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1126), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n924), .B1(new_n914), .B2(new_n898), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n912), .A2(new_n913), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n886), .A2(new_n887), .B1(new_n1138), .B2(KEYINPUT38), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1137), .B1(new_n1139), .B2(new_n924), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n933), .B2(new_n928), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n910), .A2(new_n711), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n1132), .C2(new_n1134), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1136), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1122), .B1(new_n1144), .B2(new_n979), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n711), .A2(new_n801), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n930), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1125), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1127), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1123), .B1(new_n916), .B2(new_n848), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n930), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1131), .A2(new_n932), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n1142), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1149), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n851), .A2(G330), .A3(new_n440), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n642), .A3(new_n936), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n691), .B1(new_n1144), .B2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1136), .A2(new_n1143), .A3(new_n1157), .A4(new_n1154), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1145), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(G378));
  INV_X1    g0962(.A(new_n935), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n318), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n317), .A2(new_n669), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n641), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n313), .B2(new_n318), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1165), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1165), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(KEYINPUT120), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT121), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1169), .A2(new_n1170), .A3(new_n1165), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(new_n1171), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT121), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n685), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1175), .B1(new_n918), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n917), .A2(new_n869), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n851), .A2(new_n899), .A3(new_n910), .ZN(new_n1182));
  AND4_X1   g0982(.A1(new_n1181), .A2(new_n1179), .A3(new_n1175), .A4(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1163), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1181), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1175), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1181), .A2(new_n1179), .A3(new_n1175), .A4(new_n1182), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n935), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1184), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT57), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1160), .A2(new_n1157), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1191), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n690), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1177), .A2(new_n733), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n736), .A2(G50), .A3(new_n733), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n586), .A2(G41), .ZN(new_n1198));
  AOI211_X1 g0998(.A(G50), .B(new_n1198), .C1(new_n253), .C2(new_n242), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n752), .A2(G107), .B1(new_n765), .B2(G283), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n513), .B2(new_n746), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G116), .A2(new_n809), .B1(new_n755), .B2(G77), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n763), .A2(G58), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1202), .A2(new_n948), .A3(new_n1198), .A4(new_n1203), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1201), .B(new_n1204), .C1(new_n419), .C2(new_n744), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1199), .B1(new_n1205), .B2(KEYINPUT58), .ZN(new_n1206));
  INV_X1    g1006(.A(G125), .ZN(new_n1207));
  INV_X1    g1007(.A(G132), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n768), .A2(new_n1207), .B1(new_n746), .B2(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n752), .A2(G128), .B1(new_n755), .B2(new_n1104), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n952), .B2(new_n772), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(G150), .C2(new_n760), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n253), .B(new_n242), .C1(new_n762), .C2(new_n781), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G124), .B2(new_n765), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT59), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1216), .B1(new_n1212), .B2(new_n1217), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1206), .B1(KEYINPUT58), .B2(new_n1205), .C1(new_n1214), .C2(new_n1218), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n805), .B(new_n1197), .C1(new_n1219), .C2(new_n736), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1190), .A2(new_n980), .B1(new_n1196), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1195), .A2(new_n1221), .ZN(G375));
  NAND3_X1  g1022(.A1(new_n1156), .A2(new_n1149), .A3(new_n1153), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1158), .A2(new_n1009), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n805), .B1(new_n202), .B2(new_n806), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n752), .A2(G137), .B1(new_n809), .B2(G132), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n586), .A3(new_n1203), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G159), .A2(new_n755), .B1(new_n747), .B2(new_n1104), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1228), .B1(new_n1108), .B2(new_n764), .C1(new_n283), .C2(new_n772), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1227), .B(new_n1229), .C1(G50), .C2(new_n760), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n776), .A2(G107), .B1(G116), .B2(new_n747), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1231), .A2(KEYINPUT122), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(KEYINPUT122), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G77), .A2(new_n763), .B1(new_n765), .B2(G303), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n513), .B2(new_n754), .C1(new_n450), .C2(new_n768), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n268), .A4(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1041), .B1(new_n820), .B2(new_n751), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT123), .Z(new_n1238));
  AOI21_X1  g1038(.A(new_n1230), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1225), .B1(new_n741), .B2(new_n1239), .C1(new_n1124), .C2(new_n734), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1154), .B2(new_n980), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1224), .A2(new_n1242), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT124), .Z(G381));
  NAND3_X1  g1044(.A1(new_n1195), .A2(new_n1161), .A3(new_n1221), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(G387), .A2(G390), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1038), .A2(new_n791), .A3(new_n1070), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(G381), .A2(new_n1248), .A3(G384), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1249), .ZN(G407));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  NAND2_X1  g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  AND2_X1   g1052(.A1(G387), .A2(G390), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1248), .B(new_n1252), .C1(new_n1253), .C2(new_n1247), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1099), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1255), .B(new_n978), .C1(new_n1010), .C2(new_n1031), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G387), .A2(G390), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1038), .A2(new_n791), .A3(new_n1070), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n791), .B1(new_n1038), .B2(new_n1070), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1256), .B(new_n1257), .C1(new_n1258), .C2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1254), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1195), .A2(G378), .A3(new_n1221), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1190), .A2(new_n1009), .A3(new_n1192), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1187), .A2(new_n935), .A3(new_n1188), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n935), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n980), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1196), .A2(new_n1220), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1161), .B1(new_n1263), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT125), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1190), .A2(new_n1192), .A3(new_n1009), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1221), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(KEYINPUT125), .A3(new_n1161), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1262), .A2(new_n1271), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n670), .A2(G213), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1158), .A2(new_n690), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1223), .A2(KEYINPUT60), .ZN(new_n1279));
  OR2_X1    g1079(.A1(new_n1223), .A2(KEYINPUT60), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(G384), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1242), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n691), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1279), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1223), .A2(KEYINPUT60), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1288), .B2(new_n1242), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1284), .A2(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .A4(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1277), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1273), .A2(KEYINPUT125), .A3(new_n1161), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT125), .B1(new_n1273), .B2(new_n1161), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1293), .B1(new_n1296), .B2(new_n1262), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1284), .B2(new_n1289), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1282), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1288), .A2(G384), .A3(new_n1242), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(KEYINPUT126), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1293), .A2(G2897), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1304), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1299), .A2(new_n1306), .A3(new_n1302), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1291), .B(new_n1292), .C1(new_n1297), .C2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1276), .B1(new_n1297), .B2(new_n1290), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1261), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1261), .A2(KEYINPUT61), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1297), .A2(KEYINPUT63), .A3(new_n1290), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1307), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1306), .B1(new_n1299), .B2(new_n1302), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1314), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1290), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1312), .B(new_n1313), .C1(new_n1319), .C2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1311), .A2(new_n1322), .ZN(G405));
  AND2_X1   g1123(.A1(new_n1254), .A2(new_n1260), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1161), .B1(new_n1195), .B2(new_n1221), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1290), .B1(new_n1246), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1325), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1327), .A2(new_n1245), .A3(new_n1320), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1324), .A2(new_n1326), .A3(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1324), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1329), .B1(new_n1330), .B2(KEYINPUT127), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT127), .ZN(new_n1332));
  AOI211_X1 g1132(.A(new_n1332), .B(new_n1324), .C1(new_n1326), .C2(new_n1328), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1331), .A2(new_n1333), .ZN(G402));
endmodule


