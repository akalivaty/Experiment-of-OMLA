//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT74), .ZN(new_n189));
  INV_X1    g003(.A(G101), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G104), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(G104), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G107), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n191), .A2(KEYINPUT75), .A3(KEYINPUT3), .A4(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  OAI22_X1  g015(.A1(new_n191), .A2(G104), .B1(KEYINPUT75), .B2(KEYINPUT3), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  AND4_X1   g017(.A1(KEYINPUT76), .A2(new_n201), .A3(new_n190), .A4(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n202), .B1(new_n199), .B2(new_n200), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT76), .B1(new_n205), .B2(new_n190), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n196), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G128), .ZN(new_n216));
  INV_X1    g030(.A(new_n211), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT64), .B1(new_n210), .B2(G143), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n212), .A3(G146), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n217), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n216), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n201), .A2(new_n190), .A3(new_n203), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT76), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n205), .A2(KEYINPUT76), .A3(new_n190), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(KEYINPUT77), .A3(new_n196), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n209), .A2(new_n225), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT79), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n195), .B1(new_n228), .B2(new_n229), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n216), .B1(new_n214), .B2(new_n223), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n209), .A2(new_n237), .A3(new_n225), .A4(new_n231), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT78), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G137), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT11), .A3(G134), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(G137), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n243), .A2(new_n245), .A3(new_n249), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT12), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n239), .A2(new_n240), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n209), .A2(new_n231), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT10), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n225), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n201), .A2(new_n203), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G101), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(KEYINPUT4), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n260), .A2(KEYINPUT4), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(new_n230), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT0), .B(G128), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n218), .A2(new_n220), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(new_n211), .ZN(new_n267));
  AND2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n211), .A2(new_n213), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n264), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n214), .A2(new_n268), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n271), .B(KEYINPUT67), .C1(new_n221), .C2(new_n265), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n263), .A2(new_n273), .B1(new_n236), .B2(new_n256), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n258), .A2(new_n274), .A3(new_n252), .ZN(new_n275));
  XNOR2_X1  g089(.A(G110), .B(G140), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n277), .A2(G227), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n236), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n282), .B1(new_n232), .B2(KEYINPUT79), .ZN(new_n283));
  AOI211_X1 g097(.A(KEYINPUT78), .B(new_n252), .C1(new_n283), .C2(new_n238), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT12), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n254), .B(new_n281), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n252), .B1(new_n258), .B2(new_n274), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n280), .B1(new_n288), .B2(new_n275), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT80), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n286), .B2(new_n290), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(KEYINPUT80), .A3(new_n292), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n239), .A2(new_n240), .A3(new_n251), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT78), .B1(new_n283), .B2(new_n238), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n300), .A2(KEYINPUT12), .B1(new_n301), .B2(new_n253), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n275), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n303), .A2(new_n279), .B1(new_n281), .B2(new_n288), .ZN(new_n304));
  OAI21_X1  g118(.A(G469), .B1(new_n304), .B2(G902), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n189), .B1(new_n299), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n270), .A2(new_n251), .A3(new_n272), .ZN(new_n309));
  INV_X1    g123(.A(G119), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G116), .ZN(new_n311));
  INV_X1    g125(.A(G116), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G119), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT2), .B(G113), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n315), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n242), .A2(G137), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n244), .A2(G134), .ZN(new_n321));
  OAI21_X1  g135(.A(G131), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n224), .A2(new_n250), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n309), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n219), .B1(new_n212), .B2(G146), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n210), .A2(KEYINPUT64), .A3(G143), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n211), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n265), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n269), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n330), .A2(new_n251), .A3(KEYINPUT65), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT65), .B1(new_n330), .B2(new_n251), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n250), .A2(new_n322), .ZN(new_n333));
  INV_X1    g147(.A(new_n223), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n333), .B1(new_n335), .B2(new_n216), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n331), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT66), .B1(new_n337), .B2(KEYINPUT30), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n330), .A2(new_n251), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT65), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n330), .A2(new_n251), .A3(KEYINPUT65), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n323), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT66), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n309), .A2(KEYINPUT30), .A3(new_n323), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT68), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n309), .A2(new_n323), .A3(KEYINPUT68), .A4(KEYINPUT30), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n338), .A2(new_n346), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n325), .B1(new_n351), .B2(new_n318), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT31), .ZN(new_n353));
  NOR2_X1   g167(.A1(G237), .A2(G953), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G210), .ZN(new_n355));
  XOR2_X1   g169(.A(new_n355), .B(KEYINPUT27), .Z(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT26), .B(G101), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n356), .B(new_n357), .Z(new_n358));
  NAND4_X1  g172(.A1(new_n352), .A2(KEYINPUT69), .A3(new_n353), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n349), .A2(new_n350), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n360), .B(new_n318), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n363), .A2(new_n353), .A3(new_n324), .A4(new_n358), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT69), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n324), .A3(new_n358), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n324), .A2(KEYINPUT28), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n324), .A2(KEYINPUT28), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n369), .A2(new_n370), .B1(new_n318), .B2(new_n343), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n358), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n368), .A2(KEYINPUT31), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n308), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT70), .B1(new_n375), .B2(KEYINPUT32), .ZN(new_n376));
  INV_X1    g190(.A(G472), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n363), .A2(new_n324), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n373), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n371), .B2(new_n358), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n369), .A2(new_n370), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n309), .A2(new_n323), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n318), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n358), .A2(KEYINPUT29), .ZN(new_n387));
  AOI21_X1  g201(.A(G902), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n377), .B1(new_n381), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n375), .B2(KEYINPUT32), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT70), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT32), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n368), .A2(KEYINPUT31), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n372), .A2(new_n373), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n366), .B2(new_n359), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n391), .B(new_n392), .C1(new_n396), .C2(new_n308), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n376), .A2(new_n390), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G217), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(G234), .B2(new_n293), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT23), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n310), .B2(G128), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n222), .A2(KEYINPUT23), .A3(G119), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n403), .B(new_n404), .C1(G119), .C2(new_n222), .ZN(new_n405));
  XNOR2_X1  g219(.A(G119), .B(G128), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT24), .B(G110), .Z(new_n407));
  OAI22_X1  g221(.A1(new_n405), .A2(G110), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G125), .B(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT16), .ZN(new_n410));
  INV_X1    g224(.A(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G125), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n412), .A2(KEYINPUT16), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(G146), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(new_n210), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n408), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(G146), .B1(new_n410), .B2(new_n413), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n414), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n405), .A2(G110), .B1(new_n406), .B2(new_n407), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT71), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(KEYINPUT71), .A3(new_n421), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n417), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT22), .B(G137), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n428), .B(KEYINPUT72), .Z(new_n430));
  OAI211_X1 g244(.A(new_n429), .B(new_n293), .C1(new_n425), .C2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT25), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n425), .ZN(new_n434));
  INV_X1    g248(.A(new_n430), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(KEYINPUT25), .A3(new_n293), .A4(new_n429), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n401), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n429), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n400), .A2(G902), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT73), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G214), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(G125), .ZN(new_n449));
  OR3_X1    g263(.A1(new_n330), .A2(KEYINPUT82), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n225), .A2(new_n449), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT82), .B1(new_n330), .B2(new_n449), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G224), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(G953), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT83), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n453), .B(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G122), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n263), .A2(new_n318), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT5), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n462), .B(G113), .C1(KEYINPUT5), .C2(new_n311), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n316), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n209), .B2(new_n231), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n459), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n464), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n234), .A2(KEYINPUT77), .ZN(new_n468));
  AOI211_X1 g282(.A(new_n208), .B(new_n195), .C1(new_n228), .C2(new_n229), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n458), .A3(new_n460), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n466), .A2(KEYINPUT6), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n473), .B(new_n459), .C1(new_n461), .C2(new_n465), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT81), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n458), .B1(new_n470), .B2(new_n460), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n473), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n457), .B(new_n472), .C1(new_n475), .C2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n458), .B(KEYINPUT8), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n234), .A2(new_n467), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n480), .B1(new_n465), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(KEYINPUT84), .B(new_n480), .C1(new_n465), .C2(new_n481), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT7), .B1(new_n454), .B2(G953), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n453), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n451), .B1(new_n449), .B2(new_n330), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n487), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n471), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G210), .B1(G237), .B2(G902), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n479), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n479), .B2(new_n492), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n448), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n187), .A2(new_n399), .A3(G953), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT92), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n212), .A2(G128), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n222), .A2(G143), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(new_n242), .ZN(new_n502));
  XNOR2_X1  g316(.A(G116), .B(G122), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n191), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n312), .A2(KEYINPUT14), .A3(G122), .ZN(new_n505));
  XOR2_X1   g319(.A(G116), .B(G122), .Z(new_n506));
  OAI211_X1 g320(.A(G107), .B(new_n505), .C1(new_n506), .C2(KEYINPUT14), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n502), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n501), .A2(new_n242), .ZN(new_n509));
  INV_X1    g323(.A(new_n504), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n503), .A2(new_n191), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(KEYINPUT89), .A2(KEYINPUT13), .ZN(new_n513));
  NOR2_X1   g327(.A1(KEYINPUT89), .A2(KEYINPUT13), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n499), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n242), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n499), .B(new_n500), .C1(new_n513), .C2(new_n514), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(KEYINPUT90), .A3(new_n518), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n512), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n508), .B1(new_n523), .B2(KEYINPUT91), .ZN(new_n524));
  INV_X1    g338(.A(new_n511), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n525), .A2(new_n504), .B1(new_n242), .B2(new_n501), .ZN(new_n526));
  INV_X1    g340(.A(new_n522), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT90), .B1(new_n517), .B2(new_n518), .ZN(new_n528));
  OAI211_X1 g342(.A(KEYINPUT91), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n498), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT91), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n498), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n529), .A4(new_n508), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n293), .ZN(new_n538));
  INV_X1    g352(.A(G478), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n538), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(G113), .B(G122), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n198), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(G143), .B1(new_n354), .B2(G214), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n354), .A2(G143), .A3(G214), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n249), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n547), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n549), .A2(new_n545), .A3(G131), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n414), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n449), .A2(G140), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT85), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n412), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT19), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n409), .A2(new_n553), .A3(KEYINPUT19), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n210), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT86), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(KEYINPUT86), .A3(new_n210), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n551), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n409), .B(new_n210), .ZN(new_n564));
  OAI211_X1 g378(.A(KEYINPUT18), .B(G131), .C1(new_n549), .C2(new_n545), .ZN(new_n565));
  NAND2_X1  g379(.A1(KEYINPUT18), .A2(G131), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n546), .A2(new_n547), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n544), .B1(new_n563), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n548), .A2(KEYINPUT17), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n419), .A3(new_n414), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n548), .A2(new_n550), .A3(KEYINPUT17), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n568), .B(new_n543), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G475), .A2(G902), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT87), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT20), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n579), .A2(new_n544), .ZN(new_n580));
  INV_X1    g394(.A(new_n574), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n293), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n577), .A2(new_n578), .B1(G475), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n410), .A2(G146), .A3(new_n413), .ZN(new_n584));
  INV_X1    g398(.A(new_n548), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n546), .A2(new_n249), .A3(new_n547), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT86), .B1(new_n558), .B2(new_n210), .ZN(new_n588));
  AOI211_X1 g402(.A(new_n560), .B(G146), .C1(new_n556), .C2(new_n557), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n543), .B1(new_n590), .B2(new_n568), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n576), .B1(new_n591), .B2(new_n581), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT87), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n575), .A2(KEYINPUT87), .A3(new_n576), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT20), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n583), .A2(KEYINPUT88), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT88), .B1(new_n583), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(G234), .A2(G237), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n600), .A2(G952), .A3(new_n277), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n600), .A2(G902), .A3(G953), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT21), .B(G898), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR4_X1   g418(.A1(new_n496), .A2(new_n541), .A3(new_n599), .A4(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n306), .A2(new_n398), .A3(new_n447), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT93), .B(G101), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G3));
  AND2_X1   g422(.A1(new_n364), .A2(new_n365), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n364), .A2(new_n365), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n374), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n377), .B1(new_n611), .B2(new_n293), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n612), .A2(new_n375), .A3(new_n446), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n306), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT88), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT20), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n582), .A2(G475), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n594), .B2(KEYINPUT20), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n615), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n538), .A2(new_n539), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n531), .A2(new_n621), .A3(new_n536), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT95), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n534), .A2(new_n623), .A3(new_n529), .A4(new_n508), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT94), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n498), .ZN(new_n626));
  INV_X1    g440(.A(new_n508), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n532), .B2(new_n533), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n498), .A2(new_n625), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n623), .A4(new_n529), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n536), .A2(KEYINPUT95), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n626), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n622), .B1(new_n632), .B2(KEYINPUT33), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n293), .A2(G478), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n620), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n583), .A2(new_n596), .A3(KEYINPUT88), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n619), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT96), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n448), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n479), .A2(new_n492), .ZN(new_n641));
  INV_X1    g455(.A(new_n493), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n479), .A2(new_n492), .A3(new_n493), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n604), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n639), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n614), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  XOR2_X1   g466(.A(new_n538), .B(new_n540), .Z(new_n653));
  NAND2_X1  g467(.A1(new_n583), .A2(new_n596), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n614), .A2(new_n648), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  OAI21_X1  g472(.A(G472), .B1(new_n396), .B2(G902), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n611), .A2(new_n307), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT97), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n425), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n435), .A2(KEYINPUT36), .ZN(new_n664));
  AOI211_X1 g478(.A(KEYINPUT97), .B(new_n417), .C1(new_n423), .C2(new_n424), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  OAI22_X1  g481(.A1(new_n662), .A2(new_n665), .B1(KEYINPUT36), .B2(new_n435), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n444), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n439), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n659), .A2(new_n660), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n659), .A2(KEYINPUT98), .A3(new_n660), .A4(new_n670), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n673), .A2(new_n306), .A3(new_n605), .A4(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  NAND2_X1  g491(.A1(new_n645), .A2(new_n670), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n601), .B1(new_n602), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n541), .A2(new_n596), .A3(new_n583), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT99), .Z(new_n684));
  NAND4_X1  g498(.A1(new_n306), .A2(new_n398), .A3(new_n679), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XOR2_X1   g500(.A(new_n681), .B(KEYINPUT39), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n306), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n619), .A2(new_n541), .A3(new_n636), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n670), .A2(new_n690), .A3(new_n640), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT101), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n643), .A2(new_n644), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n693), .B(KEYINPUT38), .Z(new_n694));
  NOR3_X1   g508(.A1(new_n689), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n378), .A2(new_n358), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n325), .A2(new_n358), .ZN(new_n697));
  AOI21_X1  g511(.A(G902), .B1(new_n697), .B2(new_n384), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n377), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n375), .B2(KEYINPUT32), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n376), .A2(new_n700), .A3(new_n397), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT100), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n695), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  NAND4_X1  g519(.A1(new_n619), .A2(new_n635), .A3(new_n636), .A4(new_n682), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n306), .A2(new_n398), .A3(new_n679), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  AND2_X1   g524(.A1(new_n398), .A2(new_n447), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT103), .B1(new_n297), .B2(new_n292), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n289), .B1(new_n302), .B2(new_n281), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n714), .B(G469), .C1(new_n715), .C2(G902), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n299), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n189), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n711), .A2(new_n649), .A3(new_n712), .A4(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n189), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n296), .A2(new_n298), .B1(new_n713), .B2(new_n716), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n398), .A2(new_n447), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n639), .A2(new_n648), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT104), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND2_X1  g542(.A1(new_n648), .A2(new_n655), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n312), .ZN(G18));
  NAND2_X1  g545(.A1(new_n619), .A2(new_n636), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n670), .A2(new_n653), .A3(new_n732), .A4(new_n646), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n398), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n299), .A2(new_n717), .A3(new_n721), .A4(new_n645), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n310), .ZN(G21));
  AOI22_X1  g552(.A1(new_n368), .A2(KEYINPUT31), .B1(new_n373), .B2(new_n385), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n308), .B1(new_n367), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n612), .A2(new_n446), .A3(new_n740), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n496), .A2(new_n604), .A3(new_n690), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n722), .A2(new_n741), .A3(new_n721), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  INV_X1    g558(.A(new_n736), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n367), .A2(new_n739), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n307), .ZN(new_n747));
  AOI21_X1  g561(.A(G902), .B1(new_n367), .B2(new_n374), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n747), .B(new_n670), .C1(new_n748), .C2(new_n377), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n599), .A2(new_n707), .A3(new_n635), .A4(new_n682), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n706), .A2(KEYINPUT102), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n745), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  NOR2_X1   g569(.A1(new_n660), .A2(new_n392), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n375), .A2(KEYINPUT32), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT107), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n389), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n660), .A2(new_n392), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n375), .A2(KEYINPUT32), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n758), .A2(new_n759), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n447), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n764), .A2(KEYINPUT108), .A3(new_n447), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n643), .A2(new_n721), .A3(new_n448), .A4(new_n644), .ZN(new_n770));
  NAND2_X1  g584(.A1(G469), .A2(G902), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT105), .Z(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n304), .B2(G469), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n770), .B1(new_n299), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(KEYINPUT42), .A3(new_n708), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n774), .A2(new_n398), .A3(new_n447), .A4(new_n708), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT106), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n777), .A2(KEYINPUT106), .A3(new_n778), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n769), .A2(new_n776), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n249), .ZN(G33));
  NAND4_X1  g598(.A1(new_n774), .A2(new_n398), .A3(new_n447), .A4(new_n684), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT109), .B(G134), .Z(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(G36));
  AND2_X1   g601(.A1(new_n304), .A2(KEYINPUT45), .ZN(new_n788));
  OAI21_X1  g602(.A(G469), .B1(new_n304), .B2(KEYINPUT45), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n772), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT46), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n299), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(KEYINPUT110), .A3(new_n299), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n791), .B2(KEYINPUT46), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n791), .A2(new_n797), .A3(KEYINPUT46), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n795), .A2(new_n796), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n721), .A3(new_n687), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n732), .A2(new_n635), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT43), .Z(new_n803));
  NAND2_X1  g617(.A1(new_n659), .A2(new_n660), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n803), .A2(new_n804), .A3(new_n670), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT44), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n693), .A2(new_n640), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n805), .B2(KEYINPUT44), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n801), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(new_n244), .ZN(G39));
  NAND2_X1  g626(.A1(new_n800), .A2(new_n721), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n800), .A2(KEYINPUT47), .A3(new_n721), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n809), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n398), .A2(new_n818), .A3(new_n752), .A4(new_n447), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  NAND3_X1  g635(.A1(new_n447), .A2(new_n721), .A3(new_n448), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n802), .B(new_n822), .C1(new_n718), .C2(KEYINPUT49), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT113), .ZN(new_n824));
  INV_X1    g638(.A(new_n702), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n718), .A2(KEYINPUT49), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n824), .A2(new_n694), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n398), .A2(new_n679), .ZN(new_n829));
  INV_X1    g643(.A(new_n298), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT80), .B1(new_n297), .B2(new_n292), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n305), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n684), .A3(new_n721), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n612), .A2(new_n740), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n708), .A2(new_n670), .A3(new_n834), .ZN(new_n835));
  OAI22_X1  g649(.A1(new_n829), .A2(new_n833), .B1(new_n835), .B2(new_n736), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n299), .A2(new_n773), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n439), .A2(KEYINPUT116), .A3(new_n669), .A4(new_n682), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n721), .ZN(new_n841));
  INV_X1    g655(.A(new_n669), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n438), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT116), .B1(new_n843), .B2(new_n682), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n496), .A2(new_n690), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n701), .A2(new_n839), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n709), .A2(KEYINPUT52), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n754), .A2(new_n685), .A3(KEYINPUT115), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n838), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n754), .A2(new_n685), .A3(new_n709), .A4(new_n847), .ZN(new_n851));
  XNOR2_X1  g665(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n850), .A2(KEYINPUT118), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT118), .B1(new_n850), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n743), .B1(new_n735), .B2(new_n736), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n730), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n653), .B1(new_n619), .B2(new_n636), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT114), .B1(new_n637), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n859), .A2(KEYINPUT114), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n647), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n306), .A3(new_n613), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n675), .A2(new_n606), .A3(new_n863), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n843), .A2(new_n541), .A3(new_n654), .A4(new_n681), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n306), .A2(new_n398), .A3(new_n809), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n753), .A2(new_n774), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n785), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n726), .A2(new_n858), .A3(new_n864), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n769), .A2(new_n776), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n781), .A2(new_n782), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n828), .B1(new_n856), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n709), .A2(new_n847), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n685), .A4(new_n754), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n870), .A2(new_n880), .A3(new_n873), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n875), .B1(new_n828), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT54), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n870), .A2(new_n873), .A3(KEYINPUT53), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n884), .B1(new_n856), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n850), .A2(new_n853), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n850), .A2(KEYINPUT118), .A3(new_n853), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n783), .A2(new_n869), .A3(new_n828), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(KEYINPUT120), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n878), .A2(new_n879), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n783), .A2(new_n896), .A3(new_n869), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n895), .B1(new_n897), .B2(KEYINPUT53), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n881), .A2(KEYINPUT119), .A3(new_n828), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n894), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n883), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n803), .A2(new_n601), .A3(new_n741), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n904), .A2(new_n640), .A3(new_n694), .A4(new_n719), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT50), .Z(new_n906));
  INV_X1    g720(.A(new_n601), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n718), .A2(new_n907), .A3(new_n770), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n908), .A2(new_n447), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n599), .A2(new_n635), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n825), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n908), .A2(new_n803), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n670), .A3(new_n834), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n906), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n815), .B(new_n816), .C1(new_n721), .C2(new_n718), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n904), .A2(new_n809), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT121), .Z(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n918), .A2(KEYINPUT51), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n769), .A2(new_n912), .ZN(new_n920));
  XOR2_X1   g734(.A(KEYINPUT122), .B(KEYINPUT48), .Z(new_n921));
  OR2_X1    g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n825), .A2(new_n639), .A3(new_n909), .ZN(new_n924));
  INV_X1    g738(.A(G952), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n925), .B(G953), .C1(new_n904), .C2(new_n745), .ZN(new_n926));
  AND4_X1   g740(.A1(new_n922), .A2(new_n923), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n918), .B2(KEYINPUT51), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n903), .A2(new_n919), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(G952), .A2(G953), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n827), .B1(new_n929), .B2(new_n930), .ZN(G75));
  NAND2_X1  g745(.A1(new_n894), .A2(new_n900), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(G210), .A3(G902), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n472), .B1(new_n475), .B2(new_n478), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n457), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n933), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n933), .B2(new_n934), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n277), .A2(G952), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G51));
  XNOR2_X1  g755(.A(new_n772), .B(KEYINPUT57), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n894), .A2(new_n901), .A3(new_n900), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n901), .B1(new_n894), .B2(new_n900), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n291), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n293), .B1(new_n894), .B2(new_n900), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n790), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n940), .B1(new_n946), .B2(new_n948), .ZN(G54));
  NAND3_X1  g763(.A1(new_n947), .A2(KEYINPUT58), .A3(G475), .ZN(new_n950));
  INV_X1    g764(.A(new_n575), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n940), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n947), .A2(KEYINPUT58), .A3(G475), .A4(new_n575), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G60));
  INV_X1    g769(.A(new_n633), .ZN(new_n956));
  NAND2_X1  g770(.A1(G478), .A2(G902), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT59), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n903), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n958), .ZN(new_n960));
  INV_X1    g774(.A(new_n944), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(new_n902), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n959), .A2(new_n962), .A3(new_n940), .ZN(G63));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT60), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n667), .A2(new_n668), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT123), .Z(new_n969));
  NAND3_X1  g783(.A1(new_n932), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n953), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n966), .B1(new_n894), .B2(new_n900), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(new_n441), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n964), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT124), .B1(new_n972), .B2(new_n441), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n940), .B1(new_n972), .B2(new_n969), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT124), .ZN(new_n977));
  AOI22_X1  g791(.A1(new_n886), .A2(new_n893), .B1(new_n898), .B2(new_n899), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n977), .B(new_n440), .C1(new_n978), .C2(new_n966), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT61), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n974), .A2(new_n980), .ZN(G66));
  INV_X1    g795(.A(new_n603), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n277), .B1(new_n982), .B2(G224), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n726), .A2(new_n858), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n864), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n983), .B1(new_n985), .B2(new_n277), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n935), .B1(G898), .B2(new_n277), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n986), .B(new_n987), .Z(G69));
  NAND2_X1  g802(.A1(G227), .A2(G900), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n680), .A2(G953), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n990), .A2(KEYINPUT127), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(KEYINPUT127), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n811), .B1(new_n817), .B2(new_n819), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n769), .A2(new_n846), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n801), .A2(new_n995), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n838), .A2(new_n849), .ZN(new_n997));
  AND4_X1   g811(.A1(new_n709), .A2(new_n873), .A3(new_n785), .A4(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n994), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n993), .B1(new_n999), .B2(new_n277), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n558), .B(KEYINPUT125), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n351), .B(new_n1002), .ZN(new_n1003));
  OAI211_X1 g817(.A(G953), .B(new_n989), .C1(new_n1001), .C2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n704), .A2(new_n997), .A3(new_n709), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT62), .Z(new_n1006));
  AOI21_X1  g820(.A(new_n818), .B1(new_n861), .B2(new_n860), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n711), .A2(new_n306), .A3(new_n687), .A4(new_n1007), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT126), .Z(new_n1009));
  AND3_X1   g823(.A1(new_n994), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1003), .B1(new_n1010), .B2(G953), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n989), .A2(G953), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n1011), .B(new_n1012), .C1(new_n1000), .C2(new_n1003), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1004), .A2(new_n1013), .ZN(G72));
  INV_X1    g828(.A(new_n985), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n994), .A2(new_n1006), .A3(new_n1015), .A4(new_n1009), .ZN(new_n1016));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  AOI21_X1  g832(.A(new_n696), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n363), .A2(new_n697), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n994), .A2(new_n1015), .A3(new_n996), .A4(new_n998), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1020), .B1(new_n1021), .B2(new_n1018), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n379), .A2(new_n368), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n882), .A2(new_n1018), .A3(new_n1023), .ZN(new_n1024));
  NOR4_X1   g838(.A1(new_n1019), .A2(new_n1022), .A3(new_n1024), .A4(new_n940), .ZN(G57));
endmodule


