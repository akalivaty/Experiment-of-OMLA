

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581;

  XNOR2_X1 U324 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n420) );
  XNOR2_X1 U325 ( .A(n395), .B(n394), .ZN(n396) );
  NOR2_X1 U326 ( .A1(n483), .A2(n575), .ZN(n484) );
  XNOR2_X1 U327 ( .A(n441), .B(n440), .ZN(n519) );
  XNOR2_X1 U328 ( .A(n339), .B(n403), .ZN(n517) );
  XOR2_X1 U329 ( .A(KEYINPUT74), .B(n340), .Z(n292) );
  AND2_X1 U330 ( .A1(G226GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U331 ( .A(KEYINPUT21), .B(KEYINPUT86), .Z(n294) );
  INV_X1 U332 ( .A(KEYINPUT78), .ZN(n394) );
  INV_X1 U333 ( .A(KEYINPUT32), .ZN(n345) );
  XNOR2_X1 U334 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U335 ( .A(n397), .B(n396), .ZN(n401) );
  XNOR2_X1 U336 ( .A(n377), .B(n293), .ZN(n335) );
  XNOR2_X1 U337 ( .A(n348), .B(n347), .ZN(n351) );
  NOR2_X1 U338 ( .A1(n522), .A2(n544), .ZN(n526) );
  XNOR2_X1 U339 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U340 ( .A(n407), .B(n406), .Z(n575) );
  XNOR2_X1 U341 ( .A(KEYINPUT38), .B(n487), .ZN(n497) );
  XNOR2_X1 U342 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U343 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(G197GAT), .B(G218GAT), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n294), .B(n295), .ZN(n332) );
  XOR2_X1 U346 ( .A(G155GAT), .B(n332), .Z(n301) );
  XNOR2_X1 U347 ( .A(G148GAT), .B(KEYINPUT72), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n296), .B(KEYINPUT71), .ZN(n297) );
  XOR2_X1 U349 ( .A(n297), .B(G204GAT), .Z(n299) );
  XNOR2_X1 U350 ( .A(G78GAT), .B(G106GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n353) );
  XNOR2_X1 U352 ( .A(G22GAT), .B(n353), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n307) );
  XOR2_X1 U354 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n303) );
  XNOR2_X1 U355 ( .A(G141GAT), .B(G162GAT), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n314) );
  XOR2_X1 U357 ( .A(KEYINPUT23), .B(n314), .Z(n305) );
  NAND2_X1 U358 ( .A1(G228GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U360 ( .A(n307), .B(n306), .Z(n312) );
  XOR2_X1 U361 ( .A(G211GAT), .B(KEYINPUT22), .Z(n309) );
  XNOR2_X1 U362 ( .A(KEYINPUT85), .B(KEYINPUT24), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U364 ( .A(G50GAT), .B(n310), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n462) );
  XNOR2_X1 U366 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n313), .B(G120GAT), .ZN(n433) );
  XNOR2_X1 U368 ( .A(n433), .B(n314), .ZN(n328) );
  XNOR2_X1 U369 ( .A(G1GAT), .B(G127GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n315), .B(G155GAT), .ZN(n397) );
  XOR2_X1 U371 ( .A(G29GAT), .B(G134GAT), .Z(n376) );
  XOR2_X1 U372 ( .A(n397), .B(n376), .Z(n317) );
  XNOR2_X1 U373 ( .A(G148GAT), .B(G85GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U375 ( .A(KEYINPUT5), .B(G57GAT), .Z(n319) );
  NAND2_X1 U376 ( .A1(G225GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U378 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U379 ( .A(KEYINPUT6), .B(KEYINPUT88), .Z(n323) );
  XNOR2_X1 U380 ( .A(KEYINPUT87), .B(KEYINPUT4), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n324), .B(KEYINPUT1), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n468) );
  XNOR2_X1 U385 ( .A(KEYINPUT89), .B(n468), .ZN(n515) );
  XOR2_X1 U386 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n330) );
  XNOR2_X1 U387 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n431) );
  XNOR2_X1 U389 ( .A(G176GAT), .B(G92GAT), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n331), .B(G64GAT), .ZN(n340) );
  XOR2_X1 U391 ( .A(KEYINPUT90), .B(n340), .Z(n334) );
  XNOR2_X1 U392 ( .A(G204GAT), .B(n332), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n336) );
  XOR2_X1 U394 ( .A(G36GAT), .B(G190GAT), .Z(n377) );
  XNOR2_X1 U395 ( .A(n431), .B(n337), .ZN(n339) );
  XNOR2_X1 U396 ( .A(G8GAT), .B(G183GAT), .ZN(n338) );
  XOR2_X1 U397 ( .A(n338), .B(G211GAT), .Z(n403) );
  XNOR2_X1 U398 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n292), .B(n341), .ZN(n348) );
  XOR2_X1 U400 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n343) );
  NAND2_X1 U401 ( .A1(G230GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U403 ( .A(KEYINPUT31), .B(n344), .ZN(n346) );
  XOR2_X1 U404 ( .A(KEYINPUT13), .B(KEYINPUT68), .Z(n350) );
  XNOR2_X1 U405 ( .A(G71GAT), .B(G57GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n402) );
  XNOR2_X1 U407 ( .A(n351), .B(n402), .ZN(n355) );
  XNOR2_X1 U408 ( .A(G99GAT), .B(G85GAT), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n352), .B(KEYINPUT73), .ZN(n375) );
  XOR2_X1 U410 ( .A(n353), .B(n375), .Z(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n571) );
  XOR2_X1 U412 ( .A(n571), .B(KEYINPUT41), .Z(n501) );
  INV_X1 U413 ( .A(n501), .ZN(n530) );
  XOR2_X1 U414 ( .A(G22GAT), .B(G15GAT), .Z(n392) );
  XOR2_X1 U415 ( .A(G141GAT), .B(G197GAT), .Z(n357) );
  XNOR2_X1 U416 ( .A(G29GAT), .B(G36GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U418 ( .A(n392), .B(n358), .Z(n360) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U421 ( .A(n361), .B(KEYINPUT66), .Z(n365) );
  XOR2_X1 U422 ( .A(G43GAT), .B(G50GAT), .Z(n363) );
  XNOR2_X1 U423 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n379) );
  XNOR2_X1 U425 ( .A(n379), .B(KEYINPUT30), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n373) );
  XOR2_X1 U427 ( .A(G8GAT), .B(G1GAT), .Z(n367) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(G113GAT), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U430 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n369) );
  XNOR2_X1 U431 ( .A(KEYINPUT65), .B(KEYINPUT64), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U433 ( .A(n371), .B(n370), .Z(n372) );
  XOR2_X1 U434 ( .A(n373), .B(n372), .Z(n546) );
  NAND2_X1 U435 ( .A1(n530), .A2(n546), .ZN(n374) );
  XNOR2_X1 U436 ( .A(KEYINPUT46), .B(n374), .ZN(n409) );
  XNOR2_X1 U437 ( .A(n376), .B(n375), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n383) );
  XOR2_X1 U439 ( .A(n379), .B(G92GAT), .Z(n381) );
  NAND2_X1 U440 ( .A1(G232GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U442 ( .A(n383), .B(n382), .Z(n391) );
  XOR2_X1 U443 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n385) );
  XNOR2_X1 U444 ( .A(G218GAT), .B(KEYINPUT75), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U446 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n387) );
  XNOR2_X1 U447 ( .A(G106GAT), .B(G162GAT), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U450 ( .A(n391), .B(n390), .Z(n556) );
  XNOR2_X1 U451 ( .A(n392), .B(G78GAT), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n393), .B(G64GAT), .ZN(n407) );
  NAND2_X1 U453 ( .A1(G231GAT), .A2(G233GAT), .ZN(n395) );
  XOR2_X1 U454 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n399) );
  XNOR2_X1 U455 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U457 ( .A(n401), .B(n400), .Z(n405) );
  XOR2_X1 U458 ( .A(n403), .B(n402), .Z(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U460 ( .A(KEYINPUT107), .B(n575), .Z(n560) );
  NOR2_X1 U461 ( .A1(n556), .A2(n560), .ZN(n408) );
  AND2_X1 U462 ( .A1(n409), .A2(n408), .ZN(n411) );
  XNOR2_X1 U463 ( .A(KEYINPUT47), .B(KEYINPUT108), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n411), .B(n410), .ZN(n417) );
  XOR2_X1 U465 ( .A(KEYINPUT45), .B(KEYINPUT109), .Z(n413) );
  XNOR2_X1 U466 ( .A(KEYINPUT36), .B(n556), .ZN(n578) );
  NAND2_X1 U467 ( .A1(n575), .A2(n578), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n414) );
  NOR2_X1 U469 ( .A1(n546), .A2(n414), .ZN(n415) );
  NAND2_X1 U470 ( .A1(n571), .A2(n415), .ZN(n416) );
  NAND2_X1 U471 ( .A1(n417), .A2(n416), .ZN(n419) );
  XOR2_X1 U472 ( .A(KEYINPUT110), .B(KEYINPUT48), .Z(n418) );
  XOR2_X1 U473 ( .A(n419), .B(n418), .Z(n542) );
  NAND2_X1 U474 ( .A1(n517), .A2(n542), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n422) );
  NOR2_X1 U476 ( .A1(n515), .A2(n422), .ZN(n564) );
  NAND2_X1 U477 ( .A1(n462), .A2(n564), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n423), .B(KEYINPUT55), .ZN(n442) );
  XOR2_X1 U479 ( .A(KEYINPUT20), .B(G183GAT), .Z(n425) );
  XNOR2_X1 U480 ( .A(KEYINPUT82), .B(KEYINPUT84), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n441) );
  XOR2_X1 U482 ( .A(KEYINPUT83), .B(G127GAT), .Z(n427) );
  XNOR2_X1 U483 ( .A(G134GAT), .B(G190GAT), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U485 ( .A(G43GAT), .B(G99GAT), .Z(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n437) );
  XNOR2_X1 U487 ( .A(KEYINPUT81), .B(G71GAT), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n430), .B(G176GAT), .ZN(n432) );
  XOR2_X1 U489 ( .A(n432), .B(n431), .Z(n435) );
  XNOR2_X1 U490 ( .A(G15GAT), .B(n433), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n439) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  AND2_X1 U495 ( .A1(n442), .A2(n519), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n443), .B(KEYINPUT121), .ZN(n559) );
  INV_X1 U497 ( .A(n546), .ZN(n565) );
  NOR2_X1 U498 ( .A1(n559), .A2(n565), .ZN(n446) );
  XNOR2_X1 U499 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n444), .B(KEYINPUT123), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(G1348GAT) );
  NOR2_X1 U502 ( .A1(n559), .A2(n501), .ZN(n449) );
  XNOR2_X1 U503 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n447), .B(G176GAT), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n449), .B(n448), .ZN(G1349GAT) );
  INV_X1 U506 ( .A(n556), .ZN(n454) );
  NOR2_X1 U507 ( .A1(n559), .A2(n454), .ZN(n453) );
  XNOR2_X1 U508 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n451) );
  INV_X1 U509 ( .A(G190GAT), .ZN(n450) );
  XOR2_X1 U510 ( .A(KEYINPUT34), .B(KEYINPUT94), .Z(n474) );
  NAND2_X1 U511 ( .A1(n546), .A2(n571), .ZN(n485) );
  NAND2_X1 U512 ( .A1(n454), .A2(n575), .ZN(n457) );
  XNOR2_X1 U513 ( .A(KEYINPUT16), .B(KEYINPUT80), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n455), .B(KEYINPUT79), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(n472) );
  INV_X1 U516 ( .A(n519), .ZN(n528) );
  XOR2_X1 U517 ( .A(n462), .B(KEYINPUT28), .Z(n522) );
  XNOR2_X1 U518 ( .A(KEYINPUT27), .B(n517), .ZN(n464) );
  NAND2_X1 U519 ( .A1(n464), .A2(n515), .ZN(n544) );
  NAND2_X1 U520 ( .A1(n528), .A2(n526), .ZN(n458) );
  XOR2_X1 U521 ( .A(KEYINPUT91), .B(n458), .Z(n471) );
  NAND2_X1 U522 ( .A1(n519), .A2(n517), .ZN(n459) );
  NAND2_X1 U523 ( .A1(n459), .A2(n462), .ZN(n460) );
  XNOR2_X1 U524 ( .A(n460), .B(KEYINPUT93), .ZN(n461) );
  XNOR2_X1 U525 ( .A(KEYINPUT25), .B(n461), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n519), .A2(n462), .ZN(n463) );
  XNOR2_X1 U527 ( .A(n463), .B(KEYINPUT26), .ZN(n563) );
  NAND2_X1 U528 ( .A1(n464), .A2(n563), .ZN(n465) );
  XNOR2_X1 U529 ( .A(KEYINPUT92), .B(n465), .ZN(n466) );
  NAND2_X1 U530 ( .A1(n467), .A2(n466), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U532 ( .A1(n471), .A2(n470), .ZN(n482) );
  NAND2_X1 U533 ( .A1(n472), .A2(n482), .ZN(n503) );
  NOR2_X1 U534 ( .A1(n485), .A2(n503), .ZN(n479) );
  NAND2_X1 U535 ( .A1(n479), .A2(n515), .ZN(n473) );
  XNOR2_X1 U536 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U537 ( .A(G1GAT), .B(n475), .Z(G1324GAT) );
  NAND2_X1 U538 ( .A1(n517), .A2(n479), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U541 ( .A1(n479), .A2(n519), .ZN(n477) );
  XNOR2_X1 U542 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  XOR2_X1 U543 ( .A(G22GAT), .B(KEYINPUT95), .Z(n481) );
  NAND2_X1 U544 ( .A1(n479), .A2(n522), .ZN(n480) );
  XNOR2_X1 U545 ( .A(n481), .B(n480), .ZN(G1327GAT) );
  NAND2_X1 U546 ( .A1(n578), .A2(n482), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(KEYINPUT37), .ZN(n514) );
  NOR2_X1 U548 ( .A1(n514), .A2(n485), .ZN(n486) );
  XOR2_X1 U549 ( .A(KEYINPUT97), .B(n486), .Z(n487) );
  NAND2_X1 U550 ( .A1(n497), .A2(n515), .ZN(n491) );
  XOR2_X1 U551 ( .A(KEYINPUT96), .B(KEYINPUT39), .Z(n489) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT98), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  XOR2_X1 U555 ( .A(G36GAT), .B(KEYINPUT99), .Z(n493) );
  NAND2_X1 U556 ( .A1(n497), .A2(n517), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(G1329GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT100), .Z(n495) );
  NAND2_X1 U559 ( .A1(n497), .A2(n519), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U561 ( .A(G43GAT), .B(n496), .Z(G1330GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n499) );
  NAND2_X1 U563 ( .A1(n522), .A2(n497), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  NOR2_X1 U566 ( .A1(n501), .A2(n546), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n502), .B(KEYINPUT103), .ZN(n513) );
  NOR2_X1 U568 ( .A1(n503), .A2(n513), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n504), .B(KEYINPUT104), .ZN(n510) );
  NAND2_X1 U570 ( .A1(n510), .A2(n515), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n505), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n517), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT105), .Z(n509) );
  NAND2_X1 U576 ( .A1(n510), .A2(n519), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U579 ( .A1(n522), .A2(n510), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n523), .A2(n515), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n517), .A2(n523), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n523), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n520), .B(KEYINPUT106), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  NAND2_X1 U592 ( .A1(n526), .A2(n542), .ZN(n527) );
  NOR2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n539), .A2(n546), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n529), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U597 ( .A1(n539), .A2(n530), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT111), .B(KEYINPUT50), .Z(n534) );
  NAND2_X1 U600 ( .A1(n539), .A2(n560), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n537) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U606 ( .A(KEYINPUT112), .B(n538), .Z(n541) );
  NAND2_X1 U607 ( .A1(n539), .A2(n556), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n542), .A2(n563), .ZN(n543) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(KEYINPUT115), .B(n545), .Z(n557) );
  NAND2_X1 U612 ( .A1(n557), .A2(n546), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(KEYINPUT116), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n550) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(KEYINPUT117), .B(n551), .Z(n553) );
  NAND2_X1 U619 ( .A1(n557), .A2(n530), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  XOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT119), .Z(n555) );
  NAND2_X1 U622 ( .A1(n557), .A2(n575), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n558), .ZN(G1347GAT) );
  INV_X1 U626 ( .A(n559), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n574) );
  NOR2_X1 U630 ( .A1(n565), .A2(n574), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT59), .B(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n574), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  INV_X1 U639 ( .A(n574), .ZN(n579) );
  AND2_X1 U640 ( .A1(n575), .A2(n579), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(KEYINPUT62), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

