//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  OR2_X1    g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT68), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  AOI22_X1  g032(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n465), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n468), .A2(G136), .ZN(new_n473));
  INV_X1    g048(.A(G124), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n466), .A2(new_n467), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n480));
  OAI221_X1 g055(.A(G2104), .B1(G112), .B2(new_n469), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n477), .A2(new_n482), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n469), .B2(G114), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n486), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n485), .A2(new_n487), .A3(new_n488), .A4(G2104), .ZN(new_n489));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n469), .C1(new_n460), .C2(new_n461), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n475), .A2(new_n494), .A3(G138), .A4(new_n469), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G50), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n497), .B2(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(new_n505), .B1(new_n498), .B2(new_n499), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n503), .A2(new_n505), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n509), .A2(new_n513), .ZN(G166));
  XOR2_X1   g089(.A(KEYINPUT73), .B(G89), .Z(new_n515));
  NAND2_X1  g090(.A1(new_n506), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n516), .A2(KEYINPUT74), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n500), .A2(G51), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(KEYINPUT5), .B1(new_n504), .B2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n524), .B1(new_n503), .B2(new_n505), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n519), .B(new_n520), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(KEYINPUT74), .B1(new_n516), .B2(new_n518), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n506), .A2(G90), .B1(new_n500), .B2(G52), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n528), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n534), .B1(new_n537), .B2(G651), .ZN(G171));
  NAND3_X1  g113(.A1(new_n525), .A2(G56), .A3(new_n527), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n512), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT75), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n506), .A2(G81), .B1(new_n500), .B2(G43), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n544), .B1(new_n541), .B2(KEYINPUT75), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n548), .B(KEYINPUT76), .Z(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(G65), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n503), .B2(new_n505), .ZN(new_n554));
  AND2_X1   g129(.A1(G78), .A2(G543), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT77), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n558), .B(G651), .C1(new_n554), .C2(new_n555), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n500), .A2(G53), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n500), .A2(new_n563), .A3(G53), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n562), .A2(new_n564), .B1(G91), .B2(new_n506), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n560), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  OR2_X1    g142(.A1(new_n530), .A2(new_n531), .ZN(G286));
  OR2_X1    g143(.A1(new_n509), .A2(new_n513), .ZN(G303));
  NOR2_X1   g144(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n526), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n571), .B2(G74), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n506), .A2(G87), .B1(new_n500), .B2(G49), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G288));
  AOI22_X1  g149(.A1(new_n506), .A2(G86), .B1(new_n500), .B2(G48), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n503), .B2(new_n505), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n576), .B(G651), .C1(new_n578), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G61), .B1(new_n521), .B2(new_n522), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(new_n579), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n576), .B1(new_n584), .B2(G651), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n571), .A2(G60), .ZN(new_n588));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n512), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n500), .A2(G47), .ZN(new_n591));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n507), .B2(new_n592), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n590), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(new_n506), .A2(G92), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT10), .Z(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n523), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n500), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G171), .ZN(G284));
  OAI21_X1  g179(.A(new_n603), .B1(new_n602), .B2(G171), .ZN(G321));
  NAND2_X1  g180(.A1(G299), .A2(new_n602), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G168), .B2(new_n602), .ZN(G297));
  XOR2_X1   g182(.A(G297), .B(KEYINPUT79), .Z(G280));
  INV_X1    g183(.A(new_n601), .ZN(new_n609));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n475), .A2(new_n470), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n468), .A2(G135), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n469), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(G123), .ZN(new_n625));
  OAI221_X1 g200(.A(new_n622), .B1(new_n623), .B2(new_n624), .C1(new_n625), .C2(new_n476), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND3_X1  g202(.A1(new_n620), .A2(new_n621), .A3(new_n627), .ZN(G156));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n634), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(new_n642), .A3(G14), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(G401));
  XNOR2_X1  g219(.A(G2084), .B(G2090), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(KEYINPUT17), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n648), .B1(new_n649), .B2(new_n646), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT80), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n646), .A2(new_n647), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n652), .A2(new_n645), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT18), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n646), .A2(new_n645), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n651), .B(new_n654), .C1(new_n649), .C2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2096), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1981), .B(G1986), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  INV_X1    g246(.A(new_n664), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n666), .A2(new_n667), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n675), .A3(new_n673), .ZN(new_n676));
  NAND4_X1  g251(.A1(new_n670), .A2(new_n671), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n681), .B1(new_n679), .B2(new_n682), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n661), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n677), .B(new_n678), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(new_n680), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n688), .A2(new_n660), .A3(new_n683), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  XOR2_X1   g266(.A(KEYINPUT86), .B(KEYINPUT25), .Z(new_n692));
  NAND3_X1  g267(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n468), .A2(G139), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n694), .B(new_n695), .C1(new_n469), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT87), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n699), .B2(G33), .ZN(new_n701));
  INV_X1    g276(.A(G2072), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n609), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G4), .B2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G1348), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n701), .A2(new_n702), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n703), .A2(G20), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT23), .Z(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G299), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1956), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n707), .B(new_n711), .C1(new_n702), .C2(new_n701), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n699), .A2(G32), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT90), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT26), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n470), .A2(G105), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT89), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n462), .A2(new_n469), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G129), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n468), .A2(G141), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n713), .B1(new_n723), .B2(new_n699), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT91), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G34), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n728), .A2(KEYINPUT24), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(KEYINPUT24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n699), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G160), .B2(new_n699), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT88), .B(G2084), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G27), .A2(G29), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G164), .B2(G29), .ZN(new_n736));
  INV_X1    g311(.A(G2078), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n727), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT31), .B(G11), .Z(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT30), .B(G28), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n699), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n699), .A2(G35), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT95), .ZN(new_n744));
  INV_X1    g319(.A(G162), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n747));
  INV_X1    g322(.A(G2090), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n742), .B1(new_n699), .B2(new_n626), .C1(new_n746), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n749), .B2(new_n746), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n706), .B2(new_n705), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n724), .A2(new_n726), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT92), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n699), .A2(G26), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT28), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n719), .A2(G128), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n468), .A2(G140), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT85), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n757), .A2(KEYINPUT85), .A3(new_n758), .A4(new_n760), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n756), .B1(new_n765), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2067), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n754), .A2(new_n767), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n712), .A2(new_n739), .A3(new_n752), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(G168), .A2(G16), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(KEYINPUT93), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(KEYINPUT93), .B2(new_n770), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1966), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n703), .A2(G5), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G171), .B2(new_n703), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT94), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1961), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n703), .A2(G19), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n546), .B2(new_n703), .ZN(new_n780));
  INV_X1    g355(.A(G1341), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n769), .A2(new_n774), .A3(new_n778), .A4(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G288), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(new_n703), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n703), .B2(G23), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT33), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G1976), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G22), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G166), .B2(G16), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT83), .B(G1971), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT84), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G6), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n586), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT32), .B(G1981), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n787), .B2(G1976), .ZN(new_n799));
  OR3_X1    g374(.A1(new_n794), .A2(new_n799), .A3(KEYINPUT34), .ZN(new_n800));
  OAI21_X1  g375(.A(KEYINPUT34), .B1(new_n794), .B2(new_n799), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n590), .A2(new_n593), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n802), .A2(new_n703), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n703), .B2(G24), .ZN(new_n804));
  INV_X1    g379(.A(G1986), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n699), .A2(G25), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n719), .A2(G119), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n468), .A2(G131), .ZN(new_n810));
  OR2_X1    g385(.A1(G95), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n808), .B1(new_n814), .B2(new_n699), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  XOR2_X1   g391(.A(new_n815), .B(new_n816), .Z(new_n817));
  NOR3_X1   g392(.A1(new_n806), .A2(new_n807), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n800), .A2(new_n801), .A3(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT36), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(KEYINPUT36), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n783), .B1(new_n820), .B2(new_n821), .ZN(G311));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  INV_X1    g398(.A(new_n783), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(G150));
  NAND2_X1  g400(.A1(new_n609), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  INV_X1    g403(.A(G67), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n528), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G651), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n506), .A2(G93), .B1(new_n500), .B2(G55), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n543), .B2(new_n545), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT75), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n539), .A2(new_n540), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n836), .B2(new_n512), .ZN(new_n837));
  INV_X1    g412(.A(new_n832), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n830), .B2(G651), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n837), .A2(new_n839), .A3(new_n542), .A4(new_n544), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n827), .B(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n844));
  INV_X1    g419(.A(G860), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n839), .A2(new_n845), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(G145));
  XNOR2_X1  g425(.A(G160), .B(new_n626), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G162), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n765), .A2(G164), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n723), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n765), .A2(G164), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n763), .A2(new_n764), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n493), .A2(new_n495), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n489), .A2(new_n490), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n723), .B1(new_n862), .B2(new_n853), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n698), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n855), .B1(new_n854), .B2(new_n856), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n723), .A3(new_n853), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n697), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G130), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n469), .A2(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n476), .A2(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(G142), .B2(new_n468), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n617), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n813), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n864), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n874), .B1(new_n864), .B2(new_n867), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n852), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT97), .B(G37), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n852), .B(KEYINPUT99), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n875), .B(new_n880), .C1(new_n877), .C2(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n877), .A2(new_n881), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n878), .B(new_n879), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g460(.A1(new_n839), .A2(G868), .ZN(new_n886));
  NAND2_X1  g461(.A1(G290), .A2(new_n586), .ZN(new_n887));
  XNOR2_X1  g462(.A(G288), .B(G303), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n802), .A2(G305), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n888), .B1(new_n887), .B2(new_n889), .ZN(new_n892));
  OR3_X1    g467(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT42), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n892), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(KEYINPUT101), .A3(new_n890), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n891), .B2(new_n892), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n894), .B1(new_n899), .B2(KEYINPUT42), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n841), .B(new_n612), .Z(new_n901));
  INV_X1    g476(.A(G299), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n601), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT100), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n609), .A2(G299), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n601), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n609), .B2(G299), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n908), .A2(new_n909), .B1(new_n903), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n901), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n905), .A2(new_n903), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n901), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n900), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n602), .B1(new_n900), .B2(new_n914), .ZN(new_n916));
  AOI211_X1 g491(.A(KEYINPUT102), .B(new_n886), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(KEYINPUT102), .B2(new_n918), .ZN(G295));
  AOI21_X1  g494(.A(new_n917), .B1(KEYINPUT102), .B2(new_n918), .ZN(G331));
  AND2_X1   g495(.A1(new_n896), .A2(new_n898), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  NAND2_X1  g497(.A1(G286), .A2(G301), .ZN(new_n923));
  NAND2_X1  g498(.A1(G168), .A2(G171), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n841), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n834), .A2(new_n923), .A3(new_n840), .A4(new_n924), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n913), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n926), .A2(KEYINPUT104), .A3(new_n913), .A4(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n841), .A2(new_n925), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n834), .A2(new_n840), .B1(new_n923), .B2(new_n924), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT103), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT103), .B1(new_n841), .B2(new_n925), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n911), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n921), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(new_n926), .B2(new_n927), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n908), .A2(new_n909), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n910), .A2(new_n903), .ZN(new_n944));
  OAI22_X1  g519(.A1(new_n942), .A2(new_n936), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n945), .A2(new_n899), .A3(new_n931), .A4(new_n930), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n939), .A2(new_n940), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n942), .A2(new_n929), .A3(new_n936), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n910), .A2(new_n904), .A3(new_n907), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(new_n929), .B2(KEYINPUT41), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n951), .A2(new_n928), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n921), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n953), .A2(new_n946), .A3(new_n954), .A4(new_n879), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n948), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n946), .A3(new_n879), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n939), .A2(new_n954), .A3(new_n940), .A4(new_n946), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  MUX2_X1   g535(.A(new_n956), .B(new_n960), .S(KEYINPUT44), .Z(G397));
  XNOR2_X1  g536(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n962));
  AOI21_X1  g537(.A(G1384), .B1(new_n859), .B2(new_n860), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n962), .B1(new_n963), .B2(KEYINPUT105), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n861), .A2(KEYINPUT105), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n465), .A2(G40), .A3(new_n471), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n858), .B(G2067), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n723), .B(G1996), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n814), .A2(new_n816), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n814), .A2(new_n816), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n802), .A2(new_n805), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(KEYINPUT107), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n802), .A2(new_n805), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n969), .B1(KEYINPUT107), .B2(new_n976), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n970), .A2(new_n975), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1966), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n968), .B1(new_n963), .B2(KEYINPUT45), .ZN(new_n983));
  NOR3_X1   g558(.A1(G164), .A2(G1384), .A3(new_n962), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n465), .A2(G40), .A3(new_n471), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n963), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G2084), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n985), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(G8), .B1(new_n530), .B2(new_n531), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT120), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n996), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n992), .A2(G8), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n1000), .B2(new_n993), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n985), .B2(new_n991), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1003), .A2(new_n994), .A3(new_n998), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n995), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n962), .B1(G164), .B2(G1384), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n737), .A4(new_n968), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n861), .A2(new_n965), .A3(new_n987), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n990), .A2(new_n1011), .A3(new_n968), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT121), .B(G1961), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1007), .A2(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n861), .A2(new_n965), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n986), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1007), .A2(G2078), .ZN(new_n1018));
  INV_X1    g593(.A(new_n962), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n963), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G301), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(G1981), .B1(new_n582), .B2(new_n585), .ZN(new_n1023));
  OAI21_X1  g598(.A(G651), .B1(new_n578), .B2(new_n580), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT78), .ZN(new_n1025));
  INV_X1    g600(.A(G1981), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n581), .A4(new_n575), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(KEYINPUT49), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1002), .B1(new_n968), .B2(new_n963), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT110), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n1034), .B(KEYINPUT49), .C1(new_n1023), .C2(new_n1027), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1030), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1029), .B1(new_n1037), .B2(G288), .ZN(new_n1038));
  NAND2_X1  g613(.A1(KEYINPUT109), .A2(KEYINPUT52), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1039), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1029), .B(new_n1041), .C1(new_n1037), .C2(G288), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n1043));
  NAND3_X1  g618(.A1(G288), .A2(new_n1043), .A3(new_n1037), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1036), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(G166), .B2(new_n1002), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n988), .A2(new_n748), .A3(new_n990), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n986), .B1(new_n963), .B2(KEYINPUT45), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1971), .B1(new_n1052), .B2(new_n1008), .ZN(new_n1053));
  OAI211_X1 g628(.A(G8), .B(new_n1050), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1008), .A2(new_n1009), .A3(new_n968), .ZN(new_n1055));
  INV_X1    g630(.A(G1971), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n963), .A2(new_n987), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT50), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n963), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1058), .A2(new_n748), .A3(new_n1060), .A4(new_n968), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1002), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1054), .B1(new_n1062), .B2(new_n1050), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1046), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1006), .A2(new_n1022), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n575), .A2(new_n581), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1026), .B1(new_n1068), .B2(new_n1025), .ZN(new_n1069));
  AND4_X1   g644(.A1(new_n1026), .A2(new_n1025), .A3(new_n581), .A4(new_n575), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1032), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1034), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1031), .A2(KEYINPUT110), .A3(new_n1032), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1067), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n784), .A2(new_n1037), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1027), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT112), .B(new_n1027), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1029), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1054), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1036), .A2(new_n1045), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1082), .B1(new_n1036), .B2(new_n1045), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1081), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g661(.A(new_n1002), .B(G286), .C1(new_n985), .C2(new_n991), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT63), .B1(new_n1064), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(G8), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1047), .A2(KEYINPUT113), .A3(new_n1049), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1090), .B(G8), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1092), .A2(new_n1087), .A3(KEYINPUT63), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1046), .A2(KEYINPUT111), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1094), .B1(new_n1095), .B2(new_n1083), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1080), .B(new_n1086), .C1(new_n1088), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n968), .A2(new_n963), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT115), .B(KEYINPUT58), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(new_n781), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1055), .B2(G1996), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT59), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1102), .A2(new_n546), .A3(new_n1104), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1103), .A2(KEYINPUT59), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1102), .A2(new_n546), .B1(new_n1106), .B2(new_n1104), .ZN(new_n1107));
  AOI21_X1  g682(.A(G1348), .B1(new_n988), .B2(new_n990), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1098), .A2(G2067), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n609), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1105), .A2(new_n1107), .B1(new_n1111), .B2(KEYINPUT60), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n601), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1111), .A2(new_n1113), .A3(KEYINPUT60), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT117), .B(KEYINPUT61), .Z(new_n1115));
  INV_X1    g690(.A(G1956), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n968), .B1(new_n963), .B2(new_n987), .ZN(new_n1117));
  NOR3_X1   g692(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1052), .A2(new_n1008), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n560), .A2(new_n565), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1119), .A2(new_n1121), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1115), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1112), .A2(new_n1114), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT114), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1122), .A2(new_n1131), .A3(new_n1126), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1131), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1126), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1138), .A2(KEYINPUT61), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1128), .A2(KEYINPUT118), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1135), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1134), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1132), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(new_n1138), .A3(KEYINPUT61), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT119), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1130), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1110), .A2(new_n601), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1128), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n968), .B1(new_n964), .B2(new_n966), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT122), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1154), .B(new_n968), .C1(new_n964), .C2(new_n966), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1009), .A2(new_n1018), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1153), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(G301), .B1(new_n1158), .B2(new_n1014), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1010), .A2(new_n1007), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1160), .A2(new_n1021), .A3(new_n1161), .A4(G301), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT54), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1151), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1162), .A2(KEYINPUT54), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1156), .B1(new_n1152), .B2(KEYINPUT122), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1166), .B1(new_n1155), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1165), .B(KEYINPUT123), .C1(new_n1168), .C2(G301), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1164), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1022), .B1(new_n1168), .B2(G301), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1005), .B(new_n1064), .C1(new_n1171), .C2(KEYINPUT54), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1097), .B1(new_n1150), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1066), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI211_X1 g751(.A(KEYINPUT124), .B(new_n1097), .C1(new_n1150), .C2(new_n1173), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n981), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT48), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n969), .A2(new_n978), .A3(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n969), .A2(new_n978), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1181), .A2(KEYINPUT48), .ZN(new_n1182));
  AOI211_X1 g757(.A(new_n1180), .B(new_n1182), .C1(new_n970), .C2(new_n975), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n971), .A2(new_n723), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n970), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n969), .A2(G1996), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1186), .A2(KEYINPUT125), .A3(KEYINPUT46), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT125), .B1(new_n1186), .B2(KEYINPUT46), .ZN(new_n1188));
  OAI221_X1 g763(.A(new_n1185), .B1(KEYINPUT46), .B2(new_n1186), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT47), .Z(new_n1190));
  NAND2_X1  g765(.A1(new_n971), .A2(new_n972), .ZN(new_n1191));
  OAI22_X1  g766(.A1(new_n1191), .A2(new_n974), .B1(G2067), .B2(new_n765), .ZN(new_n1192));
  AOI211_X1 g767(.A(new_n1183), .B(new_n1190), .C1(new_n970), .C2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1178), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g769(.A1(new_n658), .A2(G319), .A3(new_n643), .ZN(new_n1196));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g772(.A1(new_n658), .A2(KEYINPUT126), .A3(G319), .A4(new_n643), .ZN(new_n1199));
  AND3_X1   g773(.A1(new_n1198), .A2(new_n690), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n884), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g775(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g776(.A(KEYINPUT127), .B1(new_n956), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n1204));
  AOI211_X1 g778(.A(new_n1204), .B(new_n1201), .C1(new_n948), .C2(new_n955), .ZN(new_n1205));
  NOR2_X1   g779(.A1(new_n1203), .A2(new_n1205), .ZN(G308));
  NAND2_X1  g780(.A1(new_n956), .A2(new_n1202), .ZN(G225));
endmodule


