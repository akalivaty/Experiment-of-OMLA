

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591;

  XNOR2_X1 U326 ( .A(KEYINPUT25), .B(KEYINPUT93), .ZN(n461) );
  XNOR2_X1 U327 ( .A(KEYINPUT119), .B(n452), .ZN(n567) );
  XOR2_X1 U328 ( .A(n470), .B(KEYINPUT28), .Z(n526) );
  XOR2_X1 U329 ( .A(KEYINPUT80), .B(KEYINPUT0), .Z(n294) );
  XNOR2_X1 U330 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n440) );
  XNOR2_X1 U331 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U332 ( .A(n462), .B(n461), .ZN(n465) );
  INV_X1 U333 ( .A(KEYINPUT94), .ZN(n468) );
  NOR2_X1 U334 ( .A1(n521), .A2(n532), .ZN(n448) );
  NOR2_X1 U335 ( .A1(n470), .A2(n573), .ZN(n450) );
  NOR2_X1 U336 ( .A1(n588), .A2(n476), .ZN(n477) );
  XNOR2_X1 U337 ( .A(n317), .B(n316), .ZN(n323) );
  XNOR2_X1 U338 ( .A(n323), .B(n322), .ZN(n327) );
  INV_X1 U339 ( .A(G190GAT), .ZN(n456) );
  XOR2_X1 U340 ( .A(n434), .B(n433), .Z(n546) );
  XOR2_X1 U341 ( .A(n327), .B(n367), .Z(n530) );
  XNOR2_X1 U342 ( .A(n456), .B(KEYINPUT58), .ZN(n457) );
  XNOR2_X1 U343 ( .A(n479), .B(G29GAT), .ZN(n480) );
  XNOR2_X1 U344 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n481), .B(n480), .ZN(G1328GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n296) );
  NAND2_X1 U347 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U349 ( .A(n297), .B(KEYINPUT69), .Z(n305) );
  XOR2_X1 U350 ( .A(G15GAT), .B(G113GAT), .Z(n299) );
  XNOR2_X1 U351 ( .A(G50GAT), .B(G36GAT), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U353 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n301) );
  XNOR2_X1 U354 ( .A(G197GAT), .B(G1GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U358 ( .A(G169GAT), .B(G8GAT), .Z(n368) );
  XOR2_X1 U359 ( .A(n306), .B(n368), .Z(n310) );
  XOR2_X1 U360 ( .A(G29GAT), .B(G43GAT), .Z(n308) );
  XNOR2_X1 U361 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n422) );
  XOR2_X1 U363 ( .A(G141GAT), .B(G22GAT), .Z(n343) );
  XNOR2_X1 U364 ( .A(n422), .B(n343), .ZN(n309) );
  XOR2_X1 U365 ( .A(n310), .B(n309), .Z(n575) );
  INV_X1 U366 ( .A(n575), .ZN(n552) );
  XOR2_X1 U367 ( .A(KEYINPUT20), .B(G190GAT), .Z(n312) );
  XOR2_X1 U368 ( .A(G120GAT), .B(G71GAT), .Z(n388) );
  XOR2_X1 U369 ( .A(G15GAT), .B(G127GAT), .Z(n395) );
  XNOR2_X1 U370 ( .A(n388), .B(n395), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U372 ( .A(n313), .B(G99GAT), .Z(n317) );
  XOR2_X1 U373 ( .A(G176GAT), .B(KEYINPUT84), .Z(n315) );
  XNOR2_X1 U374 ( .A(KEYINPUT82), .B(KEYINPUT81), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U376 ( .A(G113GAT), .B(G134GAT), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n294), .B(n318), .ZN(n357) );
  XNOR2_X1 U378 ( .A(n357), .B(G169GAT), .ZN(n320) );
  AND2_X1 U379 ( .A1(G227GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U381 ( .A(G43GAT), .B(n321), .ZN(n322) );
  XOR2_X1 U382 ( .A(KEYINPUT18), .B(KEYINPUT83), .Z(n325) );
  XNOR2_X1 U383 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U385 ( .A(KEYINPUT19), .B(n326), .Z(n367) );
  XNOR2_X1 U386 ( .A(G211GAT), .B(KEYINPUT87), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n328), .B(KEYINPUT21), .ZN(n329) );
  XOR2_X1 U388 ( .A(n329), .B(KEYINPUT88), .Z(n331) );
  XNOR2_X1 U389 ( .A(G197GAT), .B(G218GAT), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n375) );
  XNOR2_X1 U391 ( .A(G148GAT), .B(KEYINPUT72), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n332), .B(KEYINPUT71), .ZN(n333) );
  XOR2_X1 U393 ( .A(n333), .B(G204GAT), .Z(n335) );
  XNOR2_X1 U394 ( .A(G78GAT), .B(G106GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n381) );
  XNOR2_X1 U396 ( .A(n375), .B(n381), .ZN(n347) );
  XOR2_X1 U397 ( .A(KEYINPUT23), .B(KEYINPUT86), .Z(n337) );
  XNOR2_X1 U398 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U400 ( .A(G50GAT), .B(G162GAT), .Z(n426) );
  XOR2_X1 U401 ( .A(n338), .B(n426), .Z(n345) );
  XNOR2_X1 U402 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n339), .B(KEYINPUT2), .ZN(n356) );
  XOR2_X1 U404 ( .A(KEYINPUT85), .B(n356), .Z(n341) );
  NAND2_X1 U405 ( .A1(G228GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U406 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n470) );
  XOR2_X1 U410 ( .A(G57GAT), .B(KEYINPUT1), .Z(n349) );
  XNOR2_X1 U411 ( .A(G1GAT), .B(G148GAT), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n365) );
  XOR2_X1 U413 ( .A(G162GAT), .B(G127GAT), .Z(n351) );
  XNOR2_X1 U414 ( .A(G141GAT), .B(G120GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n353) );
  XOR2_X1 U416 ( .A(G29GAT), .B(G85GAT), .Z(n352) );
  XNOR2_X1 U417 ( .A(n353), .B(n352), .ZN(n361) );
  XNOR2_X1 U418 ( .A(KEYINPUT6), .B(KEYINPUT4), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n354), .B(KEYINPUT89), .ZN(n355) );
  XOR2_X1 U420 ( .A(n355), .B(KEYINPUT5), .Z(n359) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n363) );
  NAND2_X1 U424 ( .A1(G225GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n467) );
  INV_X1 U427 ( .A(n467), .ZN(n519) );
  XNOR2_X1 U428 ( .A(G176GAT), .B(G92GAT), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n366), .B(G64GAT), .ZN(n387) );
  XOR2_X1 U430 ( .A(G36GAT), .B(G190GAT), .Z(n425) );
  XOR2_X1 U431 ( .A(n387), .B(n425), .Z(n370) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U434 ( .A(KEYINPUT77), .B(KEYINPUT90), .Z(n372) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U437 ( .A(n374), .B(n373), .Z(n377) );
  XNOR2_X1 U438 ( .A(n375), .B(G204GAT), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n521) );
  XOR2_X1 U440 ( .A(KEYINPUT70), .B(KEYINPUT31), .Z(n379) );
  XNOR2_X1 U441 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n392) );
  XNOR2_X1 U444 ( .A(G99GAT), .B(G85GAT), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n382), .B(KEYINPUT73), .ZN(n421) );
  INV_X1 U446 ( .A(KEYINPUT74), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n421), .B(n383), .ZN(n385) );
  NAND2_X1 U448 ( .A1(G230GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U450 ( .A(n387), .B(n386), .Z(n390) );
  XOR2_X1 U451 ( .A(G57GAT), .B(KEYINPUT13), .Z(n396) );
  XNOR2_X1 U452 ( .A(n388), .B(n396), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n578) );
  XOR2_X1 U455 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n393) );
  XNOR2_X1 U456 ( .A(n578), .B(n393), .ZN(n539) );
  NAND2_X1 U457 ( .A1(n575), .A2(n539), .ZN(n394) );
  XNOR2_X1 U458 ( .A(KEYINPUT46), .B(n394), .ZN(n414) );
  XOR2_X1 U459 ( .A(n396), .B(n395), .Z(n398) );
  XNOR2_X1 U460 ( .A(G183GAT), .B(G71GAT), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U462 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n400) );
  XNOR2_X1 U463 ( .A(KEYINPUT14), .B(KEYINPUT78), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U465 ( .A(n402), .B(n401), .Z(n404) );
  XNOR2_X1 U466 ( .A(G22GAT), .B(G211GAT), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U468 ( .A(KEYINPUT15), .B(G64GAT), .Z(n406) );
  NAND2_X1 U469 ( .A1(G231GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n413) );
  XOR2_X1 U472 ( .A(G155GAT), .B(G78GAT), .Z(n410) );
  XNOR2_X1 U473 ( .A(G1GAT), .B(G8GAT), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n411), .B(KEYINPUT79), .ZN(n412) );
  XNOR2_X1 U476 ( .A(n413), .B(n412), .ZN(n583) );
  INV_X1 U477 ( .A(n583), .ZN(n568) );
  NAND2_X1 U478 ( .A1(n414), .A2(n568), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n415), .B(KEYINPUT109), .ZN(n435) );
  XOR2_X1 U480 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n417) );
  XNOR2_X1 U481 ( .A(KEYINPUT10), .B(KEYINPUT66), .ZN(n416) );
  XNOR2_X1 U482 ( .A(n417), .B(n416), .ZN(n434) );
  XOR2_X1 U483 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n419) );
  NAND2_X1 U484 ( .A1(G232GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U486 ( .A(n420), .B(KEYINPUT65), .Z(n424) );
  XNOR2_X1 U487 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U489 ( .A(G92GAT), .B(n425), .Z(n428) );
  XNOR2_X1 U490 ( .A(G106GAT), .B(n426), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U492 ( .A(n430), .B(n429), .Z(n432) );
  XNOR2_X1 U493 ( .A(G134GAT), .B(G218GAT), .ZN(n431) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n433) );
  INV_X1 U495 ( .A(n546), .ZN(n560) );
  NAND2_X1 U496 ( .A1(n435), .A2(n560), .ZN(n438) );
  XOR2_X1 U497 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n436) );
  XNOR2_X1 U498 ( .A(KEYINPUT47), .B(n436), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n445) );
  INV_X1 U500 ( .A(KEYINPUT36), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n439), .B(n546), .ZN(n588) );
  NOR2_X1 U502 ( .A1(n568), .A2(n588), .ZN(n441) );
  NAND2_X1 U503 ( .A1(n442), .A2(n552), .ZN(n443) );
  NOR2_X1 U504 ( .A1(n578), .A2(n443), .ZN(n444) );
  NOR2_X1 U505 ( .A1(n445), .A2(n444), .ZN(n446) );
  XNOR2_X1 U506 ( .A(n446), .B(KEYINPUT48), .ZN(n532) );
  XNOR2_X1 U507 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n449) );
  NAND2_X1 U509 ( .A1(n519), .A2(n449), .ZN(n573) );
  XNOR2_X1 U510 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NOR2_X1 U511 ( .A1(n530), .A2(n451), .ZN(n452) );
  NOR2_X1 U512 ( .A1(n552), .A2(n567), .ZN(n455) );
  INV_X1 U513 ( .A(G169GAT), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n453), .B(KEYINPUT120), .ZN(n454) );
  XNOR2_X1 U515 ( .A(n455), .B(n454), .ZN(G1348GAT) );
  NOR2_X1 U516 ( .A1(n560), .A2(n567), .ZN(n458) );
  NOR2_X1 U517 ( .A1(n521), .A2(n530), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n459), .B(KEYINPUT92), .ZN(n460) );
  NOR2_X1 U519 ( .A1(n470), .A2(n460), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n530), .A2(n470), .ZN(n463) );
  XOR2_X1 U521 ( .A(n463), .B(KEYINPUT26), .Z(n550) );
  INV_X1 U522 ( .A(n550), .ZN(n574) );
  XNOR2_X1 U523 ( .A(n521), .B(KEYINPUT27), .ZN(n471) );
  NOR2_X1 U524 ( .A1(n574), .A2(n471), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n475) );
  INV_X1 U528 ( .A(n526), .ZN(n536) );
  NOR2_X1 U529 ( .A1(n471), .A2(n519), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(KEYINPUT91), .ZN(n531) );
  NOR2_X1 U531 ( .A1(n536), .A2(n531), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n473), .A2(n530), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n475), .A2(n474), .ZN(n484) );
  NAND2_X1 U534 ( .A1(n568), .A2(n484), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT37), .B(n477), .Z(n518) );
  NOR2_X1 U536 ( .A1(n552), .A2(n578), .ZN(n485) );
  NAND2_X1 U537 ( .A1(n518), .A2(n485), .ZN(n478) );
  XNOR2_X1 U538 ( .A(KEYINPUT38), .B(n478), .ZN(n502) );
  NOR2_X1 U539 ( .A1(n519), .A2(n502), .ZN(n481) );
  XNOR2_X1 U540 ( .A(KEYINPUT39), .B(KEYINPUT98), .ZN(n479) );
  NAND2_X1 U541 ( .A1(n560), .A2(n583), .ZN(n482) );
  XOR2_X1 U542 ( .A(KEYINPUT16), .B(n482), .Z(n483) );
  AND2_X1 U543 ( .A1(n484), .A2(n483), .ZN(n505) );
  NAND2_X1 U544 ( .A1(n485), .A2(n505), .ZN(n494) );
  NOR2_X1 U545 ( .A1(n519), .A2(n494), .ZN(n487) );
  XNOR2_X1 U546 ( .A(KEYINPUT34), .B(KEYINPUT95), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NOR2_X1 U549 ( .A1(n521), .A2(n494), .ZN(n489) );
  XOR2_X1 U550 ( .A(KEYINPUT96), .B(n489), .Z(n490) );
  XNOR2_X1 U551 ( .A(G8GAT), .B(n490), .ZN(G1325GAT) );
  NOR2_X1 U552 ( .A1(n530), .A2(n494), .ZN(n492) );
  XNOR2_X1 U553 ( .A(KEYINPUT97), .B(KEYINPUT35), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U555 ( .A(G15GAT), .B(n493), .Z(G1326GAT) );
  NOR2_X1 U556 ( .A1(n526), .A2(n494), .ZN(n495) );
  XOR2_X1 U557 ( .A(G22GAT), .B(n495), .Z(G1327GAT) );
  NOR2_X1 U558 ( .A1(n521), .A2(n502), .ZN(n496) );
  XOR2_X1 U559 ( .A(G36GAT), .B(n496), .Z(G1329GAT) );
  NOR2_X1 U560 ( .A1(n502), .A2(n530), .ZN(n501) );
  XOR2_X1 U561 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n498) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(KEYINPUT100), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U564 ( .A(KEYINPUT99), .B(n499), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(G1330GAT) );
  NOR2_X1 U566 ( .A1(n526), .A2(n502), .ZN(n503) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  INV_X1 U568 ( .A(n539), .ZN(n562) );
  NOR2_X1 U569 ( .A1(n575), .A2(n562), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(KEYINPUT102), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n505), .A2(n517), .ZN(n512) );
  NOR2_X1 U572 ( .A1(n519), .A2(n512), .ZN(n506) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n506), .Z(n507) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n507), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n521), .A2(n512), .ZN(n508) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n508), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n530), .A2(n512), .ZN(n510) );
  XNOR2_X1 U578 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n509) );
  XNOR2_X1 U579 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n511), .ZN(G1334GAT) );
  NOR2_X1 U581 ( .A1(n512), .A2(n526), .ZN(n516) );
  XOR2_X1 U582 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n514) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT105), .ZN(n513) );
  XNOR2_X1 U584 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U585 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n518), .A2(n517), .ZN(n525) );
  NOR2_X1 U587 ( .A1(n519), .A2(n525), .ZN(n520) );
  XOR2_X1 U588 ( .A(G85GAT), .B(n520), .Z(G1336GAT) );
  NOR2_X1 U589 ( .A1(n521), .A2(n525), .ZN(n522) );
  XOR2_X1 U590 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  NOR2_X1 U591 ( .A1(n530), .A2(n525), .ZN(n524) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(KEYINPUT107), .ZN(n523) );
  XNOR2_X1 U593 ( .A(n524), .B(n523), .ZN(G1338GAT) );
  NOR2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U595 ( .A(KEYINPUT44), .B(KEYINPUT108), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U597 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  INV_X1 U598 ( .A(n530), .ZN(n533) );
  NOR2_X1 U599 ( .A1(n532), .A2(n531), .ZN(n551) );
  NAND2_X1 U600 ( .A1(n533), .A2(n551), .ZN(n534) );
  XOR2_X1 U601 ( .A(KEYINPUT113), .B(n534), .Z(n535) );
  NOR2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n575), .A2(n547), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(KEYINPUT114), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U607 ( .A1(n547), .A2(n539), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U609 ( .A1(n583), .A2(n547), .ZN(n545) );
  XOR2_X1 U610 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n543) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n559) );
  NOR2_X1 U618 ( .A1(n552), .A2(n559), .ZN(n553) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  NOR2_X1 U620 ( .A1(n562), .A2(n559), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n568), .A2(n559), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  NOR2_X1 U629 ( .A1(n567), .A2(n562), .ZN(n566) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n564) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT59), .B(n572), .Z(n577) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n586), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n586), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n582) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT124), .Z(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n586), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n585), .ZN(G1354GAT) );
  INV_X1 U651 ( .A(n586), .ZN(n587) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

