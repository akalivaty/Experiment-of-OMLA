//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n188), .A2(G227), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G107), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n192), .A2(G107), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n194), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n202), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n203), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n206));
  INV_X1    g020(.A(new_n200), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n195), .B1(new_n207), .B2(new_n197), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n208), .B(new_n193), .C1(new_n195), .C2(new_n197), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n206), .B1(new_n209), .B2(G101), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n204), .B1(new_n205), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT64), .A2(G143), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT64), .A2(G143), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n214), .B1(new_n217), .B2(G146), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT0), .A3(G128), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n212), .B1(new_n215), .B2(new_n216), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(G143), .B2(new_n212), .ZN(new_n222));
  XOR2_X1   g036(.A(KEYINPUT0), .B(G128), .Z(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n222), .A2(new_n226), .A3(new_n223), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n220), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT64), .B(G143), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n213), .B(new_n230), .C1(new_n231), .C2(new_n212), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n229), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(new_n218), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n193), .A2(KEYINPUT82), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT81), .B1(new_n192), .B2(G107), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n192), .A3(G107), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT81), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n196), .A3(G104), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n235), .A2(new_n236), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n241), .A2(KEYINPUT83), .A3(G101), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT83), .B1(new_n241), .B2(G101), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n234), .B(new_n205), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT10), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n211), .A2(new_n228), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n212), .A2(G143), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(new_n231), .B2(new_n212), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n229), .B1(new_n213), .B2(KEYINPUT1), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n232), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n232), .B(KEYINPUT70), .C1(new_n248), .C2(new_n249), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n252), .A2(KEYINPUT10), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n205), .B1(new_n242), .B2(new_n243), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT84), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n205), .B(KEYINPUT84), .C1(new_n242), .C2(new_n243), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n254), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT11), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(KEYINPUT66), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G137), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(KEYINPUT66), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(G137), .ZN(new_n266));
  INV_X1    g080(.A(G137), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G134), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT11), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n266), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(G131), .B1(new_n265), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n269), .A2(KEYINPUT11), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n270), .B1(new_n273), .B2(new_n268), .ZN(new_n274));
  INV_X1    g088(.A(G131), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n263), .A2(new_n261), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n274), .A2(new_n275), .A3(new_n266), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n246), .A2(new_n259), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n246), .B2(new_n259), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n191), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n246), .A2(new_n259), .A3(new_n279), .ZN(new_n283));
  INV_X1    g097(.A(new_n249), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n222), .A2(new_n284), .B1(new_n218), .B2(new_n230), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n255), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n244), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT12), .B1(new_n287), .B2(new_n278), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT12), .ZN(new_n289));
  AOI211_X1 g103(.A(new_n289), .B(new_n279), .C1(new_n286), .C2(new_n244), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n283), .B(new_n190), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n282), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G469), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n283), .B1(new_n288), .B2(new_n290), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n191), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n246), .A2(new_n259), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n278), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n283), .A3(new_n190), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n295), .B1(new_n301), .B2(new_n293), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT9), .B(G234), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(G116), .B(G119), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT5), .ZN(new_n308));
  INV_X1    g122(.A(G116), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n309), .A2(KEYINPUT5), .A3(G119), .ZN(new_n310));
  INV_X1    g124(.A(G113), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT2), .B(G113), .Z(new_n313));
  AOI22_X1  g127(.A1(new_n308), .A2(new_n312), .B1(new_n313), .B2(new_n307), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n257), .A2(new_n314), .A3(new_n258), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT69), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n307), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(new_n313), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n211), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G122), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n315), .A2(new_n320), .A3(new_n322), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(KEYINPUT6), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT85), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n228), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n227), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n226), .B1(new_n222), .B2(new_n223), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n219), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT85), .A3(G125), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n232), .B(new_n328), .C1(new_n248), .C2(new_n249), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT86), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n329), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n188), .A2(G224), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(KEYINPUT87), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n329), .A2(new_n338), .A3(new_n333), .A4(new_n335), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n321), .A2(new_n343), .A3(new_n323), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n326), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n334), .A2(KEYINPUT86), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n334), .A2(KEYINPUT86), .ZN(new_n347));
  OAI22_X1  g161(.A1(new_n228), .A2(new_n328), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n338), .A2(KEYINPUT7), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n255), .A2(new_n314), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n322), .B(KEYINPUT8), .Z(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(new_n255), .B2(new_n314), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n348), .A2(new_n349), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n349), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n329), .A2(new_n333), .A3(new_n335), .A4(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n325), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n356), .A2(new_n294), .ZN(new_n357));
  OAI21_X1  g171(.A(G210), .B1(G237), .B2(G902), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n345), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n345), .B2(new_n357), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(G214), .B1(G237), .B2(G902), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT89), .ZN(new_n365));
  INV_X1    g179(.A(G237), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n366), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n366), .A2(new_n188), .A3(G214), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n231), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G131), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT17), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n275), .B(new_n367), .C1(new_n231), .C2(new_n368), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G140), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G125), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n328), .A2(G140), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT16), .ZN(new_n377));
  OR3_X1    g191(.A1(new_n328), .A2(KEYINPUT16), .A3(G140), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n377), .A2(G146), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(G146), .B1(new_n377), .B2(new_n378), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n369), .A2(KEYINPUT17), .A3(G131), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n373), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G113), .B(G122), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(new_n192), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n375), .A2(new_n376), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT88), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G125), .B(G140), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT88), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n390), .A3(G146), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n386), .A2(G146), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n369), .ZN(new_n395));
  NAND2_X1  g209(.A1(KEYINPUT18), .A2(G131), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n369), .A2(KEYINPUT18), .A3(G131), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n383), .A2(new_n385), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT19), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n388), .B2(new_n390), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n389), .A2(KEYINPUT19), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n212), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n379), .B1(new_n370), .B2(new_n372), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n385), .B1(new_n407), .B2(new_n399), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n365), .B1(new_n401), .B2(new_n408), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n393), .A2(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n398), .A2(new_n410), .B1(new_n405), .B2(new_n406), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n400), .B(KEYINPUT89), .C1(new_n411), .C2(new_n385), .ZN(new_n412));
  NOR2_X1   g226(.A1(G475), .A2(G902), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT20), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n400), .B1(new_n411), .B2(new_n385), .ZN(new_n416));
  NOR3_X1   g230(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n385), .B1(new_n383), .B2(new_n399), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n401), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n294), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G475), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n188), .A2(G952), .ZN(new_n425));
  INV_X1    g239(.A(G234), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n425), .B1(new_n426), .B2(new_n366), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AOI211_X1 g242(.A(new_n294), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(G898), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n309), .A2(G122), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G122), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT14), .B1(new_n436), .B2(G116), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n433), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n434), .A2(KEYINPUT14), .ZN(new_n439));
  MUX2_X1   g253(.A(new_n438), .B(new_n433), .S(new_n439), .Z(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G107), .ZN(new_n441));
  OR2_X1    g255(.A1(KEYINPUT64), .A2(G143), .ZN(new_n442));
  NAND2_X1  g256(.A1(KEYINPUT64), .A2(G143), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(G128), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n229), .A2(G143), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G134), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(new_n262), .A3(new_n445), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n436), .A2(G116), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n434), .A3(new_n196), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n441), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT91), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT90), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n444), .A2(KEYINPUT13), .A3(new_n445), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT13), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n442), .A2(new_n456), .A3(G128), .A4(new_n443), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G134), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n454), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n457), .A2(G134), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n444), .A2(KEYINPUT13), .A3(new_n445), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(KEYINPUT90), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n450), .A2(new_n434), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G107), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n451), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n448), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n453), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  AOI211_X1 g283(.A(KEYINPUT91), .B(new_n467), .C1(new_n459), .C2(new_n462), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n452), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n303), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(G217), .A3(new_n188), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n455), .A2(new_n454), .A3(new_n458), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT90), .B1(new_n460), .B2(new_n461), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n468), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT91), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n463), .A2(new_n453), .A3(new_n468), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n473), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n452), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n474), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G478), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(KEYINPUT15), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(KEYINPUT93), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n474), .A2(new_n482), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(KEYINPUT93), .A3(new_n294), .ZN(new_n488));
  INV_X1    g302(.A(new_n485), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n483), .A2(KEYINPUT93), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n486), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n432), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n306), .A2(new_n364), .A3(new_n493), .A4(KEYINPUT94), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT94), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n302), .A2(new_n432), .A3(new_n492), .A4(new_n304), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n345), .A2(new_n357), .ZN(new_n497));
  INV_X1    g311(.A(new_n358), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n345), .A2(new_n357), .A3(new_n358), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n362), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n495), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT32), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n278), .B(new_n219), .C1(new_n330), .C2(new_n331), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n268), .A2(new_n266), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT67), .B1(new_n506), .B2(new_n275), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n268), .A2(new_n266), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT67), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(G131), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n277), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n252), .A2(new_n511), .A3(new_n253), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n505), .A2(new_n512), .A3(KEYINPUT30), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT71), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT68), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n511), .A2(new_n516), .A3(new_n250), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n277), .A2(new_n507), .A3(new_n510), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT68), .B1(new_n285), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n505), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n505), .A2(new_n512), .A3(KEYINPUT71), .A4(KEYINPUT30), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n515), .A2(new_n522), .A3(new_n319), .A4(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n505), .A2(new_n512), .A3(new_n318), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n366), .A2(new_n188), .A3(G210), .ZN(new_n526));
  XOR2_X1   g340(.A(new_n526), .B(KEYINPUT27), .Z(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT26), .B(G101), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n527), .B(new_n528), .Z(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n530), .A2(KEYINPUT31), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n524), .A2(new_n532), .A3(new_n525), .A4(new_n529), .ZN(new_n533));
  INV_X1    g347(.A(new_n529), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT28), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n520), .A2(new_n319), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(new_n525), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n525), .A2(new_n535), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n294), .B1(new_n531), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n504), .B1(new_n541), .B2(G472), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n530), .A2(KEYINPUT31), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n533), .A3(new_n539), .ZN(new_n544));
  INV_X1    g358(.A(G472), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n544), .A2(KEYINPUT32), .A3(new_n545), .A4(new_n294), .ZN(new_n546));
  OR3_X1    g360(.A1(new_n537), .A2(new_n534), .A3(new_n538), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n524), .A2(new_n525), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n534), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT29), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n505), .A2(new_n512), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n319), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n535), .B1(new_n553), .B2(new_n525), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT72), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT72), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n538), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n529), .A2(KEYINPUT29), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n294), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G472), .B1(new_n551), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n542), .A2(new_n546), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n229), .A2(G119), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n229), .A2(G119), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT24), .B(G110), .ZN(new_n567));
  OAI22_X1  g381(.A1(new_n379), .A2(new_n380), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G119), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT74), .B1(new_n569), .B2(G128), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n563), .B1(new_n570), .B2(KEYINPUT23), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT23), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n565), .A2(KEYINPUT74), .A3(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n571), .A2(KEYINPUT75), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT75), .B1(new_n571), .B2(new_n573), .ZN(new_n575));
  OAI21_X1  g389(.A(G110), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT76), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n570), .A2(KEYINPUT23), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n573), .A3(new_n564), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT75), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(KEYINPUT75), .A3(new_n573), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT76), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(G110), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n568), .B1(new_n577), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n571), .A2(new_n573), .ZN(new_n587));
  INV_X1    g401(.A(G110), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n587), .A2(new_n588), .B1(new_n566), .B2(new_n567), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n589), .A2(new_n392), .A3(new_n379), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT77), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT22), .B(G137), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n586), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n594), .ZN(new_n596));
  INV_X1    g410(.A(new_n568), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n584), .B1(new_n583), .B2(G110), .ZN(new_n598));
  AOI211_X1 g412(.A(KEYINPUT76), .B(new_n588), .C1(new_n581), .C2(new_n582), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n590), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n596), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(G217), .B1(new_n426), .B2(G902), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT73), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n594), .B1(new_n586), .B2(new_n590), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n600), .A2(new_n601), .A3(new_n596), .ZN(new_n611));
  AOI21_X1  g425(.A(G902), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(KEYINPUT79), .B(KEYINPUT25), .C1(new_n612), .C2(KEYINPUT78), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT25), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n294), .B1(new_n595), .B2(new_n602), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT79), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT78), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n616), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n613), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n609), .B1(new_n620), .B2(new_n606), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n494), .A2(new_n503), .A3(new_n562), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  NOR2_X1   g437(.A1(new_n545), .A2(KEYINPUT95), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n541), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n541), .A2(new_n624), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n306), .A2(new_n625), .A3(new_n621), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n431), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n501), .A2(new_n362), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n484), .A2(G902), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n633), .A2(KEYINPUT96), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(KEYINPUT96), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n487), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n474), .A2(new_n482), .A3(KEYINPUT96), .A4(new_n633), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n483), .A2(G478), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n424), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n630), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n628), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT97), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  AND2_X1   g459(.A1(new_n422), .A2(G475), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n414), .A2(KEYINPUT20), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(KEYINPUT98), .B2(new_n415), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n415), .A2(KEYINPUT98), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n492), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n630), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n628), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT99), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT35), .B(G107), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  AND2_X1   g471(.A1(new_n625), .A2(new_n626), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n620), .A2(new_n606), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n600), .A2(new_n601), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n596), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n608), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT100), .B1(new_n659), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT25), .B1(new_n612), .B2(KEYINPUT79), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT79), .B1(new_n612), .B2(KEYINPUT78), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n605), .B1(new_n669), .B2(new_n613), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n670), .A2(new_n671), .A3(new_n664), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n494), .A2(new_n503), .A3(new_n658), .A4(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n428), .B1(new_n429), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n650), .A2(new_n651), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n305), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n673), .A2(new_n681), .A3(new_n364), .A4(new_n562), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  XOR2_X1   g497(.A(new_n678), .B(KEYINPUT39), .Z(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n305), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT40), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n501), .B(KEYINPUT38), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n659), .A2(new_n665), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n553), .A2(new_n525), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n530), .B1(new_n529), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n294), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G472), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n542), .A2(new_n546), .A3(new_n695), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n414), .A2(KEYINPUT20), .B1(new_n416), .B2(new_n417), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n362), .B1(new_n697), .B2(new_n646), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n492), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n689), .A2(new_n691), .A3(new_n696), .A4(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n687), .B1(new_n688), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n688), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n217), .ZN(G45));
  OAI211_X1 g517(.A(new_n424), .B(new_n679), .C1(new_n638), .C2(new_n639), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n305), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n673), .A2(new_n364), .A3(new_n562), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  AOI21_X1  g521(.A(new_n293), .B1(new_n292), .B2(new_n294), .ZN(new_n708));
  AOI211_X1 g522(.A(G469), .B(G902), .C1(new_n282), .C2(new_n291), .ZN(new_n709));
  INV_X1    g523(.A(new_n304), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n641), .A2(new_n562), .A3(new_n621), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NAND4_X1  g528(.A1(new_n653), .A2(new_n562), .A3(new_n621), .A4(new_n711), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  AND3_X1   g530(.A1(new_n711), .A2(new_n492), .A3(new_n432), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n673), .A2(new_n717), .A3(new_n364), .A4(new_n562), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  NAND2_X1  g533(.A1(new_n292), .A2(new_n294), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G469), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n721), .A2(new_n629), .A3(new_n304), .A4(new_n295), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n485), .B1(new_n483), .B2(KEYINPUT93), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n487), .A2(new_n294), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT93), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n424), .A2(new_n727), .A3(new_n362), .A4(new_n486), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n722), .A2(new_n728), .A3(new_n361), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n541), .A2(G472), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n558), .A2(new_n534), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n543), .A3(new_n533), .ZN(new_n732));
  NOR2_X1   g546(.A1(G472), .A2(G902), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT102), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n621), .A2(new_n730), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n729), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n711), .A2(new_n699), .A3(new_n501), .A4(new_n629), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n621), .A2(new_n730), .A3(new_n735), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT103), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT104), .B(G122), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G24));
  NOR2_X1   g558(.A1(new_n708), .A2(new_n709), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n304), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n502), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n704), .ZN(new_n748));
  AOI22_X1  g562(.A1(G472), .A2(new_n541), .B1(new_n732), .B2(new_n734), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n747), .A2(new_n690), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  NAND3_X1  g565(.A1(new_n499), .A2(new_n362), .A3(new_n500), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n305), .A2(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n562), .A2(new_n753), .A3(new_n621), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(KEYINPUT42), .A3(new_n748), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n562), .A2(new_n753), .A3(new_n621), .A4(new_n748), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  INV_X1    g574(.A(new_n680), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  OR2_X1    g577(.A1(new_n638), .A2(new_n639), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n423), .A3(new_n419), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT43), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT106), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n658), .A2(new_n691), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n752), .B1(new_n769), .B2(KEYINPUT44), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(KEYINPUT44), .B2(new_n769), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n297), .A2(new_n300), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT45), .ZN(new_n773));
  OAI21_X1  g587(.A(G469), .B1(new_n773), .B2(G902), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n709), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(KEYINPUT46), .B2(new_n774), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n304), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n685), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT105), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n771), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  OAI21_X1  g595(.A(new_n777), .B1(KEYINPUT107), .B2(KEYINPUT47), .ZN(new_n782));
  AND2_X1   g596(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n542), .A2(new_n546), .A3(new_n561), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n752), .A2(new_n621), .A3(new_n704), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NOR3_X1   g602(.A1(new_n766), .A2(new_n427), .A3(new_n740), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n689), .A2(new_n362), .A3(new_n746), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n791), .B(KEYINPUT113), .Z(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n792), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(KEYINPUT114), .A3(new_n792), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  INV_X1    g614(.A(new_n752), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n708), .A2(new_n709), .A3(new_n304), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n801), .B(new_n789), .C1(new_n784), .C2(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n766), .A2(new_n427), .A3(new_n746), .A4(new_n752), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n749), .A2(new_n690), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n801), .A2(new_n428), .A3(new_n621), .A4(new_n711), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n696), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n764), .A2(new_n424), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n804), .A2(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  OR3_X1    g625(.A1(new_n799), .A2(new_n800), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n621), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n785), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n804), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT48), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n808), .A2(new_n424), .A3(new_n764), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n789), .A2(new_n747), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n425), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n800), .B1(new_n799), .B2(new_n811), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n812), .B(new_n819), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n659), .A2(KEYINPUT100), .A3(new_n665), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n671), .B1(new_n670), .B2(new_n664), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n364), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n785), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n828), .A2(new_n717), .B1(new_n738), .B2(new_n741), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n830), .A3(new_n712), .A4(new_n715), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n742), .A2(new_n712), .A3(new_n715), .A4(new_n718), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT112), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n825), .A2(new_n826), .A3(new_n492), .A4(new_n650), .ZN(new_n835));
  OAI22_X1  g649(.A1(new_n785), .A2(new_n835), .B1(new_n640), .B2(new_n805), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n305), .A2(new_n752), .A3(new_n678), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n762), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n640), .B1(new_n492), .B2(new_n424), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n364), .A2(new_n840), .A3(new_n629), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n627), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n622), .A3(new_n674), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT111), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n842), .A2(new_n674), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n836), .A2(new_n837), .B1(new_n754), .B2(new_n761), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT111), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n622), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n759), .A2(KEYINPUT53), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n834), .A2(new_n844), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n305), .A2(new_n678), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n728), .A2(new_n361), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n696), .A2(new_n851), .A3(new_n691), .A4(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n682), .A2(new_n706), .A3(new_n750), .A4(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(KEYINPUT108), .B(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT109), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(KEYINPUT109), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT110), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n854), .A2(KEYINPUT109), .A3(new_n855), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT109), .B1(new_n854), .B2(new_n855), .ZN(new_n865));
  OAI211_X1 g679(.A(KEYINPUT110), .B(new_n862), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n850), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n832), .A2(new_n843), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n759), .A2(new_n846), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n854), .B(new_n861), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT53), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT110), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n866), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n869), .A2(KEYINPUT53), .A3(new_n870), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n871), .A2(new_n872), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n881), .A2(new_n882), .B1(KEYINPUT53), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n824), .A2(new_n886), .B1(G952), .B2(G953), .ZN(new_n887));
  OR4_X1    g701(.A1(new_n363), .A2(new_n765), .A3(new_n813), .A4(new_n710), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n745), .B(KEYINPUT49), .Z(new_n889));
  OR4_X1    g703(.A1(new_n696), .A2(new_n888), .A3(new_n689), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n887), .A2(new_n890), .ZN(G75));
  NOR2_X1   g705(.A1(new_n188), .A2(G952), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n873), .B1(new_n881), .B2(new_n850), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n294), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(G210), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n326), .A2(new_n344), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(new_n342), .Z(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n893), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n896), .B2(new_n899), .ZN(G51));
  AND2_X1   g715(.A1(new_n876), .A2(KEYINPUT116), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n876), .A2(KEYINPUT116), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(G469), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT57), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n292), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n895), .A2(G469), .A3(new_n773), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n892), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND3_X1  g724(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n409), .A2(new_n412), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n893), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n913), .B1(new_n912), .B2(new_n911), .ZN(G60));
  AND2_X1   g728(.A1(new_n636), .A2(new_n637), .ZN(new_n915));
  XNOR2_X1  g729(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n916));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n905), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n877), .B2(new_n885), .ZN(new_n920));
  INV_X1    g734(.A(new_n915), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n893), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n919), .A2(new_n922), .ZN(G63));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT60), .Z(new_n927));
  AOI21_X1  g741(.A(new_n925), .B1(new_n875), .B2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n834), .A2(new_n844), .A3(new_n848), .A4(new_n849), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n880), .B2(new_n866), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n925), .B(new_n927), .C1(new_n930), .C2(new_n873), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n662), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n927), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT119), .B1(new_n894), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n935), .A2(new_n936), .A3(new_n603), .A4(new_n931), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n893), .A2(KEYINPUT61), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n933), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n935), .A2(new_n603), .A3(new_n931), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT121), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n924), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n935), .A2(new_n931), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n938), .B1(new_n944), .B2(new_n662), .ZN(new_n945));
  AND4_X1   g759(.A1(new_n924), .A2(new_n945), .A3(new_n942), .A4(new_n937), .ZN(new_n946));
  XOR2_X1   g760(.A(KEYINPUT118), .B(KEYINPUT61), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n941), .A2(new_n893), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n663), .B1(new_n935), .B2(new_n931), .ZN(new_n949));
  OAI211_X1 g763(.A(KEYINPUT120), .B(new_n947), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n933), .A2(new_n893), .A3(new_n941), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT120), .B1(new_n952), .B2(new_n947), .ZN(new_n953));
  OAI22_X1  g767(.A1(new_n943), .A2(new_n946), .B1(new_n951), .B2(new_n953), .ZN(G66));
  NAND2_X1  g768(.A1(G224), .A2(G953), .ZN(new_n955));
  OAI22_X1  g769(.A1(new_n869), .A2(G953), .B1(new_n430), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT123), .ZN(new_n957));
  INV_X1    g771(.A(G898), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n897), .B1(new_n958), .B2(G953), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(G69));
  NAND3_X1  g774(.A1(new_n515), .A2(new_n522), .A3(new_n523), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT124), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n403), .A2(new_n404), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n962), .B(new_n963), .Z(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(G227), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n188), .B1(new_n965), .B2(G900), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n682), .A2(new_n706), .A3(new_n750), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n702), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT62), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n814), .A2(new_n686), .A3(new_n801), .A4(new_n840), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n780), .A2(new_n787), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n964), .A2(G953), .ZN(new_n973));
  INV_X1    g787(.A(new_n968), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n787), .A2(new_n759), .A3(new_n762), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n814), .A2(new_n852), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n779), .B1(new_n771), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n188), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI22_X1  g792(.A1(new_n972), .A2(new_n973), .B1(new_n978), .B2(new_n964), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT125), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n967), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT126), .Z(G72));
  XNOR2_X1  g797(.A(new_n548), .B(new_n529), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT63), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n892), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n548), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n972), .A2(new_n988), .A3(new_n534), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n975), .A2(new_n977), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n548), .A2(new_n529), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n987), .B1(new_n992), .B2(new_n869), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n984), .A2(new_n986), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT127), .Z(new_n995));
  AOI21_X1  g809(.A(new_n993), .B1(new_n884), .B2(new_n995), .ZN(G57));
endmodule


