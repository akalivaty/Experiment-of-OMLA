

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n515), .A2(n519), .ZN(n875) );
  BUF_X1 U550 ( .A(n694), .Z(n512) );
  NOR2_X1 U551 ( .A1(n616), .A2(n529), .ZN(n643) );
  NOR2_X1 U552 ( .A1(G651), .A2(n616), .ZN(n638) );
  BUF_X1 U553 ( .A(n694), .Z(n511) );
  AND2_X1 U554 ( .A1(n963), .A2(n817), .ZN(n513) );
  OR2_X1 U555 ( .A1(n704), .A2(n703), .ZN(n705) );
  INV_X1 U556 ( .A(n941), .ZN(n753) );
  NOR2_X1 U557 ( .A1(n676), .A2(G1384), .ZN(n768) );
  NOR2_X2 U558 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  NOR2_X1 U559 ( .A1(n803), .A2(n513), .ZN(n804) );
  NOR2_X2 U560 ( .A1(G2105), .A2(n519), .ZN(n879) );
  AND2_X1 U561 ( .A1(G137), .A2(n880), .ZN(n523) );
  INV_X1 U562 ( .A(G2104), .ZN(n519) );
  NAND2_X1 U563 ( .A1(G101), .A2(n879), .ZN(n514) );
  XNOR2_X1 U564 ( .A(n514), .B(KEYINPUT23), .ZN(n518) );
  INV_X1 U565 ( .A(G2105), .ZN(n515) );
  NOR2_X1 U566 ( .A1(G2104), .A2(n515), .ZN(n537) );
  NAND2_X1 U567 ( .A1(G125), .A2(n537), .ZN(n516) );
  XOR2_X1 U568 ( .A(KEYINPUT64), .B(n516), .Z(n517) );
  NOR2_X1 U569 ( .A1(n518), .A2(n517), .ZN(n521) );
  NAND2_X1 U570 ( .A1(n875), .A2(G113), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n525) );
  XOR2_X2 U572 ( .A(KEYINPUT17), .B(n522), .Z(n880) );
  XOR2_X1 U573 ( .A(n523), .B(KEYINPUT65), .Z(n524) );
  NOR2_X2 U574 ( .A1(n525), .A2(n524), .ZN(G160) );
  NOR2_X1 U575 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U576 ( .A1(G90), .A2(n642), .ZN(n527) );
  XOR2_X1 U577 ( .A(KEYINPUT0), .B(G543), .Z(n616) );
  INV_X1 U578 ( .A(G651), .ZN(n529) );
  NAND2_X1 U579 ( .A1(G77), .A2(n643), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U581 ( .A(n528), .B(KEYINPUT9), .ZN(n532) );
  NOR2_X1 U582 ( .A1(G543), .A2(n529), .ZN(n530) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n530), .Z(n637) );
  NAND2_X1 U584 ( .A1(G64), .A2(n637), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n535) );
  NAND2_X1 U586 ( .A1(G52), .A2(n638), .ZN(n533) );
  XNOR2_X1 U587 ( .A(KEYINPUT67), .B(n533), .ZN(n534) );
  NOR2_X1 U588 ( .A1(n535), .A2(n534), .ZN(G171) );
  AND2_X1 U589 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U590 ( .A1(G138), .A2(n880), .ZN(n536) );
  XOR2_X1 U591 ( .A(n536), .B(KEYINPUT88), .Z(n543) );
  BUF_X1 U592 ( .A(n537), .Z(n876) );
  NAND2_X1 U593 ( .A1(n876), .A2(G126), .ZN(n541) );
  NAND2_X1 U594 ( .A1(G114), .A2(n875), .ZN(n539) );
  NAND2_X1 U595 ( .A1(G102), .A2(n879), .ZN(n538) );
  AND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n676) );
  BUF_X1 U599 ( .A(n676), .Z(G164) );
  INV_X1 U600 ( .A(G132), .ZN(G219) );
  INV_X1 U601 ( .A(G82), .ZN(G220) );
  INV_X1 U602 ( .A(G57), .ZN(G237) );
  INV_X1 U603 ( .A(G120), .ZN(G236) );
  INV_X1 U604 ( .A(G69), .ZN(G235) );
  NAND2_X1 U605 ( .A1(n642), .A2(G89), .ZN(n544) );
  XNOR2_X1 U606 ( .A(n544), .B(KEYINPUT4), .ZN(n546) );
  NAND2_X1 U607 ( .A1(G76), .A2(n643), .ZN(n545) );
  NAND2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U609 ( .A(KEYINPUT5), .B(n547), .ZN(n554) );
  XNOR2_X1 U610 ( .A(KEYINPUT74), .B(KEYINPUT6), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n638), .A2(G51), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n637), .A2(G63), .ZN(n548) );
  XOR2_X1 U613 ( .A(KEYINPUT73), .B(n548), .Z(n549) );
  NAND2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U615 ( .A(n552), .B(n551), .Z(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U617 ( .A(KEYINPUT7), .B(n555), .ZN(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n556) );
  XOR2_X1 U620 ( .A(n556), .B(KEYINPUT10), .Z(n822) );
  NAND2_X1 U621 ( .A1(n822), .A2(G567), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT11), .B(n557), .Z(G234) );
  NAND2_X1 U623 ( .A1(n637), .A2(G56), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT14), .ZN(n565) );
  XNOR2_X1 U625 ( .A(KEYINPUT13), .B(KEYINPUT68), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n642), .A2(G81), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(KEYINPUT12), .ZN(n561) );
  NAND2_X1 U628 ( .A1(G68), .A2(n643), .ZN(n560) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT69), .ZN(n568) );
  NAND2_X1 U633 ( .A1(G43), .A2(n638), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n956) );
  INV_X1 U635 ( .A(G860), .ZN(n613) );
  NOR2_X1 U636 ( .A1(n956), .A2(n613), .ZN(n569) );
  XOR2_X1 U637 ( .A(KEYINPUT70), .B(n569), .Z(G153) );
  XNOR2_X1 U638 ( .A(G171), .B(KEYINPUT71), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G868), .A2(G301), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G66), .A2(n637), .ZN(n571) );
  NAND2_X1 U641 ( .A1(G92), .A2(n642), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U643 ( .A1(G54), .A2(n638), .ZN(n573) );
  NAND2_X1 U644 ( .A1(G79), .A2(n643), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U647 ( .A(KEYINPUT72), .B(KEYINPUT15), .ZN(n576) );
  XOR2_X1 U648 ( .A(n577), .B(n576), .Z(n891) );
  INV_X1 U649 ( .A(n891), .ZN(n951) );
  INV_X1 U650 ( .A(G868), .ZN(n659) );
  NAND2_X1 U651 ( .A1(n951), .A2(n659), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(G284) );
  NAND2_X1 U653 ( .A1(G65), .A2(n637), .ZN(n581) );
  NAND2_X1 U654 ( .A1(G53), .A2(n638), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G91), .A2(n642), .ZN(n583) );
  NAND2_X1 U657 ( .A1(G78), .A2(n643), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n704) );
  INV_X1 U660 ( .A(n704), .ZN(G299) );
  NOR2_X1 U661 ( .A1(G286), .A2(n659), .ZN(n586) );
  XOR2_X1 U662 ( .A(KEYINPUT75), .B(n586), .Z(n588) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n587) );
  NOR2_X1 U664 ( .A1(n588), .A2(n587), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n613), .A2(G559), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n589), .A2(n891), .ZN(n590) );
  XNOR2_X1 U667 ( .A(n590), .B(KEYINPUT16), .ZN(n591) );
  XNOR2_X1 U668 ( .A(KEYINPUT76), .B(n591), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n956), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n891), .A2(G868), .ZN(n592) );
  NOR2_X1 U671 ( .A1(G559), .A2(n592), .ZN(n593) );
  NOR2_X1 U672 ( .A1(n594), .A2(n593), .ZN(G282) );
  NAND2_X1 U673 ( .A1(G111), .A2(n875), .ZN(n596) );
  NAND2_X1 U674 ( .A1(G99), .A2(n879), .ZN(n595) );
  NAND2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n604) );
  XOR2_X1 U676 ( .A(KEYINPUT18), .B(KEYINPUT78), .Z(n598) );
  NAND2_X1 U677 ( .A1(G123), .A2(n876), .ZN(n597) );
  XNOR2_X1 U678 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U679 ( .A(KEYINPUT77), .B(n599), .ZN(n601) );
  NAND2_X1 U680 ( .A1(n880), .A2(G135), .ZN(n600) );
  NAND2_X1 U681 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U682 ( .A(KEYINPUT79), .B(n602), .Z(n603) );
  NOR2_X1 U683 ( .A1(n604), .A2(n603), .ZN(n984) );
  XNOR2_X1 U684 ( .A(G2096), .B(n984), .ZN(n605) );
  INV_X1 U685 ( .A(G2100), .ZN(n830) );
  NAND2_X1 U686 ( .A1(n605), .A2(n830), .ZN(G156) );
  NAND2_X1 U687 ( .A1(G67), .A2(n637), .ZN(n607) );
  NAND2_X1 U688 ( .A1(G93), .A2(n642), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U690 ( .A1(G55), .A2(n638), .ZN(n609) );
  NAND2_X1 U691 ( .A1(G80), .A2(n643), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n658) );
  XOR2_X1 U694 ( .A(n658), .B(KEYINPUT80), .Z(n615) );
  NAND2_X1 U695 ( .A1(n891), .A2(G559), .ZN(n612) );
  XOR2_X1 U696 ( .A(n956), .B(n612), .Z(n656) );
  NAND2_X1 U697 ( .A1(n656), .A2(n613), .ZN(n614) );
  XNOR2_X1 U698 ( .A(n615), .B(n614), .ZN(G145) );
  NAND2_X1 U699 ( .A1(G49), .A2(n638), .ZN(n618) );
  NAND2_X1 U700 ( .A1(G87), .A2(n616), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U702 ( .A1(n637), .A2(n619), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n620) );
  XOR2_X1 U704 ( .A(KEYINPUT81), .B(n620), .Z(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(G288) );
  NAND2_X1 U706 ( .A1(G88), .A2(n642), .ZN(n624) );
  NAND2_X1 U707 ( .A1(G75), .A2(n643), .ZN(n623) );
  NAND2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n638), .A2(G50), .ZN(n625) );
  XOR2_X1 U710 ( .A(KEYINPUT82), .B(n625), .Z(n626) );
  NOR2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n637), .A2(G62), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(G303) );
  INV_X1 U714 ( .A(G303), .ZN(G166) );
  NAND2_X1 U715 ( .A1(G61), .A2(n637), .ZN(n631) );
  NAND2_X1 U716 ( .A1(G86), .A2(n642), .ZN(n630) );
  NAND2_X1 U717 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n643), .A2(G73), .ZN(n632) );
  XOR2_X1 U719 ( .A(KEYINPUT2), .B(n632), .Z(n633) );
  NOR2_X1 U720 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U721 ( .A1(n638), .A2(G48), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U723 ( .A1(G60), .A2(n637), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G47), .A2(n638), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U726 ( .A(KEYINPUT66), .B(n641), .Z(n647) );
  NAND2_X1 U727 ( .A1(G85), .A2(n642), .ZN(n645) );
  NAND2_X1 U728 ( .A1(G72), .A2(n643), .ZN(n644) );
  AND2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n647), .A2(n646), .ZN(G290) );
  XNOR2_X1 U731 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n649) );
  XNOR2_X1 U732 ( .A(G288), .B(KEYINPUT85), .ZN(n648) );
  XNOR2_X1 U733 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U734 ( .A(n650), .B(KEYINPUT83), .Z(n652) );
  XOR2_X1 U735 ( .A(G299), .B(n658), .Z(n651) );
  XNOR2_X1 U736 ( .A(n652), .B(n651), .ZN(n653) );
  XOR2_X1 U737 ( .A(n653), .B(G166), .Z(n654) );
  XNOR2_X1 U738 ( .A(n654), .B(G305), .ZN(n655) );
  XNOR2_X1 U739 ( .A(n655), .B(G290), .ZN(n890) );
  XOR2_X1 U740 ( .A(n890), .B(n656), .Z(n657) );
  NOR2_X1 U741 ( .A1(n659), .A2(n657), .ZN(n661) );
  AND2_X1 U742 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U743 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2084), .A2(G2078), .ZN(n662) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U748 ( .A1(n665), .A2(G2072), .ZN(n666) );
  XNOR2_X1 U749 ( .A(KEYINPUT86), .B(n666), .ZN(G158) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U751 ( .A1(G235), .A2(G236), .ZN(n667) );
  NAND2_X1 U752 ( .A1(G108), .A2(n667), .ZN(n668) );
  NOR2_X1 U753 ( .A1(n668), .A2(G237), .ZN(n669) );
  XNOR2_X1 U754 ( .A(n669), .B(KEYINPUT87), .ZN(n910) );
  NAND2_X1 U755 ( .A1(G567), .A2(n910), .ZN(n674) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U758 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U759 ( .A1(G96), .A2(n672), .ZN(n911) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n911), .ZN(n673) );
  NAND2_X1 U761 ( .A1(n674), .A2(n673), .ZN(n826) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U763 ( .A1(n826), .A2(n675), .ZN(n825) );
  NAND2_X1 U764 ( .A1(n825), .A2(G36), .ZN(G176) );
  INV_X1 U765 ( .A(n768), .ZN(n677) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n767) );
  NOR2_X2 U767 ( .A1(n677), .A2(n767), .ZN(n710) );
  INV_X1 U768 ( .A(n710), .ZN(n694) );
  INV_X1 U769 ( .A(n511), .ZN(n696) );
  NAND2_X1 U770 ( .A1(G8), .A2(n512), .ZN(n760) );
  NOR2_X1 U771 ( .A1(G1981), .A2(G305), .ZN(n678) );
  XOR2_X1 U772 ( .A(n678), .B(KEYINPUT24), .Z(n679) );
  NOR2_X1 U773 ( .A1(n760), .A2(n679), .ZN(n765) );
  NAND2_X1 U774 ( .A1(G1996), .A2(n710), .ZN(n680) );
  XOR2_X1 U775 ( .A(KEYINPUT26), .B(n680), .Z(n681) );
  NOR2_X2 U776 ( .A1(n681), .A2(n956), .ZN(n690) );
  NAND2_X1 U777 ( .A1(G1341), .A2(n511), .ZN(n689) );
  AND2_X1 U778 ( .A1(n891), .A2(n689), .ZN(n682) );
  AND2_X1 U779 ( .A1(n690), .A2(n682), .ZN(n683) );
  XNOR2_X1 U780 ( .A(n683), .B(KEYINPUT100), .ZN(n684) );
  INV_X1 U781 ( .A(n684), .ZN(n688) );
  NOR2_X1 U782 ( .A1(n696), .A2(G1348), .ZN(n686) );
  NOR2_X1 U783 ( .A1(G2067), .A2(n512), .ZN(n685) );
  NOR2_X1 U784 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U785 ( .A1(n688), .A2(n687), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U787 ( .A1(n951), .A2(n691), .ZN(n692) );
  NAND2_X1 U788 ( .A1(n693), .A2(n692), .ZN(n701) );
  NAND2_X1 U789 ( .A1(G1956), .A2(n512), .ZN(n695) );
  XNOR2_X1 U790 ( .A(KEYINPUT99), .B(n695), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n696), .A2(G2072), .ZN(n697) );
  XNOR2_X1 U792 ( .A(KEYINPUT27), .B(n697), .ZN(n698) );
  NOR2_X1 U793 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U796 ( .A(KEYINPUT101), .B(n702), .ZN(n707) );
  XOR2_X1 U797 ( .A(KEYINPUT28), .B(n705), .Z(n706) );
  NOR2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U799 ( .A(n708), .B(KEYINPUT29), .ZN(n714) );
  INV_X1 U800 ( .A(G1961), .ZN(n950) );
  NAND2_X1 U801 ( .A1(n512), .A2(n950), .ZN(n712) );
  XNOR2_X1 U802 ( .A(G2078), .B(KEYINPUT98), .ZN(n709) );
  XNOR2_X1 U803 ( .A(n709), .B(KEYINPUT25), .ZN(n1004) );
  NAND2_X1 U804 ( .A1(n710), .A2(n1004), .ZN(n711) );
  NAND2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U806 ( .A1(G171), .A2(n716), .ZN(n713) );
  NAND2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U808 ( .A(n715), .B(KEYINPUT102), .ZN(n736) );
  NOR2_X1 U809 ( .A1(G171), .A2(n716), .ZN(n721) );
  NOR2_X1 U810 ( .A1(G1966), .A2(n760), .ZN(n739) );
  NOR2_X1 U811 ( .A1(G2084), .A2(n512), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n739), .A2(n737), .ZN(n717) );
  NAND2_X1 U813 ( .A1(G8), .A2(n717), .ZN(n718) );
  XNOR2_X1 U814 ( .A(KEYINPUT30), .B(n718), .ZN(n719) );
  NOR2_X1 U815 ( .A1(G168), .A2(n719), .ZN(n720) );
  NOR2_X1 U816 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U817 ( .A(KEYINPUT31), .B(n722), .Z(n735) );
  INV_X1 U818 ( .A(G8), .ZN(n727) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n760), .ZN(n724) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n512), .ZN(n723) );
  NOR2_X1 U821 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U822 ( .A1(n725), .A2(G303), .ZN(n726) );
  OR2_X1 U823 ( .A1(n727), .A2(n726), .ZN(n729) );
  AND2_X1 U824 ( .A1(n735), .A2(n729), .ZN(n728) );
  NAND2_X1 U825 ( .A1(n736), .A2(n728), .ZN(n733) );
  INV_X1 U826 ( .A(n729), .ZN(n731) );
  AND2_X1 U827 ( .A1(G286), .A2(G8), .ZN(n730) );
  OR2_X1 U828 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U829 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U830 ( .A(n734), .B(KEYINPUT32), .ZN(n744) );
  AND2_X1 U831 ( .A1(n736), .A2(n735), .ZN(n742) );
  NAND2_X1 U832 ( .A1(G8), .A2(n737), .ZN(n738) );
  XNOR2_X1 U833 ( .A(KEYINPUT97), .B(n738), .ZN(n740) );
  OR2_X1 U834 ( .A1(n740), .A2(n739), .ZN(n741) );
  OR2_X1 U835 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n759) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n745) );
  NOR2_X1 U839 ( .A1(n751), .A2(n745), .ZN(n947) );
  NAND2_X1 U840 ( .A1(n759), .A2(n947), .ZN(n747) );
  NAND2_X1 U841 ( .A1(G288), .A2(G1976), .ZN(n746) );
  XOR2_X1 U842 ( .A(KEYINPUT103), .B(n746), .Z(n946) );
  NAND2_X1 U843 ( .A1(n747), .A2(n946), .ZN(n748) );
  NOR2_X1 U844 ( .A1(n760), .A2(n748), .ZN(n749) );
  NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n749), .ZN(n750) );
  INV_X1 U846 ( .A(n750), .ZN(n756) );
  NAND2_X1 U847 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U848 ( .A1(n760), .A2(n752), .ZN(n754) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n941) );
  NOR2_X1 U850 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U851 ( .A1(n756), .A2(n755), .ZN(n763) );
  NOR2_X1 U852 ( .A1(G2090), .A2(G303), .ZN(n757) );
  NAND2_X1 U853 ( .A1(G8), .A2(n757), .ZN(n758) );
  NAND2_X1 U854 ( .A1(n759), .A2(n758), .ZN(n761) );
  NAND2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n766) );
  INV_X1 U858 ( .A(n766), .ZN(n805) );
  NOR2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n817) );
  XOR2_X1 U860 ( .A(G2067), .B(KEYINPUT37), .Z(n769) );
  XOR2_X1 U861 ( .A(KEYINPUT90), .B(n769), .Z(n806) );
  NAND2_X1 U862 ( .A1(n876), .A2(G128), .ZN(n770) );
  XOR2_X1 U863 ( .A(KEYINPUT93), .B(n770), .Z(n772) );
  NAND2_X1 U864 ( .A1(n875), .A2(G116), .ZN(n771) );
  NAND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U866 ( .A(KEYINPUT35), .B(n773), .ZN(n780) );
  XNOR2_X1 U867 ( .A(KEYINPUT92), .B(KEYINPUT34), .ZN(n778) );
  NAND2_X1 U868 ( .A1(n880), .A2(G140), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n879), .A2(G104), .ZN(n774) );
  XOR2_X1 U870 ( .A(KEYINPUT91), .B(n774), .Z(n775) );
  NAND2_X1 U871 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U872 ( .A(n778), .B(n777), .Z(n779) );
  NAND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U874 ( .A(KEYINPUT36), .B(n781), .Z(n857) );
  NOR2_X1 U875 ( .A1(n806), .A2(n857), .ZN(n971) );
  NAND2_X1 U876 ( .A1(n817), .A2(n971), .ZN(n812) );
  INV_X1 U877 ( .A(n817), .ZN(n800) );
  NAND2_X1 U878 ( .A1(G117), .A2(n875), .ZN(n783) );
  NAND2_X1 U879 ( .A1(G129), .A2(n876), .ZN(n782) );
  NAND2_X1 U880 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U881 ( .A1(n879), .A2(G105), .ZN(n784) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U883 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U884 ( .A(n787), .B(KEYINPUT94), .ZN(n789) );
  NAND2_X1 U885 ( .A1(G141), .A2(n880), .ZN(n788) );
  NAND2_X1 U886 ( .A1(n789), .A2(n788), .ZN(n856) );
  NAND2_X1 U887 ( .A1(G1996), .A2(n856), .ZN(n790) );
  XOR2_X1 U888 ( .A(KEYINPUT95), .B(n790), .Z(n798) );
  NAND2_X1 U889 ( .A1(G107), .A2(n875), .ZN(n792) );
  NAND2_X1 U890 ( .A1(G95), .A2(n879), .ZN(n791) );
  NAND2_X1 U891 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U892 ( .A1(G119), .A2(n876), .ZN(n794) );
  NAND2_X1 U893 ( .A1(G131), .A2(n880), .ZN(n793) );
  NAND2_X1 U894 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U895 ( .A1(n796), .A2(n795), .ZN(n860) );
  NAND2_X1 U896 ( .A1(G1991), .A2(n860), .ZN(n797) );
  NAND2_X1 U897 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U898 ( .A(KEYINPUT96), .B(n799), .Z(n982) );
  NOR2_X1 U899 ( .A1(n800), .A2(n982), .ZN(n809) );
  INV_X1 U900 ( .A(n809), .ZN(n801) );
  NAND2_X1 U901 ( .A1(n812), .A2(n801), .ZN(n803) );
  XOR2_X1 U902 ( .A(G1986), .B(KEYINPUT89), .Z(n802) );
  XNOR2_X1 U903 ( .A(G290), .B(n802), .ZN(n963) );
  NAND2_X1 U904 ( .A1(n805), .A2(n804), .ZN(n820) );
  AND2_X1 U905 ( .A1(n857), .A2(n806), .ZN(n972) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n856), .ZN(n969) );
  NOR2_X1 U907 ( .A1(G1991), .A2(n860), .ZN(n985) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U909 ( .A1(n985), .A2(n807), .ZN(n808) );
  NOR2_X1 U910 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U911 ( .A1(n969), .A2(n810), .ZN(n811) );
  XNOR2_X1 U912 ( .A(n811), .B(KEYINPUT39), .ZN(n813) );
  NAND2_X1 U913 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U914 ( .A(KEYINPUT104), .B(n814), .Z(n815) );
  NOR2_X1 U915 ( .A1(n972), .A2(n815), .ZN(n816) );
  XNOR2_X1 U916 ( .A(KEYINPUT105), .B(n816), .ZN(n818) );
  NAND2_X1 U917 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U919 ( .A(KEYINPUT40), .B(n821), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n822), .ZN(G217) );
  INV_X1 U921 ( .A(n822), .ZN(G223) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U923 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U925 ( .A1(n825), .A2(n824), .ZN(G188) );
  XOR2_X1 U926 ( .A(KEYINPUT106), .B(n826), .Z(G319) );
  XNOR2_X1 U927 ( .A(G2067), .B(G2090), .ZN(n827) );
  XNOR2_X1 U928 ( .A(n827), .B(KEYINPUT42), .ZN(n838) );
  XOR2_X1 U929 ( .A(G2678), .B(KEYINPUT43), .Z(n829) );
  XNOR2_X1 U930 ( .A(KEYINPUT109), .B(G2096), .ZN(n828) );
  XNOR2_X1 U931 ( .A(n829), .B(n828), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n830), .B(G2072), .ZN(n832) );
  XNOR2_X1 U933 ( .A(G2084), .B(G2078), .ZN(n831) );
  XNOR2_X1 U934 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U935 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U936 ( .A(KEYINPUT108), .B(KEYINPUT107), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1981), .B(G1971), .Z(n840) );
  XNOR2_X1 U940 ( .A(G1966), .B(G1956), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n841), .B(KEYINPUT41), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U945 ( .A(G2474), .B(G1976), .Z(n845) );
  XOR2_X1 U946 ( .A(G1986), .B(n950), .Z(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U949 ( .A1(G124), .A2(n876), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n848), .B(KEYINPUT44), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n849), .B(KEYINPUT110), .ZN(n851) );
  NAND2_X1 U952 ( .A1(G112), .A2(n875), .ZN(n850) );
  NAND2_X1 U953 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U954 ( .A1(G100), .A2(n879), .ZN(n853) );
  NAND2_X1 U955 ( .A1(G136), .A2(n880), .ZN(n852) );
  NAND2_X1 U956 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U957 ( .A1(n855), .A2(n854), .ZN(G162) );
  XNOR2_X1 U958 ( .A(n856), .B(G162), .ZN(n859) );
  XOR2_X1 U959 ( .A(G164), .B(n857), .Z(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n864) );
  XNOR2_X1 U961 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n860), .B(KEYINPUT48), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U965 ( .A(G160), .B(n984), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n888) );
  NAND2_X1 U967 ( .A1(G103), .A2(n879), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G139), .A2(n880), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U970 ( .A(KEYINPUT112), .B(n869), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G115), .A2(n875), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G127), .A2(n876), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n975) );
  NAND2_X1 U976 ( .A1(G118), .A2(n875), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G130), .A2(n876), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U979 ( .A1(G106), .A2(n879), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G142), .A2(n880), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U984 ( .A(n975), .B(n886), .Z(n887) );
  XNOR2_X1 U985 ( .A(n888), .B(n887), .ZN(n889) );
  NOR2_X1 U986 ( .A1(G37), .A2(n889), .ZN(G395) );
  XOR2_X1 U987 ( .A(n890), .B(G286), .Z(n893) );
  XOR2_X1 U988 ( .A(G171), .B(n891), .Z(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U990 ( .A(n894), .B(n956), .Z(n895) );
  NOR2_X1 U991 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U992 ( .A(G2451), .B(G2430), .Z(n897) );
  XNOR2_X1 U993 ( .A(G2438), .B(G2443), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n903) );
  XOR2_X1 U995 ( .A(G2435), .B(G2454), .Z(n899) );
  XNOR2_X1 U996 ( .A(G1348), .B(G1341), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n901) );
  XOR2_X1 U998 ( .A(G2446), .B(G2427), .Z(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1000 ( .A(n903), .B(n902), .Z(n904) );
  NAND2_X1 U1001 ( .A1(G14), .A2(n904), .ZN(n912) );
  NAND2_X1 U1002 ( .A1(n912), .A2(G319), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(G225) );
  XNOR2_X1 U1008 ( .A(KEYINPUT113), .B(G225), .ZN(G308) );
  XOR2_X1 U1009 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  INV_X1 U1011 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1012 ( .A1(n911), .A2(n910), .ZN(G325) );
  INV_X1 U1013 ( .A(G325), .ZN(G261) );
  INV_X1 U1014 ( .A(n912), .ZN(G401) );
  XOR2_X1 U1015 ( .A(G1966), .B(G21), .Z(n924) );
  XNOR2_X1 U1016 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n913) );
  XNOR2_X1 U1017 ( .A(n913), .B(G4), .ZN(n914) );
  XNOR2_X1 U1018 ( .A(G1348), .B(n914), .ZN(n916) );
  XNOR2_X1 U1019 ( .A(G1956), .B(G20), .ZN(n915) );
  NOR2_X1 U1020 ( .A1(n916), .A2(n915), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(G1341), .B(G19), .ZN(n918) );
  XNOR2_X1 U1022 ( .A(G1981), .B(G6), .ZN(n917) );
  NOR2_X1 U1023 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1024 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1025 ( .A(KEYINPUT60), .B(n921), .Z(n922) );
  XNOR2_X1 U1026 ( .A(n922), .B(KEYINPUT126), .ZN(n923) );
  NAND2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1028 ( .A(n925), .B(KEYINPUT127), .ZN(n928) );
  XNOR2_X1 U1029 ( .A(G5), .B(KEYINPUT124), .ZN(n926) );
  XOR2_X1 U1030 ( .A(n926), .B(G1961), .Z(n927) );
  NAND2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(G1971), .B(G22), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(G23), .B(G1976), .ZN(n929) );
  NOR2_X1 U1034 ( .A1(n930), .A2(n929), .ZN(n932) );
  XOR2_X1 U1035 ( .A(G1986), .B(G24), .Z(n931) );
  NAND2_X1 U1036 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1037 ( .A(KEYINPUT58), .B(n933), .ZN(n934) );
  NOR2_X1 U1038 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1039 ( .A(n936), .B(KEYINPUT61), .ZN(n938) );
  XNOR2_X1 U1040 ( .A(G16), .B(KEYINPUT123), .ZN(n937) );
  NAND2_X1 U1041 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1042 ( .A1(G11), .A2(n939), .ZN(n967) );
  XOR2_X1 U1043 ( .A(G16), .B(KEYINPUT56), .Z(n965) );
  XOR2_X1 U1044 ( .A(G1966), .B(G168), .Z(n940) );
  XNOR2_X1 U1045 ( .A(KEYINPUT121), .B(n940), .ZN(n942) );
  NAND2_X1 U1046 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1047 ( .A(n943), .B(KEYINPUT57), .ZN(n961) );
  XOR2_X1 U1048 ( .A(G299), .B(G1956), .Z(n945) );
  NAND2_X1 U1049 ( .A1(G1971), .A2(G303), .ZN(n944) );
  NAND2_X1 U1050 ( .A1(n945), .A2(n944), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1052 ( .A1(n949), .A2(n948), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(G171), .B(n950), .ZN(n953) );
  XOR2_X1 U1054 ( .A(G1348), .B(n891), .Z(n952) );
  NOR2_X1 U1055 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1056 ( .A1(n955), .A2(n954), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(G1341), .B(n956), .ZN(n957) );
  XNOR2_X1 U1058 ( .A(KEYINPUT122), .B(n957), .ZN(n958) );
  NOR2_X1 U1059 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n995) );
  XOR2_X1 U1064 ( .A(G2090), .B(G162), .Z(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1066 ( .A(KEYINPUT51), .B(n970), .Z(n974) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n981) );
  XOR2_X1 U1069 ( .A(G2072), .B(n975), .Z(n977) );
  XOR2_X1 U1070 ( .A(G164), .B(G2078), .Z(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1072 ( .A(KEYINPUT116), .B(n978), .Z(n979) );
  XNOR2_X1 U1073 ( .A(KEYINPUT50), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n990) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(G160), .B(G2084), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1079 ( .A(KEYINPUT115), .B(n988), .Z(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(KEYINPUT52), .B(n991), .ZN(n992) );
  INV_X1 U1082 ( .A(KEYINPUT55), .ZN(n1016) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n1016), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n993), .A2(G29), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n1020) );
  XNOR2_X1 U1086 ( .A(G2067), .B(G26), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(G33), .B(G2072), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(G1996), .B(G32), .Z(n998) );
  NAND2_X1 U1090 ( .A1(n998), .A2(G28), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(G25), .B(G1991), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(KEYINPUT118), .B(n999), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(n1004), .B(G27), .Z(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT53), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(n1008), .B(KEYINPUT119), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(G2084), .B(G34), .Z(n1009) );
  XNOR2_X1 U1100 ( .A(KEYINPUT54), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(KEYINPUT117), .B(G2090), .Z(n1012) );
  XNOR2_X1 U1103 ( .A(G35), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1016), .B(n1015), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(G29), .A2(n1017), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(n1018), .B(KEYINPUT120), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1021), .Z(G150) );
  INV_X1 U1110 ( .A(G150), .ZN(G311) );
endmodule

