//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NOR2_X1   g0011(.A1(G58), .A2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n206), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n208), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n211), .B(new_n218), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n227), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT64), .ZN(new_n245));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n220), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n245), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n206), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  OAI22_X1  g0055(.A1(new_n201), .A2(new_n206), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n226), .A2(KEYINPUT66), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G58), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT8), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(new_n226), .B2(KEYINPUT8), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT8), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(KEYINPUT67), .A3(G58), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n260), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n206), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n256), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n216), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n246), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n269), .B(new_n216), .C1(G1), .C2(new_n206), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(new_n246), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G222), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G223), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n284), .B(new_n287), .C1(G77), .C2(new_n280), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT65), .B(G226), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  AND2_X1   g0093(.A1(G1), .A2(G13), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(new_n285), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  INV_X1    g0096(.A(G45), .ZN(new_n297));
  AOI21_X1  g0097(.A(G1), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n291), .A2(new_n292), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n288), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT68), .B(G179), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n288), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n279), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT9), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n279), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT70), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n300), .A2(G200), .ZN(new_n310));
  INV_X1    g0110(.A(G190), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n300), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT71), .B1(new_n279), .B2(new_n307), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT71), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n278), .A2(new_n314), .A3(KEYINPUT9), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n312), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n309), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n306), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT16), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT78), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT3), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT78), .A3(G33), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT7), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(G20), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n329), .B1(new_n280), .B2(G20), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n220), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G159), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT77), .B1(new_n254), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(G20), .A2(G33), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT77), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(G159), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n257), .A2(new_n259), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n212), .B1(new_n340), .B2(G68), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n339), .B1(new_n341), .B2(new_n206), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n322), .B1(new_n333), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT66), .B(G58), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n213), .B1(new_n344), .B2(new_n220), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(G20), .B1(new_n335), .B2(new_n338), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n326), .A2(G33), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n325), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT7), .B1(new_n348), .B2(new_n206), .ZN(new_n349));
  INV_X1    g0149(.A(new_n330), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n280), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(G68), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n346), .A2(new_n352), .A3(KEYINPUT16), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n343), .A2(new_n270), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT79), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT8), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n262), .A2(new_n264), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n276), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n260), .A2(new_n273), .A3(new_n262), .A4(new_n264), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(new_n359), .A3(new_n355), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OR2_X1    g0163(.A1(G223), .A2(G1698), .ZN(new_n364));
  INV_X1    g0164(.A(G226), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G1698), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n347), .A2(new_n364), .A3(new_n325), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G87), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n287), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n298), .A2(new_n286), .A3(G274), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n286), .A2(G232), .A3(new_n289), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n370), .A2(new_n311), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n286), .B1(new_n367), .B2(new_n368), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(new_n372), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n354), .A2(new_n363), .A3(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT17), .ZN(new_n381));
  INV_X1    g0181(.A(new_n303), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n370), .A2(new_n382), .A3(new_n373), .ZN(new_n383));
  OAI21_X1  g0183(.A(G169), .B1(new_n376), .B2(new_n377), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n383), .A2(KEYINPUT80), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT80), .B1(new_n383), .B2(new_n384), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n353), .A2(new_n270), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n331), .A2(new_n332), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G68), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT16), .B1(new_n390), .B2(new_n346), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n363), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n387), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n387), .B2(new_n392), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G244), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n371), .B1(new_n397), .B2(new_n290), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n280), .A2(G232), .A3(new_n282), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n280), .A2(G238), .A3(G1698), .ZN(new_n400));
  INV_X1    g0200(.A(G107), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n399), .B(new_n400), .C1(new_n401), .C2(new_n280), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n398), .B1(new_n402), .B2(new_n287), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT69), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  OAI21_X1  g0206(.A(G190), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n403), .A2(new_n404), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n403), .A2(new_n404), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(G200), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT8), .B(G58), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n411), .A2(new_n254), .B1(new_n206), .B2(new_n202), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n412), .B1(new_n267), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n271), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n274), .A2(new_n202), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n276), .B2(new_n202), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n407), .A2(new_n410), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n303), .B1(new_n405), .B2(new_n406), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n408), .A2(new_n301), .A3(new_n409), .ZN(new_n422));
  INV_X1    g0222(.A(new_n419), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AND4_X1   g0224(.A1(new_n381), .A2(new_n396), .A3(new_n420), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n336), .A2(G50), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT74), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n266), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n270), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT11), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n430), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n274), .A2(KEYINPUT12), .A3(new_n220), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT12), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n273), .B2(G68), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n433), .B(new_n435), .C1(new_n276), .C2(new_n220), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT75), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n436), .A2(KEYINPUT75), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n431), .A2(new_n432), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT72), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n282), .A2(G226), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n441), .B1(new_n348), .B2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n280), .A2(KEYINPUT72), .A3(G226), .A4(new_n282), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G97), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n443), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n447), .A2(new_n287), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n371), .B1(new_n221), .B2(new_n290), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT13), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n449), .B1(new_n447), .B2(new_n287), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT13), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n440), .B1(new_n454), .B2(G169), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n451), .A2(new_n452), .ZN(new_n456));
  AOI211_X1 g0256(.A(KEYINPUT13), .B(new_n449), .C1(new_n447), .C2(new_n287), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n440), .B(G169), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n450), .A2(G179), .A3(new_n453), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n439), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n439), .B1(new_n454), .B2(G200), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n456), .A2(new_n457), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT73), .B1(new_n463), .B2(G190), .ZN(new_n464));
  AND4_X1   g0264(.A1(KEYINPUT73), .A2(new_n450), .A3(G190), .A4(new_n453), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n466), .A3(KEYINPUT76), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n461), .A2(new_n466), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT76), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n321), .A2(new_n425), .A3(new_n467), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n397), .A2(G1698), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(G238), .B2(G1698), .ZN(new_n473));
  INV_X1    g0273(.A(G116), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n473), .A2(new_n348), .B1(new_n253), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n223), .B1(new_n297), .B2(G1), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n205), .A2(new_n293), .A3(G45), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n286), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT85), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT85), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n286), .A2(new_n476), .A3(new_n477), .A4(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n287), .A2(new_n475), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n303), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT19), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n206), .B1(new_n445), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G97), .A2(G107), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n222), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n347), .A2(new_n325), .A3(new_n206), .A4(G68), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n484), .B1(new_n266), .B2(new_n228), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n270), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n413), .A2(new_n274), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n205), .A2(G33), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n273), .A2(new_n494), .A3(new_n216), .A4(new_n269), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n492), .B(new_n493), .C1(new_n413), .C2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n483), .B(new_n496), .C1(G169), .C2(new_n482), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n475), .A2(new_n287), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n479), .A2(new_n481), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G200), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n482), .A2(G190), .ZN(new_n502));
  INV_X1    g0302(.A(new_n495), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G87), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n492), .A2(new_n504), .A3(new_n493), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n205), .B(G45), .C1(new_n296), .C2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT83), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G41), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n512), .A2(KEYINPUT83), .A3(new_n205), .A4(G45), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n511), .A2(G41), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n510), .A2(new_n513), .A3(new_n295), .A4(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(G257), .B(new_n286), .C1(new_n508), .C2(new_n514), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  AND2_X1   g0319(.A1(G250), .A2(G1698), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n397), .A2(G1698), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(KEYINPUT4), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n519), .B1(new_n522), .B2(new_n348), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT82), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT82), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT4), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n280), .B2(new_n521), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n287), .B1(new_n523), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n518), .A2(new_n530), .A3(new_n303), .ZN(new_n531));
  INV_X1    g0331(.A(new_n519), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G250), .A2(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n282), .A2(G244), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n524), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n535), .B2(new_n280), .ZN(new_n536));
  XNOR2_X1  g0336(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n348), .B2(new_n534), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n286), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n516), .A2(new_n517), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n301), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n531), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n274), .A2(KEYINPUT81), .A3(new_n228), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT81), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n273), .B2(G97), .ZN(new_n545));
  AOI22_X1  g0345(.A1(G97), .A2(new_n503), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  AND2_X1   g0348(.A1(G97), .A2(G107), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(new_n486), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n401), .A2(KEYINPUT6), .A3(G97), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(G20), .B1(G77), .B2(new_n336), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n326), .A2(G33), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n206), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n329), .A2(new_n556), .B1(new_n328), .B2(new_n330), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n553), .B1(new_n557), .B2(new_n401), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n547), .B1(new_n558), .B2(new_n270), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT84), .B1(new_n542), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n552), .A2(G20), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n336), .A2(G77), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n401), .B1(new_n331), .B2(new_n332), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n270), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n546), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT84), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(new_n531), .A4(new_n541), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n539), .A2(new_n540), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G190), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n559), .B(new_n570), .C1(new_n375), .C2(new_n569), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n507), .A2(new_n560), .A3(new_n568), .A4(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n222), .A2(KEYINPUT89), .A3(G20), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT22), .B1(new_n280), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(G33), .A2(G116), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n206), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n401), .A2(KEYINPUT23), .A3(G20), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT23), .B1(new_n401), .B2(G20), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n280), .A2(KEYINPUT22), .A3(new_n574), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n573), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT22), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT89), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n585), .A2(new_n206), .A3(G87), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n348), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT23), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n206), .B2(G107), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n401), .A2(KEYINPUT23), .A3(G20), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n589), .A2(new_n590), .B1(new_n206), .B2(new_n576), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n587), .A2(new_n573), .A3(new_n582), .A4(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n270), .B1(new_n583), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n274), .A2(KEYINPUT25), .A3(new_n401), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT25), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n273), .B2(G107), .ZN(new_n597));
  AOI22_X1  g0397(.A1(G107), .A2(new_n503), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(G264), .B(new_n286), .C1(new_n508), .C2(new_n514), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(G250), .A2(G1698), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n229), .B2(G1698), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n280), .ZN(new_n603));
  NAND2_X1  g0403(.A1(G33), .A2(G294), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n600), .B1(new_n605), .B2(new_n287), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(G190), .A3(new_n516), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n602), .A2(new_n280), .B1(G33), .B2(G294), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n516), .B(new_n599), .C1(new_n608), .C2(new_n286), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G200), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n594), .A2(new_n598), .A3(new_n607), .A4(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(G179), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n606), .A2(new_n612), .A3(new_n516), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(new_n301), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n587), .A2(new_n582), .A3(new_n591), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT24), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n271), .B1(new_n616), .B2(new_n592), .ZN(new_n617));
  INV_X1    g0417(.A(new_n598), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n613), .B(new_n614), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n519), .B(new_n206), .C1(G33), .C2(new_n228), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT20), .ZN(new_n622));
  AOI22_X1  g0422(.A1(KEYINPUT86), .A2(new_n622), .B1(new_n474), .B2(G20), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n623), .A3(new_n270), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n622), .A2(KEYINPUT86), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n625), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n621), .A2(new_n623), .A3(new_n627), .A4(new_n270), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n274), .A2(G116), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(G116), .B2(new_n495), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT87), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n273), .A2(new_n474), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n503), .B2(new_n474), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT87), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(new_n626), .A4(new_n628), .ZN(new_n636));
  INV_X1    g0436(.A(G303), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n348), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n282), .A2(G264), .ZN(new_n639));
  NOR2_X1   g0439(.A1(G257), .A2(G1698), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n347), .B(new_n325), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n641), .A3(new_n287), .ZN(new_n642));
  OAI211_X1 g0442(.A(G270), .B(new_n286), .C1(new_n508), .C2(new_n514), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n516), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G200), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n632), .A2(new_n636), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT88), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n644), .A2(new_n311), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n632), .A2(new_n636), .A3(new_n645), .A4(KEYINPUT88), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n644), .A2(G169), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n632), .B2(new_n636), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT21), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n632), .A2(new_n636), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n644), .A2(new_n612), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n653), .A2(KEYINPUT21), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n620), .A2(new_n651), .A3(new_n654), .A4(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n471), .A2(new_n572), .A3(new_n658), .ZN(G372));
  AND2_X1   g0459(.A1(new_n560), .A2(new_n568), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n660), .A2(new_n571), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT90), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n505), .A2(new_n662), .ZN(new_n663));
  AND4_X1   g0463(.A1(new_n662), .A2(new_n492), .A3(new_n504), .A4(new_n493), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n501), .B(new_n502), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n665), .A2(new_n497), .A3(new_n611), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n654), .A2(new_n657), .ZN(new_n667));
  XOR2_X1   g0467(.A(new_n619), .B(KEYINPUT91), .Z(new_n668));
  OAI211_X1 g0468(.A(new_n661), .B(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n542), .A2(new_n559), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n665), .A2(new_n497), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n497), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n560), .A2(new_n568), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n507), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n672), .B1(KEYINPUT26), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n471), .B1(new_n669), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n318), .A2(new_n320), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT17), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n380), .B(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n424), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n466), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n679), .B1(new_n681), .B2(new_n461), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n383), .A2(new_n384), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n354), .B2(new_n363), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(new_n393), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n677), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n305), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n676), .A2(new_n687), .ZN(G369));
  NAND2_X1  g0488(.A1(new_n611), .A2(new_n619), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(G213), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n594), .B2(new_n598), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n689), .A2(new_n697), .B1(new_n619), .B2(new_n696), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT92), .Z(new_n699));
  INV_X1    g0499(.A(new_n667), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n695), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n668), .A2(new_n696), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n655), .A2(new_n695), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n700), .A2(new_n651), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n700), .B2(new_n705), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n699), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n704), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n209), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n487), .A2(G116), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G1), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n214), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n700), .A2(new_n619), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n718), .A2(new_n661), .A3(new_n666), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n674), .A2(KEYINPUT26), .ZN(new_n720));
  INV_X1    g0520(.A(new_n497), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g0523(.A(KEYINPUT29), .B(new_n696), .C1(new_n719), .C2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n695), .B1(new_n675), .B2(new_n669), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(new_n725), .B2(KEYINPUT29), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n569), .B1(KEYINPUT93), .B2(new_n500), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n609), .A2(new_n303), .A3(new_n644), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n727), .B(new_n728), .C1(KEYINPUT93), .C2(new_n500), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n606), .A2(new_n482), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n569), .A4(new_n656), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n569), .A3(new_n656), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n729), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT31), .B1(new_n735), .B2(new_n695), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n658), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n572), .A2(new_n695), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT94), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n660), .A2(new_n507), .A3(new_n571), .A4(new_n696), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT94), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n743), .A2(new_n658), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n739), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G330), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n726), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n717), .B1(new_n749), .B2(G1), .ZN(G364));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n216), .B1(G20), .B2(new_n301), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n251), .A2(new_n297), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n711), .A2(new_n280), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n757), .B(new_n759), .C1(new_n297), .C2(new_n215), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n209), .A2(new_n280), .ZN(new_n761));
  INV_X1    g0561(.A(G355), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(G116), .B2(new_n209), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n760), .B1(KEYINPUT95), .B2(new_n763), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n763), .A2(KEYINPUT95), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n756), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G13), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n205), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n712), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n382), .A2(G20), .A3(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n206), .A2(G190), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(KEYINPUT32), .A3(G159), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT32), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n777), .B2(new_n334), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n774), .A2(G68), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n206), .B1(new_n776), .B2(G190), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n228), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n206), .A2(new_n311), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n375), .A2(G179), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n280), .B1(new_n787), .B2(new_n222), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n775), .A2(new_n786), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n784), .B(new_n788), .C1(G107), .C2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n382), .A2(new_n375), .A3(new_n785), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n382), .A2(new_n375), .A3(new_n775), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n793), .A2(new_n340), .B1(new_n795), .B2(G77), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n782), .A2(new_n791), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n773), .A2(new_n311), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n798), .A2(KEYINPUT96), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n773), .A2(KEYINPUT96), .A3(new_n311), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n797), .B1(G50), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT97), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(KEYINPUT97), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(G326), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT33), .B(G317), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n774), .A2(new_n807), .B1(new_n793), .B2(G322), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT98), .Z(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n794), .A2(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G283), .A2(new_n790), .B1(new_n778), .B2(G329), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n812), .B(new_n348), .C1(new_n637), .C2(new_n787), .ZN(new_n813));
  INV_X1    g0613(.A(new_n783), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n811), .B(new_n813), .C1(G294), .C2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n806), .A2(new_n809), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n804), .A2(new_n805), .A3(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n766), .B(new_n772), .C1(new_n817), .C2(new_n754), .ZN(new_n818));
  INV_X1    g0618(.A(new_n753), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n707), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n708), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n772), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n707), .A2(G330), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT99), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  INV_X1    g0626(.A(KEYINPUT101), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n424), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT101), .A4(new_n423), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n830), .A2(new_n420), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n725), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n423), .A2(new_n695), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n828), .A2(new_n420), .A3(new_n833), .A4(new_n829), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n680), .A2(new_n695), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n832), .B1(new_n725), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n771), .B1(new_n837), .B2(new_n747), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n747), .B2(new_n837), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n754), .A2(new_n751), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n771), .B1(G77), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n774), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n843), .A2(new_n844), .B1(new_n474), .B2(new_n794), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G294), .B2(new_n793), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n789), .A2(new_n222), .B1(new_n777), .B2(new_n810), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n348), .B1(new_n787), .B2(new_n401), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n847), .A2(new_n848), .A3(new_n784), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n846), .B(new_n849), .C1(new_n637), .C2(new_n801), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n774), .A2(G150), .B1(new_n795), .B2(G159), .ZN(new_n851));
  INV_X1    g0651(.A(G143), .ZN(new_n852));
  INV_X1    g0652(.A(G137), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n851), .B1(new_n852), .B2(new_n792), .C1(new_n801), .C2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT34), .Z(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n280), .B1(new_n777), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT100), .Z(new_n858));
  INV_X1    g0658(.A(new_n787), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G50), .A2(new_n859), .B1(new_n790), .B2(G68), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n858), .B(new_n860), .C1(new_n344), .C2(new_n783), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n850), .B1(new_n855), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n842), .B1(new_n862), .B2(new_n754), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n752), .B2(new_n836), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n839), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(G384));
  NAND2_X1  g0666(.A1(new_n552), .A2(KEYINPUT35), .ZN(new_n867));
  OAI211_X1 g0667(.A(G116), .B(new_n217), .C1(new_n552), .C2(KEYINPUT35), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT102), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT36), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n215), .B(G77), .C1(new_n220), .C2(new_n344), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n205), .B(G13), .C1(new_n873), .C2(new_n247), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(G330), .ZN(new_n876));
  INV_X1    g0676(.A(new_n471), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n746), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT105), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n354), .A2(new_n363), .A3(new_n379), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT103), .B1(new_n881), .B2(new_n684), .ZN(new_n882));
  INV_X1    g0682(.A(new_n693), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n392), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT103), .ZN(new_n885));
  INV_X1    g0685(.A(new_n362), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(new_n360), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n348), .A2(new_n330), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n220), .B1(new_n332), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n342), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n271), .B1(new_n890), .B2(KEYINPUT16), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n887), .B1(new_n891), .B2(new_n343), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n885), .B(new_n380), .C1(new_n892), .C2(new_n683), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n882), .A2(new_n884), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n392), .B1(new_n387), .B2(new_n883), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(KEYINPUT104), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n684), .B(KEYINPUT18), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n884), .B1(new_n901), .B2(new_n381), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n894), .A2(KEYINPUT37), .B1(new_n896), .B2(new_n897), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT104), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n880), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n322), .B1(new_n342), .B2(new_n889), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n353), .A3(new_n270), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n693), .B1(new_n909), .B2(new_n363), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n387), .A2(new_n392), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT18), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n387), .A2(new_n392), .A3(new_n393), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n910), .B1(new_n914), .B2(new_n679), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n909), .A2(new_n363), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n883), .ZN(new_n917));
  INV_X1    g0717(.A(new_n916), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n917), .B(new_n380), .C1(new_n918), .C2(new_n683), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n898), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n915), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n907), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n735), .A2(new_n695), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT31), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n736), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n744), .B1(new_n743), .B2(new_n658), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n740), .A2(new_n741), .A3(KEYINPUT94), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n439), .A2(new_n695), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n461), .A2(new_n466), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n931), .B1(new_n461), .B2(new_n466), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n836), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n930), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n917), .B1(new_n396), .B2(new_n381), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n919), .A2(KEYINPUT37), .B1(new_n896), .B2(new_n897), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n880), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n922), .ZN(new_n940));
  INV_X1    g0740(.A(new_n931), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n468), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n461), .A2(new_n466), .A3(new_n931), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n942), .A2(new_n943), .B1(new_n835), .B2(new_n834), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(new_n746), .A3(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n923), .A2(new_n936), .B1(new_n935), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n876), .B1(new_n879), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n879), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT106), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT39), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n923), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n461), .A2(new_n695), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n940), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT39), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n685), .A2(new_n693), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n830), .A2(new_n695), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n832), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n942), .A2(new_n943), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n956), .B(new_n957), .C1(new_n954), .C2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n726), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n687), .B1(new_n964), .B2(new_n877), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n963), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n949), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(G1), .B1(new_n767), .B2(G20), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n967), .A2(KEYINPUT107), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n949), .B2(new_n966), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT107), .B1(new_n967), .B2(new_n968), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n875), .B1(new_n970), .B2(new_n971), .ZN(G367));
  OR3_X1    g0772(.A1(new_n663), .A2(new_n664), .A3(new_n696), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(new_n497), .A3(new_n665), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n497), .B2(new_n973), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n661), .B1(new_n559), .B2(new_n696), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n670), .A2(new_n695), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n702), .A2(new_n980), .A3(KEYINPUT42), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n660), .B1(new_n980), .B2(new_n619), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n696), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT42), .B1(new_n702), .B2(new_n980), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT108), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n986), .B1(new_n985), .B2(new_n987), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n977), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n709), .A2(new_n980), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n985), .A2(new_n987), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT108), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(new_n976), .A3(new_n988), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n991), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n992), .B1(new_n991), .B2(new_n995), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n712), .B(KEYINPUT41), .Z(new_n999));
  OR2_X1    g0799(.A1(new_n699), .A2(new_n701), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n1000), .A2(KEYINPUT110), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n1001), .A2(new_n821), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n821), .ZN(new_n1003));
  OR3_X1    g0803(.A1(new_n1002), .A2(new_n1003), .A3(new_n702), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n702), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT44), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n980), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1007), .B1(new_n704), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n702), .A2(new_n703), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(KEYINPUT44), .A3(new_n980), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n704), .A2(KEYINPUT45), .A3(new_n1008), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n1010), .B2(new_n980), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(KEYINPUT109), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n709), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n709), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(KEYINPUT109), .A3(new_n1020), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1006), .A2(new_n1019), .A3(new_n749), .A4(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n999), .B1(new_n1022), .B2(new_n749), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n998), .B1(new_n1023), .B2(new_n770), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n758), .A2(new_n240), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n756), .B1(new_n711), .B2(new_n414), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n772), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n246), .A2(new_n794), .B1(new_n792), .B2(new_n255), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G159), .B2(new_n774), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n789), .A2(new_n202), .B1(new_n777), .B2(new_n853), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n280), .B1(new_n787), .B2(new_n344), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n783), .A2(new_n220), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1029), .B(new_n1033), .C1(new_n801), .C2(new_n852), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n859), .A2(G116), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT46), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1035), .A2(new_n1036), .B1(new_n401), .B2(new_n783), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n790), .A2(G97), .ZN(new_n1039));
  INV_X1    g0839(.A(G317), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n348), .C1(new_n1040), .C2(new_n777), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G283), .B2(new_n795), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n774), .A2(G294), .B1(new_n793), .B2(G303), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1038), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n801), .A2(new_n810), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1034), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT47), .Z(new_n1047));
  INV_X1    g0847(.A(new_n754), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1027), .B1(new_n975), .B2(new_n819), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT111), .Z(new_n1050));
  NAND2_X1  g0850(.A1(new_n1024), .A2(new_n1050), .ZN(G387));
  OAI22_X1  g0851(.A1(new_n761), .A2(new_n714), .B1(G107), .B2(new_n209), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n237), .A2(new_n297), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n714), .ZN(new_n1054));
  AOI211_X1 g0854(.A(G45), .B(new_n1054), .C1(G68), .C2(G77), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n411), .A2(G50), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n759), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1052), .B1(new_n1053), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n801), .A2(new_n334), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n793), .A2(G50), .B1(new_n795), .B2(G68), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n265), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1062), .B1(new_n1063), .B2(new_n843), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n783), .A2(new_n413), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n787), .A2(new_n202), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G150), .B2(new_n778), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n280), .A3(new_n1039), .ZN(new_n1068));
  NOR4_X1   g0868(.A1(new_n1061), .A2(new_n1064), .A3(new_n1065), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n774), .A2(G311), .B1(new_n795), .B2(G303), .ZN(new_n1070));
  XOR2_X1   g0870(.A(KEYINPUT113), .B(G322), .Z(new_n1071));
  OAI221_X1 g0871(.A(new_n1070), .B1(new_n1040), .B2(new_n792), .C1(new_n801), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n859), .A2(G294), .B1(new_n814), .B2(G283), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT49), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n280), .B1(new_n778), .B2(G326), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n474), .B2(new_n789), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1069), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n771), .B1(new_n756), .B2(new_n1060), .C1(new_n1084), .C2(new_n1048), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT114), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n699), .A2(new_n819), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1006), .A2(new_n770), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1006), .A2(new_n749), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n712), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1006), .A2(new_n749), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(G393));
  AOI21_X1  g0895(.A(new_n1017), .B1(KEYINPUT115), .B2(new_n1020), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(KEYINPUT115), .B2(new_n1020), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT115), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1017), .A2(new_n1098), .A3(new_n709), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1092), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(new_n712), .A3(new_n1022), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n801), .A2(new_n1040), .B1(new_n810), .B2(new_n792), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT52), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n348), .B1(new_n789), .B2(new_n401), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1071), .A2(new_n777), .B1(new_n787), .B2(new_n844), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(G116), .C2(new_n814), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n774), .A2(G303), .B1(new_n795), .B2(G294), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n801), .A2(new_n255), .B1(new_n334), .B2(new_n792), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT51), .Z(new_n1110));
  AOI22_X1  g0910(.A1(G68), .A2(new_n859), .B1(new_n778), .B2(G143), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1111), .B(new_n280), .C1(new_n222), .C2(new_n789), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n783), .A2(new_n202), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(new_n246), .B2(new_n843), .C1(new_n411), .C2(new_n794), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1108), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n754), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n755), .B1(new_n228), .B2(new_n209), .C1(new_n759), .C2(new_n244), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n771), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n753), .B2(new_n980), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n770), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1101), .A2(new_n1122), .ZN(G390));
  INV_X1    g0923(.A(new_n836), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n747), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n961), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n932), .A2(new_n933), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(KEYINPUT116), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT116), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n961), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n723), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n718), .A2(new_n661), .A3(new_n666), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n695), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n958), .B1(new_n1135), .B2(new_n831), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n923), .B(new_n952), .C1(new_n1132), .C2(new_n1136), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n951), .A2(new_n955), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n953), .B1(new_n960), .B2(new_n961), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1126), .B(new_n1137), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n747), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n951), .A2(new_n955), .B1(new_n962), .B2(new_n952), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1137), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1145), .A2(new_n769), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n802), .A2(G128), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n787), .A2(new_n255), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT53), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n843), .B2(new_n853), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n783), .A2(new_n334), .ZN(new_n1151));
  INV_X1    g0951(.A(G125), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n280), .B1(new_n777), .B2(new_n1152), .C1(new_n246), .C2(new_n789), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n856), .A2(new_n792), .B1(new_n794), .B2(new_n1154), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n802), .A2(G283), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n774), .A2(G107), .B1(new_n795), .B2(G97), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n474), .B2(new_n792), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G68), .A2(new_n790), .B1(new_n778), .B2(G294), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(new_n348), .C1(new_n222), .C2(new_n787), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1159), .A2(new_n1113), .A3(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1147), .A2(new_n1156), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n771), .B1(new_n265), .B2(new_n841), .C1(new_n1163), .C2(new_n1048), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1138), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n751), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1146), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1125), .A2(new_n961), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n960), .B1(new_n1168), .B2(new_n1141), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1126), .B(new_n1136), .C1(new_n1125), .C2(new_n1131), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n747), .A2(new_n471), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n965), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1145), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1173), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1140), .A2(new_n1177), .A3(new_n1144), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n712), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1167), .A2(new_n1179), .ZN(G378));
  OAI21_X1  g0980(.A(new_n957), .B1(new_n962), .B2(new_n954), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1138), .B2(new_n953), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n902), .B1(new_n899), .B2(KEYINPUT104), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n904), .A2(new_n905), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT38), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n922), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n936), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n876), .B1(new_n945), .B2(new_n935), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT119), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n677), .A2(new_n305), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n278), .A2(new_n693), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n321), .B1(new_n278), .B2(new_n693), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1196), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1190), .A2(new_n1191), .A3(new_n1200), .ZN(new_n1201));
  AND4_X1   g1001(.A1(new_n1189), .A2(new_n1200), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1182), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT120), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1191), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1190), .B1(new_n1191), .B2(new_n1200), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1208), .A2(new_n963), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1203), .A2(new_n1204), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1178), .A2(new_n1174), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1208), .A2(new_n963), .A3(new_n1209), .A4(KEYINPUT120), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT57), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1178), .B2(new_n1174), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1203), .A2(new_n1210), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n713), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1211), .A2(new_n770), .A3(new_n1213), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n772), .B1(new_n246), .B2(new_n840), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n843), .A2(new_n228), .B1(new_n413), .B2(new_n794), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G107), .B2(new_n793), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n789), .A2(new_n344), .B1(new_n777), .B2(new_n844), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n348), .A2(new_n296), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(new_n1225), .A2(new_n1066), .A3(new_n1032), .A4(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1224), .B(new_n1227), .C1(new_n474), .C2(new_n801), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT117), .ZN(new_n1229));
  XOR2_X1   g1029(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1226), .B(new_n246), .C1(G33), .C2(G41), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n787), .A2(new_n1154), .B1(new_n783), .B2(new_n255), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n795), .B2(G137), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n774), .A2(G132), .B1(new_n793), .B2(G128), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n801), .C2(new_n1152), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n790), .A2(G159), .ZN(new_n1240));
  AOI211_X1 g1040(.A(G33), .B(G41), .C1(new_n778), .C2(G124), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1232), .A2(new_n1233), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1229), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(new_n1230), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1222), .B1(new_n1048), .B2(new_n1245), .C1(new_n1207), .C2(new_n752), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1221), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1220), .A2(new_n1247), .ZN(G375));
  AND2_X1   g1048(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1132), .A2(new_n751), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT121), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n280), .B1(new_n783), .B2(new_n246), .C1(new_n344), .C2(new_n789), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G159), .A2(new_n859), .B1(new_n778), .B2(G128), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT122), .Z(new_n1254));
  OAI221_X1 g1054(.A(new_n1254), .B1(new_n255), .B2(new_n794), .C1(new_n843), .C2(new_n1154), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1252), .B(new_n1255), .C1(G137), .C2(new_n793), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n802), .A2(G132), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n774), .A2(G116), .B1(new_n795), .B2(G107), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n844), .B2(new_n792), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(G97), .A2(new_n859), .B1(new_n778), .B2(G303), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1260), .B(new_n348), .C1(new_n202), .C2(new_n789), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1259), .A2(new_n1065), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n802), .A2(G294), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1256), .A2(new_n1257), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n771), .B1(G68), .B2(new_n841), .C1(new_n1264), .C2(new_n1048), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n1249), .A2(new_n769), .B1(new_n1251), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1249), .A2(new_n1173), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1177), .A2(new_n999), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(G381));
  INV_X1    g1070(.A(G390), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1269), .A3(new_n1272), .ZN(new_n1273));
  OR4_X1    g1073(.A1(G387), .A2(new_n1273), .A3(G375), .A4(G378), .ZN(G407));
  INV_X1    g1074(.A(G378), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n694), .A2(G213), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n1276), .B(KEYINPUT123), .Z(new_n1277));
  NAND4_X1  g1077(.A1(new_n1220), .A2(new_n1275), .A3(new_n1247), .A4(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(G407), .A2(G213), .A3(new_n1278), .ZN(G409));
  XNOR2_X1  g1079(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1220), .A2(G378), .A3(new_n1247), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1218), .A2(new_n770), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1282), .B(new_n1246), .C1(new_n1214), .C2(new_n999), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1275), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1277), .B1(new_n1281), .B2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1249), .A2(KEYINPUT60), .A3(new_n1173), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n712), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1175), .A2(KEYINPUT60), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1287), .B1(new_n1267), .B2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n865), .B1(new_n1289), .B2(new_n1266), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1286), .A2(new_n712), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1267), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1266), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(G384), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1276), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1295), .A2(G2897), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1290), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1290), .A2(new_n1294), .B1(G2897), .B2(new_n1277), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1280), .B1(new_n1285), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT126), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1302), .A2(KEYINPUT62), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1285), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1295), .B(new_n1305), .C1(new_n1281), .C2(new_n1284), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1304), .B1(new_n1306), .B2(KEYINPUT62), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT126), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1308), .B(new_n1280), .C1(new_n1285), .C2(new_n1299), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1301), .A2(new_n1307), .A3(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT124), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(G387), .B2(new_n1271), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(G393), .B(G396), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(G390), .A2(new_n1024), .A3(new_n1050), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G390), .B1(new_n1024), .B2(new_n1050), .ZN(new_n1317));
  OAI22_X1  g1117(.A1(new_n1312), .A2(new_n1314), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G387), .A2(new_n1271), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1319), .A2(new_n1311), .A3(new_n1315), .A4(new_n1313), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1310), .A2(new_n1321), .ZN(new_n1322));
  OR2_X1    g1122(.A1(new_n1306), .A2(KEYINPUT63), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1324));
  OAI22_X1  g1124(.A1(new_n1324), .A2(new_n1295), .B1(new_n1298), .B2(new_n1297), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1302), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT61), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1323), .A2(new_n1325), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1322), .A2(new_n1328), .ZN(G405));
  XNOR2_X1  g1129(.A(G375), .B(G378), .ZN(new_n1330));
  OR2_X1    g1130(.A1(new_n1330), .A2(new_n1302), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT127), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1318), .A2(new_n1332), .A3(new_n1320), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1330), .A2(new_n1302), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1331), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1331), .A2(new_n1334), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1332), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1337));
  OR2_X1    g1137(.A1(new_n1333), .A2(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1335), .B1(new_n1336), .B2(new_n1338), .ZN(G402));
endmodule


