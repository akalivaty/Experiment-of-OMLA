//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n205), .A2(new_n208), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G169gat), .ZN(new_n219));
  INV_X1    g018(.A(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n216), .A2(new_n218), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT25), .B1(new_n213), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT23), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n217), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  OAI211_X1 g027(.A(KEYINPUT25), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n202), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n203), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G183gat), .B2(G190gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT67), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n203), .A2(new_n209), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n235), .A2(new_n236), .B1(new_n237), .B2(G190gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n229), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT68), .B1(new_n225), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n209), .A2(KEYINPUT27), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT27), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G183gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n243), .A3(new_n210), .ZN(new_n244));
  AND2_X1   g043(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n241), .A2(new_n243), .A3(new_n210), .A4(new_n246), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT26), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n221), .A2(new_n250), .A3(new_n222), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n228), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n248), .A2(new_n249), .A3(new_n251), .A4(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT70), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n251), .A2(new_n252), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n249), .A4(new_n248), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n211), .B(new_n212), .C1(new_n206), .C2(new_n207), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n223), .A2(new_n221), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT65), .B(G176gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n218), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n259), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n236), .A2(new_n235), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n233), .A2(new_n269), .A3(new_n212), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n259), .B1(new_n218), .B2(new_n220), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n240), .A2(new_n258), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G113gat), .B(G120gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(KEYINPUT1), .ZN(new_n276));
  XOR2_X1   g075(.A(G127gat), .B(G134gat), .Z(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G227gat), .ZN(new_n281));
  INV_X1    g080(.A(G233gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n240), .A2(new_n258), .A3(new_n273), .A4(new_n278), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G15gat), .B(G43gat), .Z(new_n289));
  XNOR2_X1  g088(.A(G71gat), .B(G99gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n284), .B1(new_n280), .B2(new_n285), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(KEYINPUT33), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n285), .ZN(new_n297));
  AOI221_X4 g096(.A(new_n294), .B1(KEYINPUT33), .B2(new_n291), .C1(new_n297), .C2(new_n283), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n288), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n267), .A2(new_n272), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n300), .A2(KEYINPUT68), .B1(new_n254), .B2(new_n257), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n278), .B1(new_n301), .B2(new_n273), .ZN(new_n302));
  INV_X1    g101(.A(new_n285), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n283), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT32), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT33), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n307), .A3(new_n291), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n295), .ZN(new_n309));
  INV_X1    g108(.A(new_n287), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n286), .B(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n299), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(KEYINPUT74), .B(new_n288), .C1(new_n296), .C2(new_n298), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n319), .B(new_n288), .C1(new_n296), .C2(new_n298), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n318), .A2(KEYINPUT36), .A3(new_n320), .A4(new_n312), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT31), .B(G50gat), .ZN(new_n323));
  INV_X1    g122(.A(G106gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G228gat), .A2(G233gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G211gat), .ZN(new_n329));
  INV_X1    g128(.A(G218gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G211gat), .A2(G218gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(KEYINPUT76), .A3(new_n332), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n332), .ZN(new_n339));
  AND2_X1   g138(.A1(G197gat), .A2(G204gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(G197gat), .A2(G204gat), .ZN(new_n341));
  OAI22_X1  g140(.A1(new_n339), .A2(KEYINPUT22), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n335), .A2(new_n336), .A3(new_n342), .A4(new_n337), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT3), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349));
  INV_X1    g148(.A(G155gat), .ZN(new_n350));
  INV_X1    g149(.A(G162gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n349), .B1(new_n352), .B2(KEYINPUT2), .ZN(new_n353));
  NAND2_X1  g152(.A1(G141gat), .A2(G148gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT82), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OR2_X1    g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT82), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n359), .A3(new_n354), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n353), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT83), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n353), .A2(new_n357), .A3(new_n360), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n352), .A2(new_n349), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT80), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n349), .A2(KEYINPUT2), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n367), .A2(KEYINPUT81), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(KEYINPUT81), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n368), .A2(new_n369), .A3(new_n358), .A4(new_n354), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n362), .A2(new_n364), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT84), .B(KEYINPUT3), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT29), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI221_X1 g172(.A(new_n328), .B1(new_n348), .B2(new_n371), .C1(new_n373), .C2(new_n346), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n327), .B(KEYINPUT87), .Z(new_n375));
  NAND2_X1  g174(.A1(new_n362), .A2(new_n364), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n366), .A2(new_n370), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(new_n372), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n346), .B1(new_n378), .B2(new_n347), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n342), .A2(KEYINPUT88), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381));
  OAI221_X1 g180(.A(new_n381), .B1(new_n340), .B2(new_n341), .C1(new_n339), .C2(KEYINPUT22), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n380), .A2(new_n382), .A3(new_n335), .A4(new_n337), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n335), .A2(new_n337), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(KEYINPUT88), .A3(new_n342), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n385), .A3(new_n347), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n371), .B1(new_n386), .B2(new_n372), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n375), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n374), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G22gat), .ZN(new_n390));
  INV_X1    g189(.A(G78gat), .ZN(new_n391));
  INV_X1    g190(.A(G22gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n392), .A3(new_n388), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n391), .B1(new_n390), .B2(new_n393), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n326), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(new_n393), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G78gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n325), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G1gat), .B(G29gat), .Z(new_n402));
  XNOR2_X1  g201(.A(G57gat), .B(G85gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT4), .B1(new_n371), .B2(new_n278), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n378), .B(new_n279), .C1(new_n409), .C2(new_n371), .ZN(new_n410));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n371), .A2(KEYINPUT4), .A3(new_n278), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n408), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT5), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n376), .A2(new_n377), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n279), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n371), .A2(new_n278), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n411), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n413), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n412), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n407), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n423), .A2(new_n414), .A3(new_n411), .A4(new_n410), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n406), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(new_n424), .A3(new_n406), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n427), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n425), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(KEYINPUT86), .A3(new_n427), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n428), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G226gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(new_n282), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n300), .A2(new_n253), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT77), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n300), .A2(KEYINPUT77), .A3(new_n253), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n436), .A2(KEYINPUT77), .A3(KEYINPUT29), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n440), .A2(new_n441), .B1(new_n274), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n346), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n438), .A2(new_n347), .A3(new_n437), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n240), .A2(new_n258), .A3(new_n273), .A4(new_n436), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(G8gat), .B(G36gat), .Z(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT78), .ZN(new_n451));
  XNOR2_X1  g250(.A(G64gat), .B(G92gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n449), .A4(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT79), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n448), .B1(new_n443), .B2(new_n444), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n453), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT30), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n401), .B1(new_n434), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n322), .A2(KEYINPUT89), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT89), .B1(new_n322), .B2(new_n462), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT92), .B(KEYINPUT37), .Z(new_n465));
  NAND2_X1  g264(.A1(new_n456), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n443), .A2(new_n346), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n446), .A2(new_n447), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n444), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(KEYINPUT37), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT38), .ZN(new_n471));
  INV_X1    g270(.A(new_n453), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n466), .A2(new_n470), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n453), .B1(new_n456), .B2(new_n465), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n476), .A2(KEYINPUT93), .A3(new_n471), .A4(new_n470), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n428), .ZN(new_n479));
  INV_X1    g278(.A(new_n458), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT37), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n466), .B(new_n472), .C1(new_n481), .C2(new_n456), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n480), .B1(new_n482), .B2(KEYINPUT38), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n425), .A2(KEYINPUT91), .ZN(new_n484));
  INV_X1    g283(.A(new_n430), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n425), .A2(KEYINPUT91), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n478), .A2(new_n479), .A3(new_n483), .A4(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n484), .A2(new_n486), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n408), .A2(new_n410), .A3(new_n412), .ZN(new_n490));
  XOR2_X1   g289(.A(KEYINPUT90), .B(KEYINPUT39), .Z(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n419), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n411), .B1(new_n423), .B2(new_n410), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT39), .B1(new_n418), .B2(new_n419), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n492), .B(new_n406), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT40), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n461), .A2(new_n489), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n401), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n488), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n463), .A2(new_n464), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n318), .A2(new_n320), .A3(new_n312), .ZN(new_n501));
  INV_X1    g300(.A(new_n434), .ZN(new_n502));
  INV_X1    g301(.A(new_n461), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n498), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n487), .A2(new_n479), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT35), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n455), .A2(new_n506), .A3(new_n460), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n505), .A2(new_n401), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n314), .A2(new_n315), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n504), .A2(KEYINPUT35), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n500), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n512));
  OR2_X1    g311(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n514));
  AOI21_X1  g313(.A(G36gat), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT14), .ZN(new_n516));
  INV_X1    g315(.A(G36gat), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n516), .A2(new_n517), .A3(G29gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G43gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(G50gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT94), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT15), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G50gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(G43gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n523), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n521), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n515), .A2(new_n518), .ZN(new_n532));
  INV_X1    g331(.A(new_n525), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n512), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n533), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n529), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n538), .A2(KEYINPUT17), .A3(new_n534), .A4(new_n521), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G8gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT16), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(G1gat), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n541), .B1(new_n544), .B2(KEYINPUT95), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(G1gat), .B2(new_n542), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI221_X1 g346(.A(new_n544), .B1(KEYINPUT95), .B2(new_n541), .C1(G1gat), .C2(new_n542), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n547), .A2(KEYINPUT96), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT96), .B1(new_n547), .B2(new_n548), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n540), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(new_n548), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n554), .A2(new_n534), .A3(new_n538), .A4(new_n521), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(KEYINPUT18), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G197gat), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT11), .B(G169gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT12), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n547), .A2(new_n548), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(new_n535), .B2(new_n531), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT98), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n567), .A3(new_n555), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n553), .B(KEYINPUT13), .Z(new_n569));
  NOR2_X1   g368(.A1(new_n531), .A2(new_n535), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(KEYINPUT98), .A3(new_n554), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n558), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n552), .A2(new_n553), .A3(new_n555), .A4(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n559), .A2(new_n564), .A3(new_n572), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT99), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n574), .A2(new_n572), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n577), .A2(new_n578), .A3(new_n564), .A4(new_n559), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n559), .ZN(new_n580));
  INV_X1    g379(.A(new_n564), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n576), .A2(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n511), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G71gat), .B(G78gat), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  INV_X1    g385(.A(G71gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n586), .B1(new_n587), .B2(new_n391), .ZN(new_n588));
  XOR2_X1   g387(.A(G57gat), .B(G64gat), .Z(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n588), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n584), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n565), .B1(new_n594), .B2(new_n593), .ZN(new_n602));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n602), .B(new_n605), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n601), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(KEYINPUT41), .ZN(new_n612));
  XNOR2_X1  g411(.A(G134gat), .B(G162gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G85gat), .A2(G92gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT7), .ZN(new_n618));
  NAND2_X1  g417(.A1(G99gat), .A2(G106gat), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  INV_X1    g419(.A(G92gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(KEYINPUT8), .A2(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G99gat), .B(G106gat), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(new_n618), .A3(new_n622), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n540), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n570), .A2(new_n630), .B1(KEYINPUT41), .B2(new_n611), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n616), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n629), .A2(new_n616), .A3(new_n631), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n614), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n614), .A3(new_n634), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n610), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n640), .B(KEYINPUT103), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n628), .A2(new_n593), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n625), .A2(new_n592), .A3(new_n590), .A4(new_n627), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n628), .A2(KEYINPUT102), .A3(new_n593), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT10), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n642), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n646), .A2(new_n641), .A3(new_n647), .ZN(new_n652));
  XOR2_X1   g451(.A(G120gat), .B(G148gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT104), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n651), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n656), .B1(new_n651), .B2(new_n652), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n639), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n583), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n502), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT105), .B(G1gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1324gat));
  NOR2_X1   g465(.A1(new_n663), .A2(new_n503), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n667), .A2(KEYINPUT106), .A3(new_n541), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT106), .B1(new_n667), .B2(new_n541), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n668), .B(new_n669), .C1(new_n672), .C2(new_n673), .ZN(G1325gat));
  INV_X1    g473(.A(G15gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n322), .A2(KEYINPUT108), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n317), .A2(new_n321), .A3(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n663), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n509), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n675), .B1(new_n663), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT107), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT107), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(G1326gat));
  NOR2_X1   g484(.A1(new_n663), .A2(new_n498), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT43), .B(G22gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  NOR3_X1   g487(.A1(new_n610), .A2(new_n661), .A3(new_n638), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n583), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n690), .A2(G29gat), .A3(new_n502), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(KEYINPUT45), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n660), .A2(KEYINPUT109), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n660), .A2(KEYINPUT109), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n696), .A2(new_n582), .A3(new_n610), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n638), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n500), .B2(new_n510), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT44), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n638), .B(KEYINPUT110), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n504), .A2(KEYINPUT35), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n508), .A2(new_n509), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n488), .A2(new_n497), .A3(new_n498), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n676), .A2(new_n708), .A3(new_n462), .A4(new_n678), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n704), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n698), .B1(new_n701), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G29gat), .B1(new_n713), .B2(new_n502), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n691), .A2(KEYINPUT45), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n692), .A2(new_n714), .A3(new_n715), .ZN(G1328gat));
  OAI21_X1  g515(.A(G36gat), .B1(new_n713), .B2(new_n503), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n583), .A2(new_n517), .A3(new_n461), .A4(new_n689), .ZN(new_n718));
  AND2_X1   g517(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n717), .B(new_n721), .C1(new_n719), .C2(new_n718), .ZN(G1329gat));
  NAND3_X1  g521(.A1(new_n583), .A2(new_n509), .A3(new_n689), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n723), .A2(new_n522), .B1(KEYINPUT112), .B2(KEYINPUT47), .ZN(new_n724));
  INV_X1    g523(.A(new_n679), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n712), .A2(G43gat), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n724), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n724), .B2(new_n726), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(G1330gat));
  NOR2_X1   g529(.A1(new_n498), .A2(new_n527), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n322), .A2(new_n462), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT89), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n708), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n707), .B1(new_n735), .B2(new_n463), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n703), .B1(new_n736), .B2(new_n699), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n697), .B(new_n731), .C1(new_n737), .C2(new_n710), .ZN(new_n738));
  INV_X1    g537(.A(new_n582), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n736), .A2(new_n739), .A3(new_n401), .A4(new_n689), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n527), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n743));
  NOR3_X1   g542(.A1(new_n742), .A2(KEYINPUT114), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT114), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n712), .A2(new_n731), .B1(new_n527), .B2(new_n740), .ZN(new_n746));
  INV_X1    g545(.A(new_n743), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n742), .A2(KEYINPUT48), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(G1331gat));
  NOR2_X1   g549(.A1(new_n639), .A2(new_n739), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n696), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT115), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n707), .A2(new_n709), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n434), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g557(.A(new_n503), .B(new_n755), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1333gat));
  NOR3_X1   g560(.A1(new_n755), .A2(G71gat), .A3(new_n681), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n756), .A2(new_n725), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(G71gat), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g564(.A1(new_n755), .A2(new_n498), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(new_n391), .ZN(G1335gat));
  NOR2_X1   g566(.A1(new_n739), .A2(new_n610), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n754), .A2(new_n699), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n754), .A2(KEYINPUT51), .A3(new_n699), .A4(new_n768), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n660), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n620), .A3(new_n434), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n710), .B1(new_n700), .B2(KEYINPUT44), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n768), .A2(new_n661), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT116), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779));
  INV_X1    g578(.A(new_n777), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n779), .B(new_n780), .C1(new_n737), .C2(new_n710), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n778), .A2(new_n434), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n775), .B1(new_n782), .B2(new_n620), .ZN(G1336gat));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n696), .A2(new_n621), .A3(new_n461), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n776), .A2(new_n503), .A3(new_n777), .ZN(new_n786));
  OAI221_X1 g585(.A(new_n784), .B1(new_n773), .B2(new_n785), .C1(new_n786), .C2(new_n621), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n785), .B1(new_n771), .B2(new_n772), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n778), .A2(new_n461), .A3(new_n781), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(G92gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n790), .B2(new_n784), .ZN(G1337gat));
  INV_X1    g590(.A(G99gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n774), .A2(new_n792), .A3(new_n509), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n778), .A2(new_n725), .A3(new_n781), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(new_n792), .ZN(G1338gat));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n796), .A2(KEYINPUT117), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n696), .A2(new_n324), .A3(new_n401), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n776), .A2(new_n498), .A3(new_n777), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(G106gat), .ZN(new_n800));
  OAI221_X1 g599(.A(new_n797), .B1(new_n773), .B2(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AOI211_X1 g600(.A(KEYINPUT117), .B(new_n798), .C1(new_n771), .C2(new_n772), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n778), .A2(new_n401), .A3(new_n781), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(G106gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n804), .B2(new_n796), .ZN(G1339gat));
  NAND2_X1  g604(.A1(new_n576), .A2(new_n579), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n553), .B1(new_n552), .B2(new_n555), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n569), .B1(new_n568), .B2(new_n571), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n563), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT118), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n811), .B(new_n563), .C1(new_n807), .C2(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n806), .A2(new_n661), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n646), .A2(new_n647), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n650), .B1(new_n816), .B2(new_n649), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n641), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n818), .A2(KEYINPUT54), .A3(new_n651), .ZN(new_n819));
  INV_X1    g618(.A(new_n656), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n651), .B2(KEYINPUT54), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n815), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n821), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(KEYINPUT54), .A3(new_n651), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n657), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n814), .B1(new_n582), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n638), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n822), .A2(new_n657), .A3(new_n825), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n576), .A2(new_n579), .B1(new_n810), .B2(new_n812), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n702), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n610), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n639), .A2(new_n739), .A3(new_n661), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n401), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n681), .A2(new_n502), .A3(new_n461), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n739), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n830), .A2(new_n834), .ZN(new_n843));
  INV_X1    g642(.A(new_n610), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n836), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n498), .A2(new_n501), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n502), .A2(new_n461), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n582), .A2(G113gat), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n842), .A2(G113gat), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT119), .ZN(G1340gat));
  AND3_X1   g652(.A1(new_n841), .A2(G120gat), .A3(new_n696), .ZN(new_n854));
  AOI21_X1  g653(.A(G120gat), .B1(new_n850), .B2(new_n661), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(G1341gat));
  OAI21_X1  g655(.A(G127gat), .B1(new_n840), .B2(new_n844), .ZN(new_n857));
  INV_X1    g656(.A(G127gat), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n850), .A2(new_n858), .A3(new_n610), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1342gat));
  INV_X1    g659(.A(G134gat), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n841), .B2(new_n699), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n850), .A2(new_n861), .A3(new_n699), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n863), .A2(new_n865), .A3(KEYINPUT120), .A4(new_n866), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1343gat));
  OAI21_X1  g670(.A(new_n401), .B1(new_n835), .B2(new_n836), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n679), .A2(new_n849), .ZN(new_n873));
  NOR4_X1   g672(.A1(new_n872), .A2(new_n873), .A3(G141gat), .A4(new_n582), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(KEYINPUT58), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n699), .B1(new_n827), .B2(KEYINPUT121), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n814), .B(new_n877), .C1(new_n582), .C2(new_n826), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n876), .A2(new_n878), .B1(new_n702), .B2(new_n833), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n846), .B1(new_n879), .B2(new_n610), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n401), .A2(KEYINPUT57), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n880), .A2(new_n882), .B1(new_n872), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n582), .A3(new_n873), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886));
  OAI21_X1  g685(.A(G141gat), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR4_X1   g686(.A1(new_n884), .A2(KEYINPUT123), .A3(new_n582), .A4(new_n873), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n875), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(new_n884), .B2(new_n873), .ZN(new_n891));
  INV_X1    g690(.A(new_n873), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n582), .A2(new_n826), .ZN(new_n893));
  AOI221_X4 g692(.A(new_n660), .B1(new_n810), .B2(new_n812), .C1(new_n576), .C2(new_n579), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT121), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n638), .A3(new_n878), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n834), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n844), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n881), .B1(new_n898), .B2(new_n846), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n847), .B2(new_n401), .ZN(new_n900));
  OAI211_X1 g699(.A(KEYINPUT122), .B(new_n892), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n891), .A2(new_n901), .A3(new_n739), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n874), .B1(new_n902), .B2(G141gat), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n889), .B1(new_n903), .B2(new_n904), .ZN(G1344gat));
  NAND3_X1  g704(.A1(new_n891), .A2(new_n901), .A3(new_n661), .ZN(new_n906));
  INV_X1    g705(.A(G148gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(KEYINPUT59), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n873), .A2(new_n660), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n831), .A2(new_n699), .A3(new_n832), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(new_n876), .B2(new_n878), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n846), .B1(new_n914), .B2(new_n610), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT57), .B1(new_n915), .B2(new_n401), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n881), .B1(new_n845), .B2(new_n846), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI211_X1 g717(.A(new_n910), .B(new_n911), .C1(new_n918), .C2(G148gat), .ZN(new_n919));
  INV_X1    g718(.A(new_n913), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n610), .B1(new_n896), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n401), .B1(new_n921), .B2(new_n836), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n917), .B1(new_n922), .B2(new_n883), .ZN(new_n923));
  INV_X1    g722(.A(new_n912), .ZN(new_n924));
  OAI21_X1  g723(.A(G148gat), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT124), .B1(new_n925), .B2(KEYINPUT59), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n909), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n872), .A2(new_n873), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n907), .A3(new_n661), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1345gat));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n350), .A3(new_n610), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n891), .A2(new_n901), .A3(new_n610), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n350), .ZN(G1346gat));
  NAND3_X1  g732(.A1(new_n928), .A2(new_n351), .A3(new_n699), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT125), .Z(new_n935));
  AND3_X1   g734(.A1(new_n891), .A2(new_n901), .A3(new_n702), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n351), .ZN(G1347gat));
  NOR2_X1   g736(.A1(new_n503), .A2(new_n434), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n847), .A2(new_n848), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(G169gat), .B1(new_n939), .B2(new_n739), .ZN(new_n940));
  AND4_X1   g739(.A1(new_n498), .A2(new_n847), .A3(new_n509), .A4(new_n938), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n582), .A2(new_n219), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(G1348gat));
  AOI21_X1  g742(.A(G176gat), .B1(new_n939), .B2(new_n661), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n695), .A2(new_n216), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n941), .B2(new_n945), .ZN(G1349gat));
  AOI21_X1  g745(.A(new_n209), .B1(new_n941), .B2(new_n610), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n610), .A2(new_n241), .A3(new_n243), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n939), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g748(.A(KEYINPUT126), .B(KEYINPUT60), .Z(new_n950));
  XNOR2_X1  g749(.A(new_n949), .B(new_n950), .ZN(G1350gat));
  AOI21_X1  g750(.A(new_n210), .B1(new_n941), .B2(new_n699), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT61), .Z(new_n953));
  NAND3_X1  g752(.A1(new_n939), .A2(new_n210), .A3(new_n702), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1351gat));
  INV_X1    g754(.A(new_n872), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n679), .A2(new_n938), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  XOR2_X1   g758(.A(KEYINPUT127), .B(G197gat), .Z(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n739), .A3(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(new_n923), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(new_n957), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(new_n582), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n964), .B2(new_n960), .ZN(G1352gat));
  NOR3_X1   g764(.A1(new_n958), .A2(G204gat), .A3(new_n660), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT62), .ZN(new_n967));
  OAI21_X1  g766(.A(G204gat), .B1(new_n963), .B2(new_n695), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1353gat));
  NAND3_X1  g768(.A1(new_n959), .A2(new_n329), .A3(new_n610), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n962), .A2(new_n610), .A3(new_n957), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  OAI21_X1  g773(.A(G218gat), .B1(new_n963), .B2(new_n638), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n330), .A3(new_n702), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1355gat));
endmodule


