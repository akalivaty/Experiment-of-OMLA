//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  AOI21_X1  g006(.A(G143), .B1(new_n190), .B2(G214), .ZN(new_n193));
  OAI21_X1  g007(.A(G131), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G214), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(new_n191), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT17), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT94), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n206), .B1(new_n210), .B2(new_n204), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n211), .B(G146), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n194), .A2(new_n199), .A3(KEYINPUT94), .A4(new_n200), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n197), .A2(new_n191), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT17), .A3(G131), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n203), .A2(new_n212), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G113), .B(G122), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n192), .A2(new_n193), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT18), .A2(G131), .ZN(new_n221));
  XNOR2_X1  g035(.A(G125), .B(G140), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n210), .A2(G146), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n220), .A2(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n214), .A2(KEYINPUT18), .A3(G131), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n216), .A2(new_n219), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n219), .B1(new_n216), .B2(new_n228), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n189), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G475), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT19), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n210), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n222), .A2(KEYINPUT19), .ZN(new_n236));
  AOI21_X1  g050(.A(G146), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI211_X1 g051(.A(G146), .B(new_n206), .C1(new_n210), .C2(new_n204), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n194), .A2(new_n199), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n240), .A2(new_n241), .B1(new_n226), .B2(new_n227), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT93), .B1(new_n242), .B2(new_n219), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n235), .A2(new_n236), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n241), .B(new_n238), .C1(G146), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n228), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT93), .ZN(new_n247));
  INV_X1    g061(.A(new_n219), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n229), .A2(new_n243), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G475), .A2(G902), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT20), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT20), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n250), .B2(new_n251), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n233), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G952), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(G234), .B2(G237), .ZN(new_n259));
  AOI211_X1 g073(.A(new_n189), .B(new_n257), .C1(G234), .C2(G237), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT21), .B(G898), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G128), .B(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT13), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n265), .A2(KEYINPUT13), .A3(G143), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n264), .A2(new_n268), .B1(new_n267), .B2(new_n263), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT68), .B(G116), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G122), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT95), .B(G122), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G116), .ZN(new_n273));
  INV_X1    g087(.A(G107), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n271), .B2(new_n273), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n269), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n263), .B(G134), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT96), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n263), .B(new_n267), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT96), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n283), .A3(new_n275), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n271), .A2(KEYINPUT14), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n271), .A2(KEYINPUT14), .B1(G116), .B2(new_n272), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n274), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n278), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT76), .B(G217), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT9), .B(G234), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n289), .A2(new_n290), .A3(G953), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n291), .B(new_n278), .C1(new_n284), .C2(new_n287), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n189), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT15), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(G478), .ZN(new_n298));
  INV_X1    g112(.A(G478), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n295), .B(new_n189), .C1(KEYINPUT15), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OR3_X1    g115(.A1(new_n256), .A2(new_n262), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G113), .ZN(new_n303));
  INV_X1    g117(.A(G116), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(G119), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(KEYINPUT68), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT68), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G116), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n310), .A3(G119), .ZN(new_n311));
  INV_X1    g125(.A(new_n305), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n307), .B1(new_n313), .B2(new_n306), .ZN(new_n314));
  NAND2_X1  g128(.A1(KEYINPUT2), .A2(G113), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT2), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(new_n303), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND4_X1   g135(.A1(KEYINPUT69), .A2(new_n321), .A3(new_n312), .A4(new_n311), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n305), .B1(new_n270), .B2(G119), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT69), .B1(new_n323), .B2(new_n321), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n314), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n274), .A2(G104), .ZN(new_n326));
  AND2_X1   g140(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n327));
  NOR2_X1   g141(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G101), .ZN(new_n330));
  XNOR2_X1  g144(.A(G104), .B(G107), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n329), .B(new_n330), .C1(new_n327), .C2(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n331), .A2(new_n330), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n325), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT69), .ZN(new_n336));
  INV_X1    g150(.A(new_n320), .ZN(new_n337));
  NOR3_X1   g151(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n315), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n336), .B1(new_n313), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n323), .A2(KEYINPUT69), .A3(new_n321), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n323), .A2(KEYINPUT5), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n340), .A2(new_n341), .B1(new_n342), .B2(new_n307), .ZN(new_n343));
  INV_X1    g157(.A(new_n334), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n335), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G122), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT8), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n196), .A2(G146), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT65), .B1(new_n223), .B2(G143), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT65), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n196), .A3(G146), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n349), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G128), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n223), .A2(G143), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n196), .A2(G146), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n208), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT0), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(new_n265), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n358), .A2(new_n359), .B1(KEYINPUT0), .B2(G128), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT64), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n364), .A3(new_n265), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n353), .A2(new_n365), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n257), .A2(G224), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT88), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT89), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n363), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(KEYINPUT7), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n378), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n363), .A2(new_n372), .A3(new_n380), .A4(new_n376), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n346), .A2(new_n348), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n332), .A2(KEYINPUT4), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  OR2_X1    g198(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n385), .A2(new_n386), .B1(G104), .B2(new_n274), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n218), .A2(G107), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n327), .B1(new_n326), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G101), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n329), .B1(new_n331), .B2(new_n327), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT82), .B1(new_n393), .B2(G101), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n384), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  OAI22_X1  g209(.A1(new_n322), .A2(new_n324), .B1(new_n321), .B2(new_n323), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n397), .A3(G101), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n340), .A2(new_n341), .ZN(new_n401));
  AND4_X1   g215(.A1(new_n400), .A2(new_n401), .A3(new_n344), .A4(new_n314), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n343), .B2(new_n344), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n399), .B(new_n347), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n382), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n189), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT90), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n408));
  INV_X1    g222(.A(new_n347), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(KEYINPUT6), .A3(new_n404), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n363), .A2(new_n372), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(new_n374), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(new_n414), .A3(new_n409), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT90), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n405), .A2(new_n417), .A3(new_n189), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n407), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT91), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n405), .B2(new_n189), .ZN(new_n421));
  AOI211_X1 g235(.A(KEYINPUT90), .B(G902), .C1(new_n382), .C2(new_n404), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT91), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n416), .ZN(new_n425));
  OAI21_X1  g239(.A(G210), .B1(G237), .B2(G902), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(KEYINPUT92), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n420), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n423), .A2(new_n426), .A3(new_n416), .ZN(new_n429));
  AOI211_X1 g243(.A(new_n188), .B(new_n302), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT11), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n267), .B2(G137), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n267), .A2(G137), .ZN(new_n433));
  INV_X1    g247(.A(G137), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(KEYINPUT11), .A3(G134), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G131), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT66), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n432), .A2(new_n435), .A3(new_n198), .A4(new_n433), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n436), .A2(KEYINPUT66), .A3(G131), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n371), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n267), .A2(G137), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n434), .A2(G134), .ZN(new_n444));
  OAI21_X1  g258(.A(G131), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n362), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT30), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n442), .A2(new_n447), .A3(KEYINPUT30), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n396), .A3(new_n451), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n340), .A2(new_n341), .B1(new_n339), .B2(new_n313), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n442), .A3(new_n447), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT70), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT70), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n453), .A2(new_n456), .A3(new_n442), .A4(new_n447), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT26), .B(G101), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n190), .A2(G210), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n452), .A2(new_n455), .A3(new_n457), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT31), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n455), .A2(new_n457), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT31), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n466), .A2(new_n467), .A3(new_n463), .A4(new_n452), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT28), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n455), .B2(new_n457), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n454), .A2(new_n469), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n448), .A2(new_n396), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n462), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n468), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(G472), .A2(G902), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT72), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT32), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT72), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n475), .A2(new_n480), .A3(new_n476), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(KEYINPUT32), .A3(new_n476), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT73), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n448), .A2(new_n484), .A3(new_n396), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n448), .B2(new_n396), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n455), .B(new_n457), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT28), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n463), .A2(KEYINPUT29), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n471), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT74), .ZN(new_n491));
  INV_X1    g305(.A(new_n471), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(new_n487), .B2(KEYINPUT28), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT74), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n489), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n452), .A2(new_n455), .A3(new_n457), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT29), .B1(new_n496), .B2(new_n462), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n471), .A2(new_n472), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n463), .B(new_n498), .C1(new_n466), .C2(new_n469), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n491), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n501), .A2(KEYINPUT75), .A3(G472), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT75), .B1(new_n501), .B2(G472), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n482), .B(new_n483), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n265), .A2(G119), .ZN(new_n505));
  INV_X1    g319(.A(G119), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G128), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT24), .B(G110), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT23), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n506), .B2(G128), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n265), .A2(KEYINPUT23), .A3(G119), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n510), .B1(G110), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n211), .A2(new_n223), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n515), .B1(new_n516), .B2(new_n239), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n238), .A2(new_n224), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n508), .A2(new_n509), .ZN(new_n519));
  INV_X1    g333(.A(G110), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n512), .A2(new_n513), .A3(new_n520), .A4(new_n507), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT77), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  AND4_X1   g337(.A1(KEYINPUT77), .A2(new_n522), .A3(new_n224), .A4(new_n238), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n517), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT78), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT22), .B(G137), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT79), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n529), .B(new_n530), .Z(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT78), .B(new_n517), .C1(new_n523), .C2(new_n524), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT80), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n527), .A2(KEYINPUT80), .A3(new_n532), .A4(new_n533), .ZN(new_n537));
  INV_X1    g351(.A(new_n525), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n531), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n536), .A2(new_n189), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT25), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n534), .A2(new_n535), .B1(new_n531), .B2(new_n538), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n189), .A4(new_n537), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n289), .B1(G234), .B2(new_n189), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n542), .A2(new_n537), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n545), .A2(G902), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G469), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G140), .ZN(new_n553));
  INV_X1    g367(.A(G227), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(G953), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n553), .B(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n440), .A2(new_n441), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n344), .A2(KEYINPUT10), .A3(new_n362), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n390), .A2(new_n391), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n393), .A2(KEYINPUT82), .A3(G101), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n383), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n398), .A2(new_n371), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n355), .A2(KEYINPUT83), .ZN(new_n566));
  INV_X1    g380(.A(new_n353), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n356), .A2(KEYINPUT84), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT84), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n358), .A2(new_n569), .A3(KEYINPUT1), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(G128), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT83), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n353), .A2(new_n573), .A3(new_n354), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n566), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT10), .B1(new_n575), .B2(new_n344), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n559), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT86), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n353), .A2(new_n354), .B1(new_n357), .B2(new_n360), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n334), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n564), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n582), .B1(new_n395), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n575), .A2(new_n344), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n581), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(KEYINPUT86), .A3(new_n559), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n584), .A2(new_n558), .A3(new_n586), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n557), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n334), .A2(new_n580), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n558), .B1(new_n585), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT12), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT85), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n594), .B1(new_n558), .B2(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n593), .A2(new_n596), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n590), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n599), .A2(new_n600), .A3(new_n556), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n552), .B(new_n189), .C1(new_n591), .C2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n600), .A2(new_n556), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n589), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n590), .B1(new_n597), .B2(new_n598), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n556), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n606), .A3(G469), .ZN(new_n607));
  NAND2_X1  g421(.A1(G469), .A2(G902), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n602), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G221), .B1(new_n290), .B2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n430), .A2(new_n504), .A3(new_n551), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  INV_X1    g428(.A(new_n262), .ZN(new_n615));
  AND4_X1   g429(.A1(new_n426), .A2(new_n407), .A3(new_n416), .A4(new_n418), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n426), .B1(new_n423), .B2(new_n416), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n187), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n288), .A2(KEYINPUT97), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT33), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n295), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n293), .A2(new_n619), .A3(KEYINPUT33), .A4(new_n294), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n621), .A2(G478), .A3(new_n189), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n296), .A2(new_n299), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n256), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n481), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n480), .B1(new_n475), .B2(new_n476), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n475), .A2(new_n189), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(G472), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n630), .A2(new_n609), .A3(new_n610), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n627), .A2(new_n633), .A3(new_n551), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  XNOR2_X1  g450(.A(new_n252), .B(KEYINPUT20), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n301), .A3(new_n233), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n618), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n633), .A3(new_n551), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  AOI21_X1  g456(.A(new_n188), .B1(new_n428), .B2(new_n429), .ZN(new_n643));
  INV_X1    g457(.A(new_n302), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n527), .A2(new_n533), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT36), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n531), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n527), .B(new_n533), .C1(KEYINPUT36), .C2(new_n532), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n647), .A2(new_n548), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n546), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n633), .A2(new_n643), .A3(new_n644), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  OAI211_X1 g468(.A(new_n651), .B(new_n187), .C1(new_n616), .C2(new_n617), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n501), .A2(G472), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT75), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n501), .A2(KEYINPUT75), .A3(G472), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n482), .A2(new_n483), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n655), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n259), .B1(new_n260), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n638), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n665), .A2(new_n609), .A3(new_n610), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XOR2_X1   g482(.A(new_n664), .B(KEYINPUT39), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n612), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT99), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n428), .A2(new_n429), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT38), .Z(new_n675));
  AND3_X1   g489(.A1(new_n487), .A2(KEYINPUT98), .A3(new_n462), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT98), .B1(new_n487), .B2(new_n462), .ZN(new_n677));
  INV_X1    g491(.A(new_n464), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n679), .B2(G902), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n661), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n545), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n540), .B2(KEYINPUT25), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n649), .B1(new_n684), .B2(new_n544), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n256), .A2(new_n301), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n187), .A3(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n675), .A2(new_n682), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n673), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  INV_X1    g504(.A(new_n664), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n256), .A2(new_n625), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT100), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n256), .A2(new_n625), .A3(new_n694), .A4(new_n691), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n611), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n662), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  AOI21_X1  g513(.A(KEYINPUT86), .B1(new_n587), .B2(new_n559), .ZN(new_n700));
  AOI211_X1 g514(.A(new_n578), .B(new_n558), .C1(new_n584), .C2(new_n586), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n590), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n599), .ZN(new_n703));
  AOI22_X1  g517(.A1(new_n702), .A2(new_n556), .B1(new_n703), .B2(new_n603), .ZN(new_n704));
  OAI21_X1  g518(.A(G469), .B1(new_n704), .B2(G902), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n610), .A3(new_n602), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n504), .A2(new_n627), .A3(new_n551), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT41), .B(G113), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT101), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n708), .B(new_n710), .ZN(G15));
  NAND4_X1  g525(.A1(new_n504), .A2(new_n639), .A3(new_n551), .A4(new_n707), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT102), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NOR2_X1   g528(.A1(new_n706), .A2(new_n302), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT103), .B1(new_n662), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n655), .ZN(new_n717));
  AND4_X1   g531(.A1(KEYINPUT103), .A2(new_n504), .A3(new_n717), .A4(new_n715), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n506), .ZN(G21));
  AND4_X1   g534(.A1(new_n615), .A2(new_n705), .A3(new_n610), .A4(new_n602), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n465), .B(new_n468), .C1(new_n493), .C2(new_n463), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n476), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n546), .A2(new_n632), .A3(new_n723), .A4(new_n549), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n426), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n419), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n188), .B1(new_n727), .B2(new_n429), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n721), .A2(new_n725), .A3(new_n728), .A4(new_n686), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n187), .B(new_n686), .C1(new_n616), .C2(new_n617), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n705), .A2(new_n615), .A3(new_n610), .A4(new_n602), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(KEYINPUT104), .A3(new_n725), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  AND2_X1   g551(.A1(new_n707), .A2(new_n728), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n632), .A2(new_n723), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT105), .B1(new_n739), .B2(new_n685), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n631), .A2(G472), .B1(new_n722), .B2(new_n476), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n651), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n696), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  AOI21_X1  g560(.A(new_n550), .B1(new_n660), .B2(new_n661), .ZN(new_n747));
  INV_X1    g561(.A(new_n696), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n428), .A2(new_n187), .A3(new_n429), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n607), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n604), .A2(new_n606), .A3(KEYINPUT106), .A4(G469), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n602), .A3(new_n608), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n610), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n747), .A2(new_n748), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n749), .A2(new_n754), .A3(new_n696), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n477), .B(KEYINPUT32), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n550), .B1(new_n660), .B2(new_n759), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n756), .A2(new_n757), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT107), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n198), .ZN(G33));
  NAND3_X1  g577(.A1(new_n747), .A2(new_n665), .A3(new_n755), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  INV_X1    g579(.A(new_n625), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n256), .ZN(new_n767));
  NOR2_X1   g581(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n768));
  NAND2_X1  g582(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n767), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n767), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n630), .A2(new_n632), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n651), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT110), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n604), .A2(new_n606), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n552), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n779), .B2(new_n778), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n608), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n602), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(KEYINPUT108), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n602), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT108), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n781), .A2(new_n608), .ZN(new_n787));
  OAI22_X1  g601(.A1(new_n785), .A2(new_n786), .B1(KEYINPUT46), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n610), .B(new_n669), .C1(new_n784), .C2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n749), .B1(new_n774), .B2(new_n775), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n777), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  OAI21_X1  g607(.A(new_n610), .B1(new_n784), .B2(new_n788), .ZN(new_n794));
  XOR2_X1   g608(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT47), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(KEYINPUT111), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n610), .B(new_n799), .C1(new_n784), .C2(new_n788), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n504), .A2(new_n749), .A3(new_n551), .A4(new_n696), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n796), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  AND4_X1   g617(.A1(new_n551), .A2(new_n767), .A3(new_n187), .A4(new_n610), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n705), .A2(new_n602), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT49), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n675), .A2(new_n682), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n772), .A2(new_n259), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n749), .A2(new_n706), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n760), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT48), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n551), .A2(new_n682), .A3(new_n259), .A4(new_n809), .ZN(new_n814));
  INV_X1    g628(.A(new_n626), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n808), .A2(new_n725), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n258), .B1(new_n818), .B2(new_n738), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n813), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n817), .A2(new_n187), .A3(new_n706), .ZN(new_n821));
  NOR2_X1   g635(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n675), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n740), .A2(new_n743), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n811), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n821), .A2(new_n675), .ZN(new_n827));
  XOR2_X1   g641(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n828));
  AOI21_X1  g642(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n814), .A2(new_n233), .A3(new_n637), .A4(new_n766), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n829), .A2(KEYINPUT51), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n610), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n805), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n796), .ZN(new_n834));
  INV_X1    g648(.A(new_n800), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n817), .A2(new_n749), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n820), .B1(new_n831), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n833), .B(KEYINPUT113), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n834), .B2(new_n835), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n837), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n829), .A2(new_n842), .A3(new_n830), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n844), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n839), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT104), .B1(new_n734), .B2(new_n725), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n732), .A2(new_n733), .A3(new_n724), .A4(new_n730), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n708), .B(new_n712), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n638), .A2(new_n626), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n262), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n633), .A2(new_n643), .A3(new_n854), .A4(new_n551), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n504), .A2(new_n551), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n643), .A2(new_n612), .A3(new_n644), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n652), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n719), .A2(new_n851), .A3(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n504), .B(new_n717), .C1(new_n697), .C2(new_n666), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n732), .A2(new_n651), .A3(new_n664), .ZN(new_n861));
  INV_X1    g675(.A(new_n754), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n681), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n860), .A2(new_n863), .A3(new_n745), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n860), .A2(new_n863), .A3(new_n745), .A4(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n256), .A2(new_n301), .A3(new_n664), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n610), .A2(new_n609), .A3(new_n651), .A4(new_n869), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n744), .A2(new_n862), .B1(new_n504), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n764), .B1(new_n871), .B2(new_n749), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n761), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n859), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n613), .A2(KEYINPUT53), .A3(new_n652), .A4(new_n855), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n761), .A2(new_n872), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT112), .ZN(new_n879));
  INV_X1    g693(.A(new_n851), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n504), .A2(new_n717), .A3(new_n715), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT103), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n881), .B(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n879), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n719), .A2(new_n851), .A3(KEYINPUT112), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n878), .B(new_n868), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n876), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n874), .B(KEYINPUT53), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(new_n887), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n848), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(G952), .A2(G953), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n807), .B1(new_n891), .B2(new_n892), .ZN(G75));
  NOR2_X1   g707(.A1(new_n257), .A2(G952), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n189), .B1(new_n876), .B2(new_n886), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(G210), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n411), .A2(new_n415), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n413), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n895), .A2(new_n427), .ZN(new_n901));
  XNOR2_X1  g715(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n894), .B(new_n900), .C1(new_n901), .C2(new_n903), .ZN(G51));
  NAND2_X1  g718(.A1(new_n876), .A2(new_n886), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(KEYINPUT117), .A3(new_n888), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT54), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n608), .B(KEYINPUT57), .Z(new_n910));
  NAND3_X1  g724(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT118), .ZN(new_n912));
  INV_X1    g726(.A(new_n704), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n907), .A2(new_n914), .A3(new_n909), .A4(new_n910), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n895), .B(new_n780), .C1(new_n779), .C2(new_n778), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n894), .B1(new_n916), .B2(new_n917), .ZN(G54));
  NAND2_X1  g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT119), .Z(new_n920));
  NAND3_X1  g734(.A1(new_n895), .A2(new_n250), .A3(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n921), .A2(KEYINPUT120), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(KEYINPUT120), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n250), .B1(new_n895), .B2(new_n920), .ZN(new_n924));
  NOR4_X1   g738(.A1(new_n922), .A2(new_n923), .A3(new_n894), .A4(new_n924), .ZN(G60));
  INV_X1    g739(.A(new_n894), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n299), .A2(new_n189), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n890), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n621), .A2(new_n622), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND4_X1   g746(.A1(new_n931), .A2(new_n907), .A3(new_n909), .A4(new_n929), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(G63));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT60), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n876), .B2(new_n886), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n647), .A2(new_n648), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n894), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n935), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n938), .A2(new_n547), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n940), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n942), .B(new_n944), .Z(G66));
  INV_X1    g759(.A(new_n859), .ZN(new_n946));
  NAND2_X1  g760(.A1(G224), .A2(G953), .ZN(new_n947));
  OAI22_X1  g761(.A1(new_n946), .A2(G953), .B1(new_n261), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n897), .B1(G898), .B2(new_n257), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n948), .B(new_n949), .Z(G69));
  OAI21_X1  g764(.A(G953), .B1(new_n554), .B2(new_n663), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT124), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n954));
  NOR4_X1   g768(.A1(new_n671), .A2(new_n856), .A3(new_n749), .A4(new_n853), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n956), .A2(new_n792), .A3(new_n802), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n860), .A2(new_n745), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n689), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n689), .A2(KEYINPUT62), .A3(new_n960), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n958), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n450), .A2(new_n451), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(new_n244), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n967), .A2(G953), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n954), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n760), .A2(new_n728), .A3(new_n686), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n802), .B1(new_n789), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n792), .A2(new_n960), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n792), .A2(KEYINPUT125), .A3(new_n960), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n764), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n761), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT126), .Z(new_n983));
  AOI21_X1  g797(.A(G953), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n967), .B1(G900), .B2(new_n257), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n971), .B(new_n973), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n984), .A2(new_n985), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n972), .B1(new_n987), .B2(new_n970), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n986), .A2(new_n988), .ZN(G72));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  INV_X1    g805(.A(new_n965), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(new_n946), .ZN(new_n993));
  INV_X1    g807(.A(new_n496), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n994), .A2(new_n462), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n980), .A2(new_n859), .A3(new_n983), .ZN(new_n997));
  AOI211_X1 g811(.A(new_n463), .B(new_n496), .C1(new_n997), .C2(new_n991), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n994), .A2(new_n463), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n991), .B1(new_n999), .B2(new_n678), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n926), .B1(new_n889), .B2(new_n1000), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n996), .A2(new_n998), .A3(new_n1001), .ZN(G57));
endmodule


