//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n194));
  OR3_X1    g008(.A1(new_n192), .A2(KEYINPUT16), .A3(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT73), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n195), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT73), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n194), .A2(new_n195), .A3(new_n201), .A4(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  OR2_X1    g017(.A1(KEYINPUT68), .A2(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT68), .A2(G128), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n204), .A2(G119), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G119), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT24), .B(G110), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G110), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT23), .B1(new_n207), .B2(G119), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(new_n208), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .A4(new_n205), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n203), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n209), .B1(new_n206), .B2(new_n208), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n213), .A2(new_n214), .A3(new_n211), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n196), .A2(KEYINPUT74), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT74), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n194), .A2(new_n195), .A3(new_n222), .A4(G146), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n191), .A2(new_n193), .A3(new_n199), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n220), .A2(new_n221), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G953), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(G221), .A3(G234), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n228), .B(KEYINPUT75), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT22), .B(G137), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n217), .A2(new_n225), .A3(new_n231), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT25), .B1(new_n235), .B2(new_n188), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n217), .A2(new_n225), .A3(new_n231), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n231), .B1(new_n217), .B2(new_n225), .ZN(new_n238));
  OAI211_X1 g052(.A(KEYINPUT25), .B(new_n188), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n189), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT76), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n188), .B1(new_n237), .B2(new_n238), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n239), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT76), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n189), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n189), .A2(G902), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n235), .A2(KEYINPUT77), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n235), .A2(KEYINPUT77), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n242), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(G472), .A2(G902), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT11), .A3(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n259), .A3(new_n263), .A4(new_n260), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(KEYINPUT67), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n261), .A2(new_n266), .A3(G131), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT66), .A2(G143), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(G146), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n199), .A2(G143), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n272), .A2(KEYINPUT0), .A3(G128), .A4(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT0), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(new_n207), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n277), .A2(new_n278), .B1(KEYINPUT0), .B2(G128), .ZN(new_n279));
  AOI21_X1  g093(.A(G146), .B1(new_n270), .B2(new_n271), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n199), .A2(G143), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n265), .A2(new_n267), .A3(new_n274), .A4(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n284));
  INV_X1    g098(.A(G116), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(G119), .ZN(new_n286));
  INV_X1    g100(.A(G119), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(G116), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G113), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT2), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G113), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n287), .A2(G116), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n285), .A2(G119), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT69), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n289), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(G116), .B(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n260), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n256), .A2(G137), .ZN(new_n305));
  OAI21_X1  g119(.A(G131), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(KEYINPUT66), .A2(G143), .ZN(new_n307));
  NOR2_X1   g121(.A1(KEYINPUT66), .A2(G143), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n199), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n281), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n204), .A2(new_n205), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n273), .A2(KEYINPUT1), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n272), .A2(new_n273), .A3(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n264), .B(new_n306), .C1(new_n313), .C2(new_n315), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n283), .A2(new_n303), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT26), .B(G101), .ZN(new_n318));
  INV_X1    g132(.A(G237), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n227), .A3(G210), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n318), .B(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT71), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n283), .A2(new_n303), .A3(new_n316), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT71), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n323), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n283), .A2(new_n316), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT64), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT30), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n333));
  AOI211_X1 g147(.A(KEYINPUT64), .B(new_n333), .C1(new_n283), .C2(new_n316), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n302), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT31), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n329), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n303), .B1(new_n283), .B2(new_n316), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT28), .B1(new_n317), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT28), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n326), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n324), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n336), .B1(new_n329), .B2(new_n335), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n254), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT32), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT32), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n348), .B(new_n254), .C1(new_n344), .C2(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n339), .A2(KEYINPUT29), .A3(new_n323), .A4(new_n341), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n188), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT72), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(KEYINPUT72), .A3(new_n188), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n323), .B1(new_n335), .B2(new_n326), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n357), .B1(new_n342), .B2(new_n324), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n354), .B(new_n355), .C1(new_n356), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G472), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n253), .B1(new_n350), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G475), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n319), .A2(new_n227), .A3(G143), .A4(G214), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT66), .B(G143), .ZN(new_n364));
  INV_X1    g178(.A(G214), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n365), .A2(G237), .A3(G953), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n363), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(G131), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT17), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT87), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(new_n367), .B2(G131), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n319), .A2(new_n227), .A3(G214), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n270), .A3(new_n271), .ZN(new_n374));
  AOI211_X1 g188(.A(KEYINPUT87), .B(new_n263), .C1(new_n374), .C2(new_n363), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n369), .B(new_n370), .C1(new_n372), .C2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n203), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n367), .A2(G131), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT87), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n367), .A2(new_n371), .A3(G131), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(KEYINPUT17), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n376), .A2(new_n377), .A3(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n192), .A2(G140), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n190), .A2(G125), .ZN(new_n384));
  OAI21_X1  g198(.A(G146), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n224), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT18), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(new_n263), .ZN(new_n388));
  OAI221_X1 g202(.A(new_n386), .B1(new_n367), .B2(new_n388), .C1(new_n378), .C2(new_n387), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G113), .B(G122), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n382), .A2(new_n393), .A3(new_n389), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n362), .B1(new_n397), .B2(new_n188), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT89), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n378), .A2(new_n387), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n386), .B1(new_n367), .B2(new_n388), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n221), .A2(new_n223), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT19), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n383), .B2(new_n384), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT19), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n199), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT88), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(KEYINPUT88), .A3(new_n199), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n404), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n369), .B1(new_n372), .B2(new_n375), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n403), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n400), .B1(new_n415), .B2(new_n393), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT88), .B1(new_n408), .B2(new_n199), .ZN(new_n417));
  AOI211_X1 g231(.A(new_n410), .B(G146), .C1(new_n406), .C2(new_n407), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n221), .B(new_n223), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n368), .B1(new_n379), .B2(new_n380), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n389), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT89), .A3(new_n394), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n416), .A2(new_n396), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n424));
  NOR2_X1   g238(.A1(G475), .A2(G902), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(new_n423), .B2(new_n425), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n399), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT90), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n399), .B(new_n431), .C1(new_n426), .C2(new_n428), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n307), .A2(new_n308), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G128), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n204), .A2(G143), .A3(new_n205), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n437), .A2(new_n256), .ZN(new_n438));
  XNOR2_X1  g252(.A(G116), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT91), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n440), .A2(G107), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(G107), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n438), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT13), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n435), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n434), .A2(KEYINPUT13), .A3(G128), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(new_n436), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n447), .A2(new_n448), .A3(G134), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n447), .B2(G134), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n443), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n285), .A2(KEYINPUT14), .A3(G122), .ZN(new_n452));
  INV_X1    g266(.A(new_n439), .ZN(new_n453));
  OAI211_X1 g267(.A(G107), .B(new_n452), .C1(new_n453), .C2(KEYINPUT14), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n437), .A2(new_n256), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n441), .B(new_n454), .C1(new_n438), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT9), .B(G234), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n458), .A2(new_n187), .A3(G953), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n451), .A2(new_n456), .A3(new_n459), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G478), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n463), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(G234), .A2(G237), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n467), .A2(G952), .A3(new_n227), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n467), .A2(G902), .A3(G953), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(G898), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G469), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n265), .A2(new_n267), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n478));
  INV_X1    g292(.A(G107), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n479), .A3(G104), .ZN(new_n480));
  INV_X1    g294(.A(G101), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n392), .A2(G107), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n477), .A2(new_n480), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n392), .A2(G107), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n479), .A2(G104), .ZN(new_n485));
  OAI21_X1  g299(.A(G101), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT1), .ZN(new_n488));
  OAI21_X1  g302(.A(G128), .B1(new_n280), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n272), .A2(new_n273), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n272), .A2(new_n273), .A3(new_n314), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n483), .A2(new_n486), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n494), .A2(new_n313), .A3(new_n315), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n476), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT12), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT10), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n315), .B1(new_n490), .B2(new_n489), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n498), .B1(new_n499), .B2(new_n487), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n494), .B(KEYINPUT10), .C1(new_n315), .C2(new_n313), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G101), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(KEYINPUT4), .A3(new_n483), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT4), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n505), .A3(G101), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n504), .A2(new_n274), .A3(new_n282), .A4(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n500), .A2(new_n475), .A3(new_n501), .A4(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G110), .B(G140), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n227), .A2(G227), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n476), .B(new_n513), .C1(new_n493), .C2(new_n495), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n497), .A2(new_n508), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT78), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n501), .B(new_n507), .C1(new_n493), .C2(KEYINPUT10), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n476), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n508), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n511), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n515), .A2(new_n516), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n474), .B(new_n188), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n497), .A2(new_n508), .A3(new_n514), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n511), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n512), .A3(new_n508), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(G469), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n474), .A2(new_n188), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G221), .B1(new_n458), .B2(G902), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n433), .A2(new_n473), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT85), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT84), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT83), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n227), .A2(G224), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT7), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT82), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n281), .B1(new_n364), .B2(new_n199), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n204), .A2(new_n205), .B1(new_n273), .B2(KEYINPUT1), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n492), .B(new_n192), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT80), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n311), .A2(new_n312), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n280), .B2(new_n281), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT80), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n548), .A2(new_n549), .A3(new_n192), .A4(new_n492), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n542), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n192), .B1(new_n282), .B2(new_n274), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n546), .A2(new_n542), .A3(new_n550), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n541), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n502), .A2(G101), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n505), .A2(new_n557), .B1(new_n299), .B2(new_n301), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n504), .ZN(new_n559));
  INV_X1    g373(.A(new_n301), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT69), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT69), .B1(new_n296), .B2(new_n297), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT5), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G113), .B1(new_n296), .B2(KEYINPUT5), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n560), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n494), .ZN(new_n567));
  INV_X1    g381(.A(G122), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G110), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n211), .A2(G122), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n559), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n546), .A2(new_n550), .ZN(new_n574));
  INV_X1    g388(.A(new_n552), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n541), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT5), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n289), .B2(new_n298), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n301), .B(new_n487), .C1(new_n578), .C2(new_n564), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT8), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT8), .B1(new_n569), .B2(new_n570), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT5), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n301), .B1(new_n583), .B2(new_n564), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n582), .B1(new_n494), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT81), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n579), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n586), .B1(new_n579), .B2(new_n585), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n573), .B(new_n576), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n538), .B(new_n188), .C1(new_n556), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n574), .A2(new_n575), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(new_n539), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n559), .A2(new_n567), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n571), .B(KEYINPUT79), .Z(new_n595));
  AOI22_X1  g409(.A1(new_n573), .A2(KEYINPUT6), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n594), .A2(KEYINPUT6), .A3(new_n595), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n593), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n579), .A2(new_n585), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT81), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n558), .A2(new_n504), .B1(new_n566), .B2(new_n494), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n601), .A2(new_n587), .B1(new_n602), .B2(new_n572), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n554), .A2(new_n551), .A3(new_n552), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n603), .B(new_n576), .C1(new_n604), .C2(new_n541), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n538), .B1(new_n605), .B2(new_n188), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n537), .B1(new_n599), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G210), .B1(G237), .B2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n188), .B1(new_n556), .B2(new_n590), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT83), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n611), .A2(KEYINPUT84), .A3(new_n598), .A4(new_n591), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n607), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n611), .A2(new_n608), .A3(new_n598), .A4(new_n591), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(G214), .B1(G237), .B2(G902), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n536), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n616), .ZN(new_n618));
  AOI211_X1 g432(.A(KEYINPUT85), .B(new_n618), .C1(new_n613), .C2(new_n614), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n361), .B(new_n535), .C1(new_n617), .C2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G101), .ZN(G3));
  NOR2_X1   g435(.A1(new_n464), .A2(new_n188), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n463), .B2(new_n464), .ZN(new_n623));
  INV_X1    g437(.A(new_n462), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n459), .B1(new_n451), .B2(new_n456), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT33), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n461), .A2(new_n627), .A3(new_n462), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(G478), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n422), .A2(new_n396), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT89), .B1(new_n421), .B2(new_n394), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n425), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n427), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n431), .B1(new_n638), .B2(new_n399), .ZN(new_n639));
  AOI211_X1 g453(.A(KEYINPUT90), .B(new_n398), .C1(new_n636), .C2(new_n637), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n631), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT93), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT93), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n433), .A2(new_n643), .A3(new_n631), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n609), .B1(new_n599), .B2(new_n606), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n618), .B1(new_n646), .B2(new_n614), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n471), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n188), .B1(new_n344), .B2(new_n345), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(G472), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n346), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n652), .A2(new_n534), .A3(new_n253), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n645), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  INV_X1    g470(.A(new_n465), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n463), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n463), .A2(new_n657), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n634), .A2(new_n635), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n660), .B(new_n399), .C1(new_n428), .C2(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n662), .A2(new_n648), .A3(new_n471), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n653), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NOR2_X1   g480(.A1(new_n231), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n226), .B(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT94), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n668), .A2(new_n669), .A3(new_n249), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n669), .B1(new_n668), .B2(new_n249), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n242), .A2(new_n248), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT95), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT95), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n242), .A2(new_n675), .A3(new_n248), .A4(new_n672), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n652), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n535), .B(new_n677), .C1(new_n617), .C2(new_n619), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  AOI22_X1  g494(.A1(new_n350), .A2(new_n360), .B1(new_n674), .B2(new_n676), .ZN(new_n681));
  INV_X1    g495(.A(new_n533), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n524), .B2(new_n531), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n469), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n468), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n399), .B(new_n687), .C1(new_n661), .C2(new_n428), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n466), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n681), .A2(new_n683), .A3(new_n647), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XNOR2_X1  g505(.A(new_n687), .B(KEYINPUT39), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT97), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT40), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n615), .B(KEYINPUT38), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n674), .A2(new_n676), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n618), .B1(new_n658), .B2(new_n659), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n433), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n330), .A2(new_n331), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n333), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT30), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n303), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n326), .A2(new_n327), .A3(new_n323), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n327), .B1(new_n326), .B2(new_n323), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n338), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n323), .B1(new_n709), .B2(new_n326), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n188), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G472), .ZN(new_n712));
  INV_X1    g526(.A(new_n349), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT31), .B1(new_n704), .B2(new_n707), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n343), .A3(new_n337), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n348), .B1(new_n715), .B2(new_n254), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n712), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT96), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT96), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n350), .A2(new_n719), .A3(new_n712), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n695), .A2(new_n700), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n364), .ZN(G45));
  INV_X1    g537(.A(new_n687), .ZN(new_n724));
  AOI211_X1 g538(.A(new_n724), .B(new_n630), .C1(new_n430), .C2(new_n432), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n681), .A2(new_n725), .A3(new_n683), .A4(new_n647), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  OAI21_X1  g541(.A(new_n360), .B1(new_n713), .B2(new_n716), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n188), .B1(new_n522), .B2(new_n523), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G469), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n533), .A3(new_n524), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT98), .ZN(new_n732));
  INV_X1    g546(.A(new_n253), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT98), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n730), .A2(new_n734), .A3(new_n533), .A4(new_n524), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n728), .A2(new_n732), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n645), .A2(new_n736), .A3(new_n649), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT41), .B(G113), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G15));
  NAND2_X1  g553(.A1(new_n736), .A2(new_n663), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G116), .ZN(G18));
  INV_X1    g555(.A(KEYINPUT99), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n639), .A2(new_n640), .ZN(new_n743));
  INV_X1    g557(.A(new_n473), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n730), .A2(new_n533), .A3(new_n524), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n743), .A2(new_n744), .A3(new_n647), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n697), .A2(new_n728), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n742), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n648), .A2(new_n731), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n433), .A2(new_n473), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n681), .A2(new_n749), .A3(new_n750), .A4(KEYINPUT99), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  AND2_X1   g567(.A1(new_n732), .A2(new_n735), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n646), .A2(new_n614), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(new_n698), .C1(new_n639), .C2(new_n640), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n471), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT101), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n650), .A2(G472), .B1(new_n715), .B2(new_n254), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n247), .B1(new_n246), .B2(new_n189), .ZN(new_n760));
  INV_X1    g574(.A(new_n189), .ZN(new_n761));
  AOI211_X1 g575(.A(KEYINPUT76), .B(new_n761), .C1(new_n245), .C2(new_n239), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT100), .B1(new_n763), .B2(new_n252), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n242), .A2(KEYINPUT100), .A3(new_n248), .A4(new_n252), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n758), .B(new_n759), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT100), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n253), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n765), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n758), .B1(new_n771), .B2(new_n759), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n754), .B(new_n757), .C1(new_n768), .C2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  NAND3_X1  g588(.A1(new_n725), .A2(new_n749), .A3(new_n677), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G125), .ZN(G27));
  AND2_X1   g590(.A1(new_n614), .A2(new_n616), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n613), .A2(new_n777), .A3(new_n683), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n725), .A2(new_n361), .A3(new_n778), .A4(KEYINPUT102), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n613), .A2(new_n777), .A3(new_n683), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n347), .A2(new_n349), .B1(G472), .B2(new_n359), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n782), .A2(new_n783), .A3(new_n253), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT102), .B1(new_n784), .B2(new_n725), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT104), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n350), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n347), .A2(KEYINPUT104), .A3(new_n349), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n360), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n771), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n725), .A2(KEYINPUT42), .A3(new_n778), .ZN(new_n791));
  OAI22_X1  g605(.A1(new_n781), .A2(new_n785), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G131), .ZN(G33));
  NAND3_X1  g607(.A1(new_n361), .A2(new_n778), .A3(new_n689), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  INV_X1    g609(.A(KEYINPUT107), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n526), .A2(KEYINPUT45), .A3(new_n527), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT105), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT45), .B1(new_n526), .B2(new_n527), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n474), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n529), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(KEYINPUT106), .A3(KEYINPUT46), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n524), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT106), .B1(new_n801), .B2(KEYINPUT46), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n796), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n801), .A2(KEYINPUT46), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n801), .A2(KEYINPUT46), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT106), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(KEYINPUT107), .A3(new_n524), .A4(new_n802), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n805), .A2(new_n806), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(new_n533), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n692), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT108), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n743), .A2(new_n631), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT43), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n433), .A2(KEYINPUT43), .A3(new_n630), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n652), .A4(new_n697), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT44), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT109), .Z(new_n821));
  AND2_X1   g635(.A1(new_n613), .A2(new_n777), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n818), .B2(new_n819), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n814), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G137), .ZN(G39));
  INV_X1    g640(.A(KEYINPUT47), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(KEYINPUT110), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n811), .A2(new_n533), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n811), .B2(new_n533), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n783), .A2(new_n725), .A3(new_n253), .A4(new_n822), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G140), .ZN(G42));
  NAND2_X1  g650(.A1(new_n730), .A2(new_n524), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(KEYINPUT49), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n837), .A2(KEYINPUT49), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n815), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n721), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n764), .A2(new_n766), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n842), .A2(new_n618), .A3(new_n682), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n696), .A2(new_n840), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n811), .A2(new_n533), .A3(new_n829), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n846), .B(new_n847), .C1(new_n812), .C2(new_n831), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT114), .B1(new_n830), .B2(new_n832), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n848), .B(new_n849), .C1(new_n533), .C2(new_n837), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n816), .A2(new_n817), .A3(new_n468), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n768), .A2(new_n772), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n853), .A2(new_n822), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(KEYINPUT115), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n731), .A2(new_n616), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n696), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n852), .A3(new_n851), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT50), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n853), .A2(KEYINPUT50), .A3(new_n857), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n862), .B1(new_n860), .B2(new_n861), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n823), .A2(new_n731), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n733), .A2(new_n841), .A3(new_n865), .A4(new_n468), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n743), .A3(new_n630), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n851), .A2(new_n677), .A3(new_n865), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n863), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n855), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT115), .B1(new_n850), .B2(new_n854), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n845), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n853), .A2(new_n749), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT118), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n851), .A2(new_n865), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT48), .ZN(new_n877));
  OR4_X1    g691(.A1(KEYINPUT119), .A2(new_n876), .A3(new_n877), .A4(new_n790), .ZN(new_n878));
  XNOR2_X1  g692(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(new_n876), .B2(new_n790), .ZN(new_n880));
  INV_X1    g694(.A(G952), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n881), .B(G953), .C1(new_n866), .C2(new_n645), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n875), .A2(new_n878), .A3(new_n880), .A4(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n869), .B(KEYINPUT117), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n860), .A2(new_n861), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n884), .A2(new_n845), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n837), .A2(new_n533), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n854), .B1(new_n833), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n883), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n873), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n652), .A2(new_n534), .A3(new_n253), .A4(new_n471), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT111), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n743), .B2(new_n660), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n430), .A2(new_n893), .A3(new_n432), .A4(new_n660), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n641), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n892), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n617), .A2(new_n619), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n620), .B(new_n678), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n660), .A2(new_n688), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n681), .A2(new_n683), .A3(new_n822), .A4(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n725), .A2(new_n677), .A3(new_n778), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n902), .A3(new_n794), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n662), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n649), .B(new_n736), .C1(new_n645), .C2(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n906), .A2(new_n752), .A3(new_n773), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n904), .A2(new_n907), .A3(new_n792), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n683), .A2(new_n763), .A3(new_n672), .A4(new_n687), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n756), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n721), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(new_n726), .A3(new_n690), .A4(new_n775), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT52), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n891), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT112), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n790), .A2(new_n791), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n779), .A2(new_n780), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n784), .A2(new_n725), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT102), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n917), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n906), .A2(new_n752), .A3(new_n773), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n737), .A2(new_n773), .A3(new_n740), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n925), .A2(KEYINPUT112), .A3(new_n792), .A4(new_n752), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n690), .A2(new_n775), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n927), .A2(KEYINPUT52), .A3(new_n726), .A4(new_n911), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT52), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n912), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n899), .A2(new_n891), .A3(new_n903), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n924), .A2(new_n926), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n914), .A2(new_n915), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n922), .A2(new_n923), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n935), .A2(new_n931), .A3(KEYINPUT53), .A4(new_n904), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n915), .B1(new_n914), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT113), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n903), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n430), .A2(new_n432), .A3(new_n660), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT111), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n941), .A2(new_n641), .A3(new_n895), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n942), .B(new_n892), .C1(new_n619), .C2(new_n617), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(new_n620), .A3(new_n678), .A4(new_n943), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n944), .A2(new_n922), .A3(new_n923), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT53), .B1(new_n945), .B2(new_n931), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n908), .A2(new_n913), .A3(new_n891), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT54), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT113), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n914), .A2(new_n933), .A3(new_n915), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n890), .B1(new_n938), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(G952), .A2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n844), .B1(new_n952), .B2(new_n953), .ZN(G75));
  AOI21_X1  g768(.A(new_n188), .B1(new_n914), .B2(new_n933), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT56), .B1(new_n955), .B2(G210), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n596), .A2(new_n597), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n593), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT55), .Z(new_n959));
  XNOR2_X1  g773(.A(new_n956), .B(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n227), .A2(G952), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT120), .Z(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n960), .A2(new_n963), .ZN(G51));
  INV_X1    g778(.A(KEYINPUT121), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n950), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n914), .A2(new_n933), .A3(KEYINPUT121), .A4(new_n915), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n914), .A2(new_n933), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n966), .B(new_n967), .C1(new_n915), .C2(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n529), .B(KEYINPUT57), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n523), .B2(new_n522), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n955), .A2(new_n798), .A3(new_n800), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n961), .B1(new_n972), .B2(new_n973), .ZN(G54));
  AND3_X1   g788(.A1(new_n955), .A2(KEYINPUT58), .A3(G475), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n975), .A2(new_n423), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n423), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n961), .ZN(G60));
  XNOR2_X1  g792(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(new_n622), .Z(new_n980));
  NAND3_X1  g794(.A1(new_n938), .A2(new_n951), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n626), .A2(new_n628), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n980), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n963), .B1(new_n969), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT123), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n983), .A2(new_n986), .A3(KEYINPUT123), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G63));
  NAND2_X1  g805(.A1(G217), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT124), .Z(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT60), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n914), .B2(new_n933), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n250), .A2(new_n251), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n962), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(new_n668), .B2(new_n995), .ZN(new_n998));
  XOR2_X1   g812(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(G66));
  INV_X1    g814(.A(new_n470), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n227), .B1(new_n1001), .B2(G224), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n923), .A2(new_n899), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT126), .Z(new_n1004));
  AOI21_X1  g818(.A(new_n1002), .B1(new_n1004), .B2(new_n227), .ZN(new_n1005));
  INV_X1    g819(.A(G898), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n957), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1005), .B(new_n1007), .ZN(G69));
  AOI21_X1  g822(.A(new_n227), .B1(G227), .B2(G900), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n702), .A2(new_n703), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(new_n408), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G900), .A2(G953), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n927), .A2(new_n726), .ZN(new_n1014));
  AND4_X1   g828(.A1(new_n792), .A2(new_n835), .A3(new_n794), .A4(new_n1014), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n790), .A2(new_n756), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n814), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n825), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1012), .B(new_n1013), .C1(new_n1018), .C2(G953), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n722), .A2(new_n1014), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1020), .A2(KEYINPUT62), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT127), .Z(new_n1022));
  AND4_X1   g836(.A1(new_n361), .A2(new_n942), .A3(new_n694), .A4(new_n822), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1023), .B1(new_n1020), .B2(KEYINPUT62), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1022), .A2(new_n825), .A3(new_n835), .A4(new_n1024), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n1025), .A2(new_n227), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n1010), .B(new_n1019), .C1(new_n1026), .C2(new_n1012), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1019), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1012), .B1(new_n1025), .B2(new_n227), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1009), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1027), .A2(new_n1030), .ZN(G72));
  NAND2_X1  g845(.A1(G472), .A2(G902), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n1032), .B(KEYINPUT63), .Z(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(new_n1025), .B2(new_n1004), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n324), .B1(new_n335), .B2(new_n326), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1033), .B1(new_n1018), .B2(new_n1004), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n1037), .A2(new_n335), .A3(new_n326), .A4(new_n324), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n914), .A2(new_n936), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n708), .A2(new_n356), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1033), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n961), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  AND3_X1   g857(.A1(new_n1036), .A2(new_n1038), .A3(new_n1043), .ZN(G57));
endmodule


