//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n542, new_n543, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT64), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G101), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(G137), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT66), .B1(new_n461), .B2(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n458), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT65), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n460), .A2(new_n475), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n462), .A2(new_n472), .B1(new_n478), .B2(G2105), .ZN(G160));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n463), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI221_X1 g057(.A(new_n482), .B1(new_n481), .B2(new_n480), .C1(G112), .C2(new_n471), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n467), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n467), .A2(new_n471), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND3_X1  g064(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n490));
  NAND2_X1  g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n463), .A2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G102), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n471), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n460), .A2(KEYINPUT4), .A3(G138), .A4(new_n471), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n493), .A2(new_n495), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT68), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(G543), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(new_n506), .B1(KEYINPUT5), .B2(new_n502), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(G543), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n510), .A2(new_n516), .ZN(G166));
  AND2_X1   g092(.A1(new_n507), .A2(new_n511), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G89), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n522));
  INV_X1    g097(.A(new_n515), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G51), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n519), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  AOI22_X1  g101(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n509), .ZN(new_n528));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n512), .A2(new_n529), .B1(new_n530), .B2(new_n515), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(G171));
  AOI22_X1  g107(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n509), .ZN(new_n534));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  INV_X1    g110(.A(G43), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n512), .A2(new_n535), .B1(new_n536), .B2(new_n515), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  AND3_X1   g114(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G36), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n540), .A2(new_n543), .ZN(G188));
  INV_X1    g119(.A(G53), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT9), .B1(new_n515), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT9), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n511), .A2(new_n547), .A3(G53), .A4(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n507), .A2(G91), .A3(new_n511), .ZN(new_n550));
  XOR2_X1   g125(.A(KEYINPUT69), .B(G65), .Z(new_n551));
  AOI22_X1  g126(.A1(new_n507), .A2(new_n551), .B1(G78), .B2(G543), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n549), .B(new_n550), .C1(new_n509), .C2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n552), .A2(new_n509), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n556), .A2(KEYINPUT70), .A3(new_n550), .A4(new_n549), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(G299));
  INV_X1    g133(.A(G171), .ZN(G301));
  OR2_X1    g134(.A1(new_n510), .A2(new_n516), .ZN(G303));
  NAND2_X1  g135(.A1(new_n518), .A2(G87), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n523), .A2(G49), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G288));
  AOI22_X1  g139(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n565), .A2(new_n509), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n523), .A2(G48), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n518), .A2(G86), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(G305));
  AOI22_X1  g146(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n509), .ZN(new_n573));
  INV_X1    g148(.A(G85), .ZN(new_n574));
  INV_X1    g149(.A(G47), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n512), .A2(new_n574), .B1(new_n575), .B2(new_n515), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G290));
  NAND2_X1  g153(.A1(G301), .A2(G868), .ZN(new_n579));
  NAND2_X1  g154(.A1(G79), .A2(G543), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT72), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n503), .A2(new_n506), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G66), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT73), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n588), .B(new_n581), .C1(new_n584), .C2(new_n585), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(G651), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n523), .A2(G54), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n507), .A2(G92), .A3(new_n511), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n579), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n579), .B1(new_n595), .B2(G868), .ZN(G321));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G299), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G297));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G280));
  XNOR2_X1  g176(.A(KEYINPUT74), .B(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(G860), .B2(new_n602), .ZN(G148));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n538), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n486), .A2(G123), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT75), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n484), .A2(G135), .ZN(new_n610));
  NOR2_X1   g185(.A1(G99), .A2(G2105), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(new_n471), .B2(G111), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(G2096), .Z(new_n614));
  NAND2_X1  g189(.A1(new_n460), .A2(new_n494), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(KEYINPUT15), .B(G2435), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT77), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(G2427), .B(G2430), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2451), .B(G2454), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2443), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2446), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n627), .A2(new_n630), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n627), .A2(new_n630), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n634), .A2(G14), .A3(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT78), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g215(.A1(new_n634), .A2(KEYINPUT78), .A3(G14), .A4(new_n637), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n647), .B2(KEYINPUT18), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n645), .A2(new_n646), .ZN(new_n650));
  AOI21_X1  g225(.A(KEYINPUT18), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  MUX2_X1   g226(.A(new_n648), .B(new_n644), .S(new_n651), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT79), .B(G2096), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(G227));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  AOI22_X1  g240(.A1(new_n663), .A2(KEYINPUT20), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n659), .A3(new_n662), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n666), .B(new_n668), .C1(KEYINPUT20), .C2(new_n663), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT80), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G1991), .Z(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1986), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n671), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G229));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(G29), .B2(G32), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n484), .A2(G141), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT90), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n682));
  NAND3_X1  g257(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  AOI22_X1  g259(.A1(new_n486), .A2(G129), .B1(G105), .B2(new_n494), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g263(.A1(new_n681), .A2(KEYINPUT92), .A3(new_n684), .A4(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(new_n679), .B(new_n678), .S(new_n692), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT27), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  OAI21_X1  g271(.A(KEYINPUT23), .B1(new_n599), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(G20), .ZN(new_n698));
  MUX2_X1   g273(.A(KEYINPUT23), .B(new_n697), .S(new_n698), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G1956), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n691), .A2(G26), .ZN(new_n701));
  OR2_X1    g276(.A1(G104), .A2(G2105), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n702), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT85), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n486), .A2(G128), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n484), .A2(G140), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n701), .B1(new_n707), .B2(G29), .ZN(new_n708));
  MUX2_X1   g283(.A(new_n701), .B(new_n708), .S(KEYINPUT28), .Z(new_n709));
  XOR2_X1   g284(.A(KEYINPUT86), .B(G2067), .Z(new_n710));
  XOR2_X1   g285(.A(new_n709), .B(new_n710), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n696), .A2(G19), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n538), .B2(new_n696), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(G1341), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n691), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n691), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G2090), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G5), .A2(G16), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G171), .B2(G16), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(G1961), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n691), .A2(G27), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G164), .B2(new_n691), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G2078), .ZN(new_n725));
  NOR4_X1   g300(.A1(new_n711), .A2(new_n719), .A3(new_n722), .A4(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n699), .A2(G1956), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT24), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n691), .B1(new_n728), .B2(G34), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(KEYINPUT88), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n729), .A2(KEYINPUT88), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n730), .B(new_n731), .C1(new_n728), .C2(G34), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G160), .B2(G29), .ZN(new_n733));
  OAI22_X1  g308(.A1(new_n717), .A2(G2090), .B1(G2084), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(G2084), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT89), .Z(new_n736));
  NOR2_X1   g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AND4_X1   g312(.A1(new_n700), .A2(new_n726), .A3(new_n727), .A4(new_n737), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT87), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G2105), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n484), .A2(G139), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n494), .A2(G103), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT25), .Z(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  MUX2_X1   g320(.A(G33), .B(new_n745), .S(G29), .Z(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(G2072), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n696), .A2(G21), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G168), .B2(new_n696), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT94), .B(G1966), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT31), .B(G11), .ZN(new_n752));
  INV_X1    g327(.A(G28), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(KEYINPUT30), .B2(new_n753), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n613), .B2(new_n691), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G1961), .B2(new_n721), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n751), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT95), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT84), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G4), .B2(G16), .ZN(new_n761));
  OR3_X1    g336(.A1(new_n760), .A2(G4), .A3(G16), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n761), .B(new_n762), .C1(new_n763), .C2(new_n696), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1348), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n738), .A2(new_n747), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n577), .A2(new_n696), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n696), .B2(G24), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT82), .B(G1986), .Z(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n691), .A2(G25), .ZN(new_n772));
  OR2_X1    g347(.A1(G95), .A2(G2105), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT81), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n463), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n775), .B1(new_n774), .B2(new_n773), .C1(G107), .C2(new_n471), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n484), .A2(G131), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n486), .A2(G119), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n772), .B1(new_n780), .B2(new_n691), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT35), .B(G1991), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n770), .A2(new_n771), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n696), .A2(G23), .ZN(new_n785));
  INV_X1    g360(.A(G288), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n696), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT33), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT33), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G1976), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n788), .A2(G1976), .A3(new_n789), .ZN(new_n793));
  INV_X1    g368(.A(G1971), .ZN(new_n794));
  NOR2_X1   g369(.A1(G166), .A2(new_n696), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n696), .B2(G22), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(G6), .A2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G305), .B2(new_n696), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT32), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT83), .B(G1981), .Z(new_n801));
  AOI21_X1  g376(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n796), .A2(new_n794), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n784), .B1(new_n805), .B2(KEYINPUT34), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n781), .A2(new_n782), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT34), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n802), .A2(new_n803), .A3(new_n808), .A4(new_n804), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(KEYINPUT36), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n806), .A2(new_n812), .A3(new_n807), .A4(new_n809), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n695), .B(new_n766), .C1(new_n811), .C2(new_n813), .ZN(G311));
  AOI21_X1  g389(.A(new_n766), .B1(new_n811), .B2(new_n813), .ZN(new_n815));
  INV_X1    g390(.A(new_n695), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(G150));
  AOI22_X1  g392(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n509), .ZN(new_n819));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n512), .A2(new_n820), .B1(new_n821), .B2(new_n515), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n595), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n538), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n819), .A2(new_n822), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n534), .B2(new_n537), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT39), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n827), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n825), .B1(new_n833), .B2(G860), .ZN(G145));
  INV_X1    g409(.A(G37), .ZN(new_n835));
  INV_X1    g410(.A(new_n707), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n741), .A2(new_n837), .A3(new_n742), .A4(new_n744), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n688), .A2(new_n689), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n838), .B1(new_n688), .B2(new_n689), .ZN(new_n841));
  OAI21_X1  g416(.A(G164), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n841), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n843), .A2(new_n500), .A3(new_n839), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n836), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n486), .A2(G130), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n484), .A2(G142), .ZN(new_n848));
  NOR2_X1   g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n616), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n780), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n842), .A2(new_n844), .A3(new_n836), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n846), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n853), .B1(new_n857), .B2(new_n845), .ZN(new_n858));
  XNOR2_X1  g433(.A(G162), .B(G160), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n613), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n856), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n856), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n860), .B1(new_n858), .B2(new_n863), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n835), .B(new_n862), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g442(.A(new_n604), .B(new_n831), .Z(new_n868));
  AND2_X1   g443(.A1(new_n590), .A2(new_n591), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n869), .A2(new_n594), .B1(new_n555), .B2(new_n557), .ZN(new_n870));
  NOR2_X1   g445(.A1(G299), .A2(new_n763), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n595), .A2(new_n555), .A3(new_n557), .ZN(new_n875));
  NAND2_X1  g450(.A1(G299), .A2(new_n763), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n875), .A2(new_n877), .A3(new_n876), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n880), .B1(new_n883), .B2(new_n879), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n874), .B1(new_n884), .B2(new_n868), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n885), .A2(KEYINPUT42), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(KEYINPUT42), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(G303), .A2(new_n786), .ZN(new_n889));
  NOR2_X1   g464(.A1(G166), .A2(G288), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n569), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(new_n570), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n569), .A2(KEYINPUT71), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(G305), .B1(new_n889), .B2(new_n890), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n895), .A2(new_n896), .A3(new_n577), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n577), .B1(new_n895), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n888), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n886), .A2(new_n887), .A3(new_n899), .ZN(new_n902));
  OAI21_X1  g477(.A(G868), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(G868), .B2(new_n829), .ZN(G295));
  OAI21_X1  g479(.A(new_n903), .B1(G868), .B2(new_n829), .ZN(G331));
  XOR2_X1   g480(.A(KEYINPUT99), .B(KEYINPUT44), .Z(new_n906));
  NAND3_X1  g481(.A1(new_n828), .A2(new_n830), .A3(G301), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(G301), .B1(new_n828), .B2(new_n830), .ZN(new_n909));
  OAI21_X1  g484(.A(G286), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n831), .A2(G171), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(G168), .A3(new_n907), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n910), .A2(new_n912), .A3(KEYINPUT100), .A4(new_n872), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n912), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(new_n884), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n915), .B2(new_n873), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n916), .A2(new_n917), .A3(new_n899), .A4(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT41), .B1(new_n870), .B2(new_n871), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n879), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n880), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n915), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n925), .A2(new_n899), .A3(new_n919), .A4(new_n913), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT101), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n919), .A3(new_n913), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n900), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n920), .A2(new_n927), .A3(new_n835), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n883), .B1(new_n912), .B2(new_n910), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n915), .A2(new_n873), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n900), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n920), .A2(new_n927), .A3(new_n935), .A4(new_n835), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n906), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n936), .B2(KEYINPUT43), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n926), .B(new_n917), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n941), .A2(new_n942), .A3(new_n835), .A4(new_n929), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n940), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n940), .B2(new_n943), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n938), .B1(new_n945), .B2(new_n946), .ZN(G397));
  INV_X1    g522(.A(KEYINPUT50), .ZN(new_n948));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  INV_X1    g524(.A(new_n491), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n460), .B2(G126), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n495), .B1(new_n951), .B2(new_n471), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n498), .A2(new_n499), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n948), .B(new_n949), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT106), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n500), .A2(new_n956), .A3(new_n948), .A4(new_n949), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n948), .B1(new_n500), .B2(new_n949), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n462), .A2(new_n472), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n478), .A2(G2105), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(G40), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G2084), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n958), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1966), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(G160), .B(G40), .C1(new_n967), .C2(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n498), .A2(new_n499), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n492), .A2(G2105), .B1(G102), .B2(new_n494), .ZN(new_n972));
  AOI21_X1  g547(.A(G1384), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(KEYINPUT45), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n966), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n965), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G8), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n978));
  INV_X1    g553(.A(G8), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n977), .B(new_n978), .C1(new_n979), .C2(G168), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(KEYINPUT118), .ZN(new_n981));
  NOR2_X1   g556(.A1(G168), .A2(new_n979), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n979), .B1(new_n965), .B2(new_n975), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT118), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT119), .B1(new_n986), .B2(KEYINPUT51), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT119), .ZN(new_n988));
  AOI211_X1 g563(.A(new_n988), .B(new_n978), .C1(new_n981), .C2(new_n985), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n980), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n976), .A2(new_n982), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n968), .B1(new_n500), .B2(new_n949), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(new_n962), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n973), .A2(KEYINPUT45), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n993), .B1(new_n997), .B2(G2078), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n993), .A2(G2078), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  OR3_X1    g575(.A1(new_n970), .A2(new_n974), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n958), .A2(new_n963), .ZN(new_n1002));
  INV_X1    g577(.A(G1961), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n998), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT62), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(G171), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT58), .B(G1341), .Z(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n962), .B2(new_n967), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT116), .B(new_n1008), .C1(new_n962), .C2(new_n967), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n960), .A2(G40), .A3(new_n961), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n967), .A2(new_n969), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT115), .B(G1996), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1013), .A2(new_n996), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1011), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n538), .A2(KEYINPUT117), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1017), .A2(KEYINPUT59), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT59), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n954), .B(KEYINPUT110), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n963), .ZN(new_n1023));
  INV_X1    g598(.A(G1956), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n553), .B(KEYINPUT57), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT56), .B(G2072), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n995), .A2(new_n996), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1956), .B1(new_n1022), .B2(new_n963), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1029), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1026), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(new_n1033), .A3(KEYINPUT61), .ZN(new_n1034));
  INV_X1    g609(.A(G1348), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1002), .A2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n962), .A2(G2067), .A3(new_n967), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n763), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1348), .B1(new_n958), .B2(new_n963), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1040), .A2(new_n1037), .A3(new_n595), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT60), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OR4_X1    g617(.A1(KEYINPUT60), .A2(new_n1040), .A3(new_n763), .A4(new_n1037), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1021), .A2(new_n1034), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1030), .A2(KEYINPUT113), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1025), .A2(new_n1046), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1039), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1048), .B(new_n595), .C1(new_n1040), .C2(new_n1037), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1033), .A2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1045), .B(new_n1047), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1044), .A2(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1005), .A2(G171), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1004), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1002), .A2(KEYINPUT121), .A3(new_n1003), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1013), .A2(KEYINPUT122), .A3(new_n1014), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n994), .B2(new_n962), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1059), .A2(new_n1061), .A3(new_n996), .A4(new_n999), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT123), .ZN(new_n1063));
  OAI211_X1 g638(.A(G40), .B(G160), .C1(new_n973), .C2(new_n968), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1000), .B1(new_n1064), .B2(new_n1060), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n996), .A4(new_n1059), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1058), .A2(new_n1068), .A3(new_n998), .ZN(new_n1069));
  OAI211_X1 g644(.A(KEYINPUT54), .B(new_n1054), .C1(new_n1069), .C2(G301), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1058), .A2(new_n1068), .A3(G301), .A4(new_n998), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1005), .A2(G171), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT61), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1053), .A2(new_n1070), .A3(new_n1075), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n992), .A2(new_n1007), .A3(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n990), .B(new_n991), .C1(new_n1006), .C2(new_n1072), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G166), .A2(new_n979), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT55), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1002), .A2(G2090), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n997), .A2(new_n794), .ZN(new_n1086));
  AOI211_X1 g661(.A(new_n979), .B(new_n1084), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1981), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n566), .B2(KEYINPUT108), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n565), .A2(new_n509), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(G86), .B2(new_n518), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n567), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT108), .ZN(new_n1093));
  OAI21_X1  g668(.A(G1981), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n569), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT109), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1092), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT49), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n962), .A2(new_n967), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(new_n979), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT49), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1092), .A2(new_n1095), .A3(new_n1096), .A4(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n786), .A2(G1976), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1100), .A2(KEYINPUT107), .A3(KEYINPUT52), .A4(new_n1104), .ZN(new_n1105));
  OAI221_X1 g680(.A(G8), .B1(G288), .B2(new_n791), .C1(new_n962), .C2(new_n967), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT107), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(G288), .A2(new_n1108), .A3(new_n791), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1105), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1103), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1087), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1086), .B1(new_n1023), .B2(G2090), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G8), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1084), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT111), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(KEYINPUT111), .A3(new_n1084), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1113), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT124), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1080), .A2(new_n1081), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1087), .A2(new_n1103), .A3(new_n1111), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n977), .A2(G286), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1113), .A2(new_n1118), .A3(new_n1119), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT112), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1115), .A2(KEYINPUT111), .A3(new_n1084), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT111), .B1(new_n1115), .B2(new_n1084), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1130), .A2(KEYINPUT112), .A3(new_n1113), .A4(new_n1124), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1127), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1084), .B1(new_n1134), .B2(new_n979), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1113), .A2(KEYINPUT63), .A3(new_n1124), .A4(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1103), .A2(new_n791), .A3(new_n786), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(G1981), .B2(new_n569), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1133), .A2(new_n1136), .B1(new_n1100), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1122), .A2(new_n1123), .A3(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n707), .B(G2067), .Z(new_n1141));
  INV_X1    g716(.A(new_n690), .ZN(new_n1142));
  INV_X1    g717(.A(G1996), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1014), .A2(new_n962), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT105), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1145), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(G1996), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1147), .B1(new_n690), .B2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n779), .B(new_n782), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(new_n1146), .ZN(new_n1153));
  OR2_X1    g728(.A1(G290), .A2(G1986), .ZN(new_n1154));
  NAND2_X1  g729(.A1(G290), .A2(G1986), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(KEYINPUT104), .A3(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1156), .B(new_n1145), .C1(KEYINPUT104), .C2(new_n1155), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1140), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1149), .B(KEYINPUT46), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1142), .A2(new_n1141), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1160), .B1(new_n1146), .B2(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n1162), .B(KEYINPUT47), .Z(new_n1163));
  NOR3_X1   g738(.A1(new_n1151), .A2(new_n782), .A3(new_n779), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n707), .A2(G2067), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1146), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1154), .A2(new_n1148), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT48), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n1153), .A2(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1163), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1159), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g746(.A1(new_n866), .A2(new_n676), .ZN(new_n1173));
  OAI21_X1  g747(.A(G319), .B1(new_n655), .B2(new_n656), .ZN(new_n1174));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n1175));
  XNOR2_X1  g749(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  AND3_X1   g750(.A1(new_n1176), .A2(new_n642), .A3(KEYINPUT126), .ZN(new_n1177));
  AOI21_X1  g751(.A(KEYINPUT126), .B1(new_n1176), .B2(new_n642), .ZN(new_n1178));
  NOR2_X1   g752(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OR2_X1    g753(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n1180));
  AOI211_X1 g754(.A(new_n1173), .B(new_n1179), .C1(new_n931), .C2(new_n1180), .ZN(G308));
  AOI21_X1  g755(.A(new_n1179), .B1(new_n931), .B2(new_n1180), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n1182), .A2(new_n676), .A3(new_n866), .ZN(G225));
endmodule


