//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n553, new_n555, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1243, new_n1244;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT66), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  OR2_X1    g038(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n467), .A3(G137), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G101), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n466), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OAI221_X1 g057(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n480), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n466), .A2(new_n467), .A3(G138), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n464), .B2(new_n465), .ZN(new_n492));
  AND2_X1   g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n467), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n495), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(KEYINPUT70), .B1(new_n495), .B2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OR3_X1    g073(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n490), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(G543), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n509), .A2(G651), .B1(new_n513), .B2(G50), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n504), .B(new_n506), .C1(new_n510), .C2(new_n511), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT71), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n516), .A2(G88), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n514), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT73), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n526), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n528), .B(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n516), .A2(G89), .A3(new_n520), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n513), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n507), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G651), .B1(new_n513), .B2(G52), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n516), .A2(G90), .A3(new_n520), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n507), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n547), .A2(G651), .B1(new_n513), .B2(G43), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n516), .A2(G81), .A3(new_n520), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G188));
  XOR2_X1   g133(.A(KEYINPUT75), .B(KEYINPUT9), .Z(new_n559));
  NAND4_X1  g134(.A1(new_n559), .A2(G53), .A3(G543), .A4(new_n517), .ZN(new_n560));
  NOR2_X1   g135(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n512), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G651), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n516), .A2(G91), .A3(new_n520), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(G299));
  NAND3_X1  g144(.A1(new_n516), .A2(G87), .A3(new_n520), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n513), .A2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(G288));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n507), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(new_n513), .B2(G48), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n516), .A2(G86), .A3(new_n520), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n576), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(new_n576), .A3(new_n581), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT78), .B1(new_n587), .B2(new_n566), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n516), .A2(G85), .A3(new_n520), .ZN(new_n589));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n507), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n592), .A2(new_n593), .A3(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n513), .A2(G47), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n588), .A2(new_n589), .A3(new_n594), .A4(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n516), .A2(G92), .A3(new_n520), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n507), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g179(.A(KEYINPUT79), .B(new_n600), .C1(new_n507), .C2(new_n601), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n604), .A2(G651), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n513), .A2(G54), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n516), .A2(new_n520), .A3(new_n608), .A4(G92), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n599), .A2(new_n606), .A3(new_n607), .A4(new_n609), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(KEYINPUT80), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(KEYINPUT80), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n597), .B1(new_n613), .B2(G868), .ZN(G284));
  XNOR2_X1  g189(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n611), .A2(new_n612), .ZN(new_n622));
  OAI21_X1  g197(.A(G868), .B1(new_n622), .B2(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n551), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT82), .Z(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g201(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n464), .A2(new_n465), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n631), .A2(G123), .A3(new_n467), .ZN(new_n632));
  OR2_X1    g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(G2104), .B(new_n633), .C1(new_n466), .C2(G111), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n467), .A2(G135), .A3(new_n472), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n630), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT84), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  INV_X1    g216(.A(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2430), .Z(new_n644));
  OAI21_X1  g219(.A(KEYINPUT14), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT83), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(new_n644), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n648), .B1(new_n646), .B2(new_n649), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT16), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  OR3_X1    g229(.A1(new_n650), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n650), .B2(new_n651), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n640), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT85), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n640), .A3(new_n656), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(G401));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT86), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT17), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n665), .B2(new_n664), .ZN(new_n672));
  INV_X1    g247(.A(new_n666), .ZN(new_n673));
  OR3_X1    g248(.A1(new_n664), .A2(new_n667), .A3(new_n665), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT88), .B(G2096), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n683), .A2(new_n685), .A3(new_n687), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n690), .B(new_n691), .C1(new_n689), .C2(new_n688), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n692), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT89), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G4), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n613), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(KEYINPUT93), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT93), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n704), .B(new_n701), .C1(new_n613), .C2(new_n700), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G1348), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n703), .A2(G1348), .A3(new_n705), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n700), .A2(G21), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G168), .B2(new_n700), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(KEYINPUT96), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(KEYINPUT96), .ZN(new_n714));
  OAI21_X1  g289(.A(G1966), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT97), .ZN(new_n716));
  NAND2_X1  g291(.A1(G171), .A2(G16), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G5), .B2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G1961), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n636), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G29), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT30), .B(G28), .Z(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(G29), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n631), .A2(G129), .A3(new_n467), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT26), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(KEYINPUT95), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n731), .A2(new_n472), .A3(G105), .A4(G2104), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n467), .A2(G141), .A3(new_n472), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n725), .A2(new_n728), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  MUX2_X1   g310(.A(G32), .B(new_n735), .S(G29), .Z(new_n736));
  XOR2_X1   g311(.A(KEYINPUT27), .B(G1996), .Z(new_n737));
  AOI21_X1  g312(.A(new_n724), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G1341), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n551), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G16), .B2(G19), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n720), .B(new_n738), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n739), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n719), .B2(new_n718), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT31), .B(G11), .Z(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G27), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G164), .B2(new_n746), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2078), .ZN(new_n749));
  NOR4_X1   g324(.A1(new_n742), .A2(new_n744), .A3(new_n745), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n736), .A2(new_n737), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n713), .A2(new_n714), .ZN(new_n752));
  INV_X1    g327(.A(G1966), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT99), .B(KEYINPUT23), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n700), .A2(G20), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n617), .B2(new_n700), .ZN(new_n758));
  INV_X1    g333(.A(G1956), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT94), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(G115), .A2(G2104), .ZN(new_n764));
  INV_X1    g339(.A(G127), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n480), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(KEYINPUT94), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(new_n631), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT25), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n484), .A2(G139), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  MUX2_X1   g348(.A(G33), .B(new_n773), .S(G29), .Z(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G2072), .Z(new_n775));
  NAND4_X1  g350(.A1(new_n750), .A2(new_n754), .A3(new_n760), .A4(new_n775), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n710), .A2(new_n716), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n746), .A2(G26), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n631), .A2(G128), .A3(new_n467), .ZN(new_n779));
  OR2_X1    g354(.A1(G104), .A2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(G2104), .B(new_n780), .C1(new_n466), .C2(G116), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n467), .A2(G140), .A3(new_n472), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n778), .B1(new_n783), .B2(new_n746), .ZN(new_n784));
  MUX2_X1   g359(.A(new_n778), .B(new_n784), .S(KEYINPUT28), .Z(new_n785));
  INV_X1    g360(.A(G2067), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(KEYINPUT24), .A2(G34), .ZN(new_n788));
  NAND2_X1  g363(.A1(KEYINPUT24), .A2(G34), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n788), .A2(new_n746), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G160), .B2(new_n746), .ZN(new_n791));
  INV_X1    g366(.A(G2084), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G35), .ZN(new_n794));
  OAI21_X1  g369(.A(KEYINPUT98), .B1(new_n794), .B2(G29), .ZN(new_n795));
  OR3_X1    g370(.A1(new_n794), .A2(KEYINPUT98), .A3(G29), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n795), .B(new_n796), .C1(G162), .C2(new_n746), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT29), .B(G2090), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n777), .A2(new_n787), .A3(new_n793), .A4(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G290), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G16), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G16), .B2(G24), .ZN(new_n803));
  INV_X1    g378(.A(G1986), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n481), .A2(G119), .ZN(new_n808));
  OAI221_X1 g383(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n484), .A2(G131), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G29), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G25), .B2(G29), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT35), .B(G1991), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT90), .Z(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n814), .A2(new_n817), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n807), .A2(new_n819), .A3(new_n820), .A4(KEYINPUT92), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n700), .A2(G22), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G166), .B2(new_n700), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(G1971), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n700), .A2(G23), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n700), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT33), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G1976), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(KEYINPUT33), .ZN(new_n830));
  INV_X1    g405(.A(G1976), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n823), .A2(G1971), .ZN(new_n833));
  AND4_X1   g408(.A1(new_n824), .A2(new_n829), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n585), .A2(G16), .ZN(new_n835));
  NOR2_X1   g410(.A1(G6), .A2(G16), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT32), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT32), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n835), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G1981), .ZN(new_n843));
  INV_X1    g418(.A(G1981), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n839), .A2(new_n844), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n834), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n847), .B1(new_n834), .B2(new_n846), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n805), .B(new_n821), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT36), .ZN(new_n852));
  INV_X1    g427(.A(new_n821), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n834), .A2(new_n846), .ZN(new_n854));
  INV_X1    g429(.A(new_n847), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n853), .B1(new_n856), .B2(new_n848), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT36), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n858), .A3(new_n805), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n800), .B1(new_n852), .B2(new_n859), .ZN(G311));
  INV_X1    g435(.A(new_n710), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n776), .A2(new_n716), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n861), .A2(new_n862), .A3(new_n793), .A4(new_n799), .ZN(new_n863));
  INV_X1    g438(.A(new_n787), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n851), .A2(KEYINPUT36), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n858), .B1(new_n857), .B2(new_n805), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(G150));
  NAND2_X1  g443(.A1(new_n613), .A2(G559), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  XOR2_X1   g445(.A(KEYINPUT101), .B(G93), .Z(new_n871));
  NAND3_X1  g446(.A1(new_n516), .A2(new_n520), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n513), .A2(G55), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n504), .A2(new_n506), .A3(G67), .ZN(new_n874));
  NAND2_X1  g449(.A1(G80), .A2(G543), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT100), .B1(new_n876), .B2(G651), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n878));
  AOI211_X1 g453(.A(new_n878), .B(new_n566), .C1(new_n874), .C2(new_n875), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n872), .B(new_n873), .C1(new_n877), .C2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT102), .ZN(new_n881));
  INV_X1    g456(.A(new_n875), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n518), .B2(G67), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n878), .B1(new_n883), .B2(new_n566), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n876), .A2(KEYINPUT100), .A3(G651), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n886), .A2(new_n887), .A3(new_n872), .A4(new_n873), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n881), .A2(new_n551), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n551), .B1(new_n881), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n870), .B(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(KEYINPUT103), .A3(KEYINPUT39), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n895));
  AOI21_X1  g470(.A(G860), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n892), .B2(new_n895), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n880), .A2(G860), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT104), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(G145));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n500), .B(new_n628), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n484), .A2(G142), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n481), .A2(G130), .ZN(new_n910));
  OAI21_X1  g485(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n913), .B(new_n914), .C1(G118), .C2(new_n466), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n484), .A2(KEYINPUT106), .A3(G142), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n909), .A2(new_n910), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n783), .A2(new_n735), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n728), .A2(new_n734), .A3(new_n733), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n725), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n918), .A2(new_n921), .A3(new_n811), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n811), .B1(new_n918), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n917), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n918), .A2(new_n921), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n812), .ZN(new_n926));
  INV_X1    g501(.A(new_n917), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n918), .A2(new_n921), .A3(new_n811), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n470), .ZN(new_n931));
  INV_X1    g506(.A(new_n474), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n721), .ZN(new_n934));
  NAND2_X1  g509(.A1(G160), .A2(new_n636), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n486), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n935), .A3(G162), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n768), .A2(new_n631), .B1(G139), .B2(new_n484), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n940), .B2(new_n771), .ZN(new_n941));
  AND4_X1   g516(.A1(new_n939), .A2(new_n769), .A3(new_n771), .A4(new_n772), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n937), .B(new_n938), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n773), .A2(KEYINPUT105), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n939), .A3(new_n771), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n934), .A2(new_n935), .A3(G162), .ZN(new_n946));
  AOI21_X1  g521(.A(G162), .B1(new_n934), .B2(new_n935), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n944), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n930), .A2(new_n943), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n930), .B1(new_n943), .B2(new_n948), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n906), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n943), .A2(new_n948), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n924), .A2(new_n929), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n905), .A3(new_n949), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n952), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n952), .A2(KEYINPUT108), .A3(new_n953), .A4(new_n957), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n960), .B2(new_n962), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n904), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n960), .A2(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(KEYINPUT40), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n965), .A2(new_n969), .ZN(G395));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n613), .A2(new_n891), .A3(new_n620), .ZN(new_n972));
  OAI22_X1  g547(.A1(new_n622), .A2(G559), .B1(new_n889), .B2(new_n890), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n599), .A2(new_n609), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n975), .A2(new_n617), .A3(new_n607), .A4(new_n606), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n610), .A2(G299), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n971), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n980), .A3(KEYINPUT41), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n610), .A2(G299), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n610), .A2(G299), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT41), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT41), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n976), .A2(new_n985), .A3(new_n977), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(KEYINPUT111), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n974), .A2(new_n981), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n978), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n972), .A2(KEYINPUT110), .A3(new_n973), .A4(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n979), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT42), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n514), .A2(new_n993), .A3(new_n521), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n993), .B1(new_n514), .B2(new_n521), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n583), .B(new_n584), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n996), .ZN(new_n998));
  INV_X1    g573(.A(new_n584), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n998), .B(new_n994), .C1(new_n999), .C2(new_n582), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n588), .A2(new_n594), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n589), .A2(new_n595), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n573), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n826), .A2(G290), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT113), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1001), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1007), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(new_n997), .A3(new_n1000), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT42), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n979), .A2(new_n988), .A3(new_n1014), .A4(new_n990), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n992), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1013), .B1(new_n992), .B2(new_n1015), .ZN(new_n1017));
  OAI21_X1  g592(.A(G868), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G868), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n880), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(G295));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1020), .ZN(G331));
  XNOR2_X1  g597(.A(G171), .B(G286), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n889), .B2(new_n890), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n884), .A2(new_n885), .B1(G55), .B2(new_n513), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n887), .B1(new_n1025), .B2(new_n872), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n880), .A2(KEYINPUT102), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n550), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n881), .A2(new_n551), .A3(new_n888), .ZN(new_n1029));
  XNOR2_X1  g604(.A(G286), .B(G301), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(new_n981), .A3(new_n987), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1024), .A2(new_n1031), .A3(new_n989), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1013), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n953), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1013), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT43), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT114), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1034), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1024), .A2(new_n1031), .B1(new_n984), .B2(new_n986), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(new_n1035), .A3(new_n953), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1044), .A2(KEYINPUT43), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(KEYINPUT43), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1039), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT43), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1051), .B2(new_n1044), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT44), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1054), .ZN(G397));
  NAND3_X1  g630(.A1(new_n931), .A2(new_n932), .A3(G40), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1384), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT45), .B1(new_n500), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n783), .A2(new_n786), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n919), .A2(G2067), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n811), .A2(new_n816), .ZN(new_n1064));
  INV_X1    g639(.A(G1996), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n735), .B(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1060), .B1(new_n1067), .B2(new_n1061), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1060), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1063), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(new_n735), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(KEYINPUT46), .A3(new_n1065), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT46), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1060), .B2(G1996), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  XOR2_X1   g650(.A(new_n1075), .B(KEYINPUT47), .Z(new_n1076));
  NAND2_X1  g651(.A1(new_n801), .A2(new_n804), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(new_n1060), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT127), .ZN(new_n1079));
  XOR2_X1   g654(.A(new_n1079), .B(KEYINPUT48), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n812), .A2(new_n817), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1081), .A2(new_n1064), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1069), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n1068), .B(new_n1076), .C1(new_n1080), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n500), .A2(new_n1058), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT45), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n1058), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1057), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n753), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1056), .B1(new_n1088), .B2(KEYINPUT50), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n500), .A2(new_n1095), .A3(new_n1058), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(new_n792), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1087), .B1(new_n1098), .B2(G286), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1093), .A2(G168), .A3(new_n1097), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G8), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1087), .B1(new_n1100), .B2(G8), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT62), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1971), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1092), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(G2090), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(G303), .A2(G8), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT55), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(G8), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1096), .A2(KEYINPUT120), .ZN(new_n1114));
  INV_X1    g689(.A(G2090), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n500), .A2(new_n1116), .A3(new_n1095), .A4(new_n1058), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1094), .A2(new_n1114), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1113), .B1(new_n1106), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1112), .B1(new_n1111), .B2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(G160), .A2(new_n500), .A3(G40), .A4(new_n1058), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(G8), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT115), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(new_n1124), .A3(G8), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n580), .A2(new_n581), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n566), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(G1981), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n580), .A2(new_n1130), .A3(G1981), .A4(new_n581), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(KEYINPUT119), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT49), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1126), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n570), .A2(G1976), .A3(new_n571), .A4(new_n572), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT116), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1121), .A2(new_n1124), .A3(G8), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1124), .B1(new_n1121), .B2(G8), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT52), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT117), .B(G1976), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT52), .B1(G288), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1126), .A2(new_n1146), .A3(new_n1140), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1138), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1120), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1091), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1150), .A2(new_n1059), .A3(new_n1056), .ZN(new_n1151));
  INV_X1    g726(.A(G2078), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(KEYINPUT53), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1092), .B2(G2078), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1107), .A2(new_n719), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1153), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(G301), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1103), .ZN(new_n1159));
  AOI21_X1  g734(.A(G168), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1160));
  OAI211_X1 g735(.A(G8), .B(new_n1100), .C1(new_n1160), .C2(new_n1087), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1104), .A2(new_n1149), .A3(new_n1158), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(G288), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1138), .A2(new_n831), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n580), .A2(new_n844), .A3(new_n581), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1166), .A2(new_n1167), .B1(new_n1125), .B2(new_n1123), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1108), .A2(KEYINPUT121), .A3(G8), .A4(new_n1110), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1110), .A2(KEYINPUT121), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1088), .A2(KEYINPUT50), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1171), .A2(new_n1057), .A3(new_n1096), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1172), .A2(new_n1115), .B1(new_n1092), .B2(new_n1105), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1170), .B1(new_n1173), .B2(new_n1113), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1169), .A2(new_n1174), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1138), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1101), .A2(G286), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1168), .B1(new_n1178), .B2(KEYINPUT63), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1119), .A2(new_n1111), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1098), .A2(new_n1181), .A3(G8), .A4(G168), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1112), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1176), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1164), .A2(new_n1179), .A3(new_n1184), .ZN(new_n1185));
  OR3_X1    g760(.A1(new_n1092), .A2(KEYINPUT124), .A3(G1996), .ZN(new_n1186));
  XOR2_X1   g761(.A(KEYINPUT58), .B(G1341), .Z(new_n1187));
  NAND2_X1  g762(.A1(new_n1121), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT124), .B1(new_n1092), .B2(G1996), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1186), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n551), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT59), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1190), .A2(new_n1193), .A3(new_n551), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g770(.A(G299), .B(KEYINPUT122), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT57), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1094), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n759), .ZN(new_n1201));
  XNOR2_X1  g776(.A(KEYINPUT56), .B(G2072), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1151), .A2(new_n1202), .ZN(new_n1203));
  AND3_X1   g778(.A1(new_n1201), .A2(KEYINPUT123), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(KEYINPUT123), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1199), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1198), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1206), .A2(new_n1208), .A3(KEYINPUT61), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n1210));
  AND2_X1   g785(.A1(new_n1207), .A2(new_n1198), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1207), .A2(new_n1198), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1210), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1121), .A2(G2067), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1214), .B1(new_n1107), .B2(new_n707), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1215), .B1(new_n613), .B2(KEYINPUT60), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n613), .A2(KEYINPUT60), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1216), .B(new_n1217), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1195), .A2(new_n1209), .A3(new_n1213), .A4(new_n1218), .ZN(new_n1219));
  OR3_X1    g794(.A1(new_n1211), .A2(new_n622), .A3(new_n1215), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1219), .A2(new_n1206), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1151), .A2(new_n1223), .A3(G2078), .ZN(new_n1224));
  AND2_X1   g799(.A1(new_n1224), .A2(new_n1156), .ZN(new_n1225));
  NAND4_X1  g800(.A1(new_n1151), .A2(KEYINPUT125), .A3(KEYINPUT53), .A4(new_n1152), .ZN(new_n1226));
  NAND4_X1  g801(.A1(new_n1225), .A2(KEYINPUT126), .A3(new_n1155), .A4(new_n1226), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1226), .A2(new_n1224), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1228));
  INV_X1    g803(.A(KEYINPUT126), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1227), .A2(new_n1230), .A3(G171), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT54), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1232), .B1(new_n1157), .B2(G301), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g809(.A1(new_n1228), .A2(G171), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1232), .B1(new_n1158), .B2(new_n1235), .ZN(new_n1236));
  AND4_X1   g811(.A1(new_n1222), .A2(new_n1234), .A3(new_n1149), .A4(new_n1236), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1185), .B1(new_n1221), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g813(.A(new_n1084), .B1(G1986), .B2(G290), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1060), .B1(new_n1239), .B2(new_n1077), .ZN(new_n1240));
  OAI21_X1  g815(.A(new_n1086), .B1(new_n1238), .B2(new_n1240), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g816(.A(G227), .B(G229), .C1(new_n960), .C2(new_n962), .ZN(new_n1243));
  AOI21_X1  g817(.A(new_n462), .B1(new_n658), .B2(new_n660), .ZN(new_n1244));
  AND3_X1   g818(.A1(new_n1048), .A2(new_n1243), .A3(new_n1244), .ZN(G308));
  NAND3_X1  g819(.A1(new_n1048), .A2(new_n1243), .A3(new_n1244), .ZN(G225));
endmodule


