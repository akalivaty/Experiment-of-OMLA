//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G113gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT67), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n208), .B1(new_n205), .B2(new_n207), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n203), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n206), .A2(KEYINPUT68), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G120gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n204), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT69), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(new_n206), .B2(G113gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n210), .B(new_n202), .C1(new_n217), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n224), .B1(new_n227), .B2(KEYINPUT2), .ZN(new_n228));
  INV_X1    g027(.A(G148gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G141gat), .ZN(new_n230));
  INV_X1    g029(.A(G141gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G148gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT77), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(new_n230), .B2(new_n232), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n228), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n232), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G155gat), .B(G162gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT4), .B1(new_n223), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n240), .B1(new_n237), .B2(new_n238), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n231), .A2(G148gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n229), .A2(G141gat), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT77), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n245), .B1(new_n250), .B2(new_n228), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n251), .A2(new_n252), .A3(new_n213), .A4(new_n222), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n244), .A2(KEYINPUT79), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n251), .A2(new_n255), .B1(new_n213), .B2(new_n222), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT78), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n257), .B1(new_n243), .B2(KEYINPUT3), .ZN(new_n258));
  AOI211_X1 g057(.A(KEYINPUT78), .B(new_n255), .C1(new_n236), .C2(new_n242), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G225gat), .A2(G233gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n223), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT79), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n262), .A2(new_n263), .A3(new_n252), .A4(new_n251), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n254), .A2(new_n260), .A3(new_n261), .A4(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT5), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n223), .B(new_n243), .ZN(new_n267));
  INV_X1    g066(.A(new_n261), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT78), .B1(new_n251), .B2(new_n255), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n243), .A2(new_n257), .A3(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n268), .B1(new_n273), .B2(new_n256), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT80), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n275), .B(KEYINPUT4), .C1(new_n223), .C2(new_n243), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n244), .A2(KEYINPUT80), .A3(new_n253), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n274), .A2(new_n266), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT0), .B(G57gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(G85gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(G1gat), .B(G29gat), .ZN(new_n282));
  XOR2_X1   g081(.A(new_n281), .B(new_n282), .Z(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n279), .A2(KEYINPUT6), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT81), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n279), .A2(new_n284), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n270), .A2(new_n278), .A3(new_n283), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n283), .B1(new_n270), .B2(new_n278), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n292), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n287), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G211gat), .ZN(new_n295));
  INV_X1    g094(.A(G218gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G197gat), .ZN(new_n298));
  INV_X1    g097(.A(G204gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(G197gat), .A2(G204gat), .ZN(new_n301));
  OAI22_X1  g100(.A1(KEYINPUT22), .A2(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G211gat), .B(G218gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G226gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G183gat), .ZN(new_n307));
  INV_X1    g106(.A(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(KEYINPUT24), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT23), .ZN(new_n313));
  INV_X1    g112(.A(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n310), .A2(KEYINPUT24), .ZN(new_n318));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT23), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n311), .A2(new_n317), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT64), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(KEYINPUT64), .A3(new_n322), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT65), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT65), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n329), .B1(G169gat), .B2(G176gat), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n327), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(new_n322), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n332), .A2(new_n311), .A3(new_n318), .A4(new_n317), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n325), .A2(new_n326), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT28), .ZN(new_n335));
  NAND2_X1  g134(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n335), .B(new_n308), .C1(new_n336), .C2(KEYINPUT27), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(KEYINPUT27), .B2(new_n336), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT27), .B(G183gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n308), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(KEYINPUT28), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n316), .A2(KEYINPUT26), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n328), .A2(new_n330), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n312), .B(new_n342), .C1(new_n343), .C2(KEYINPUT26), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n344), .A3(new_n310), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n334), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n306), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n305), .B1(new_n334), .B2(new_n345), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n304), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n306), .ZN(new_n351));
  INV_X1    g150(.A(new_n303), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n302), .B(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT29), .B1(new_n334), .B2(new_n345), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n351), .B(new_n353), .C1(new_n306), .C2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356));
  INV_X1    g155(.A(G64gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G92gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n350), .A2(new_n355), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n350), .A2(new_n355), .A3(KEYINPUT30), .A4(new_n361), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n361), .B1(new_n350), .B2(new_n355), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT75), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n368));
  AOI211_X1 g167(.A(new_n368), .B(new_n361), .C1(new_n350), .C2(new_n355), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n364), .B(new_n365), .C1(new_n367), .C2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT82), .B1(new_n294), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n287), .A2(new_n291), .A3(new_n293), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n366), .B(KEYINPUT75), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n364), .A2(new_n365), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT31), .B(G22gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G228gat), .A2(G233gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n304), .A2(KEYINPUT29), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n243), .B1(new_n380), .B2(KEYINPUT3), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n251), .B2(new_n255), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n353), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(G50gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n353), .A2(new_n347), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n251), .B1(new_n385), .B2(new_n255), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n382), .A2(new_n353), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G50gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n379), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n383), .A2(G50gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n389), .ZN(new_n394));
  INV_X1    g193(.A(new_n379), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n391), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n392), .B1(new_n391), .B2(new_n396), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n326), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n311), .A2(new_n318), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n319), .B1(KEYINPUT23), .B2(new_n312), .ZN(new_n402));
  NOR4_X1   g201(.A1(new_n401), .A2(new_n331), .A3(new_n322), .A4(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT64), .B1(new_n321), .B2(new_n322), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n400), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n341), .A2(new_n310), .A3(new_n344), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n262), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G227gat), .ZN(new_n408));
  INV_X1    g207(.A(G233gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n334), .A2(new_n223), .A3(new_n345), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT32), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  XOR2_X1   g214(.A(G71gat), .B(G99gat), .Z(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT70), .ZN(new_n417));
  XOR2_X1   g216(.A(G15gat), .B(G43gat), .Z(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n413), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n412), .B(KEYINPUT32), .C1(new_n414), .C2(new_n419), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n411), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n223), .B1(new_n334), .B2(new_n345), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n425), .B1(new_n428), .B2(new_n410), .ZN(new_n429));
  OAI221_X1 g228(.A(new_n424), .B1(new_n408), .B2(new_n409), .C1(new_n426), .C2(new_n427), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT72), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n421), .A2(new_n422), .A3(new_n430), .A4(new_n429), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n423), .A2(KEYINPUT72), .A3(new_n431), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n399), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n371), .A2(new_n376), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT35), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(KEYINPUT85), .A3(KEYINPUT35), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n370), .A2(KEYINPUT83), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n374), .A2(new_n375), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n432), .A2(KEYINPUT73), .A3(new_n434), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT73), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n423), .A2(new_n448), .A3(new_n431), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT35), .ZN(new_n452));
  INV_X1    g251(.A(new_n399), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n372), .A4(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n441), .A2(new_n442), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n350), .A2(new_n355), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT84), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT38), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n350), .A2(new_n355), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT37), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n360), .A3(new_n457), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n459), .B(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n294), .A3(new_n362), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT39), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n267), .A2(new_n268), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n277), .A2(new_n260), .A3(new_n276), .ZN(new_n467));
  AOI211_X1 g266(.A(new_n465), .B(new_n466), .C1(new_n268), .C2(new_n467), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n467), .A2(new_n465), .A3(new_n268), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n468), .A2(new_n284), .A3(new_n469), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n470), .A2(KEYINPUT40), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n292), .B1(new_n470), .B2(KEYINPUT40), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n443), .A2(new_n445), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n464), .A2(new_n473), .A3(new_n453), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n371), .A2(new_n376), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n399), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n435), .A2(new_n436), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT36), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n478), .B(KEYINPUT74), .C1(KEYINPUT36), .C2(new_n450), .ZN(new_n479));
  OR3_X1    g278(.A1(new_n450), .A2(KEYINPUT74), .A3(KEYINPUT36), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n474), .A2(new_n476), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n455), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT11), .B(G169gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(G197gat), .ZN(new_n484));
  XOR2_X1   g283(.A(G113gat), .B(G141gat), .Z(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT12), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(KEYINPUT90), .A2(KEYINPUT18), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT88), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT16), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(G1gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n491), .B(KEYINPUT88), .ZN(new_n496));
  INV_X1    g295(.A(G1gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(KEYINPUT89), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(G8gat), .ZN(new_n500));
  INV_X1    g299(.A(G8gat), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n495), .A2(KEYINPUT89), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G29gat), .ZN(new_n504));
  INV_X1    g303(.A(G36gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT14), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT14), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n506), .B(new_n508), .C1(new_n504), .C2(new_n505), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n389), .A2(G43gat), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT86), .B(G43gat), .Z(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G50gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n389), .A2(G43gat), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n510), .A2(KEYINPUT15), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT87), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n514), .A2(new_n520), .A3(new_n517), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n509), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT17), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n519), .A2(new_n521), .A3(new_n525), .A4(new_n522), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n503), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n503), .A2(new_n523), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n490), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n530), .ZN(new_n532));
  NOR4_X1   g331(.A1(new_n527), .A2(new_n528), .A3(new_n532), .A4(new_n489), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n530), .B(KEYINPUT13), .ZN(new_n535));
  INV_X1    g334(.A(new_n503), .ZN(new_n536));
  INV_X1    g335(.A(new_n523), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n503), .A2(new_n523), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n488), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  NOR4_X1   g341(.A1(new_n531), .A2(new_n533), .A3(new_n540), .A4(new_n487), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  OR2_X1    g347(.A1(G71gat), .A2(G78gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT9), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n548), .B(new_n549), .C1(new_n545), .C2(new_n550), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT7), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  INV_X1    g357(.A(G85gat), .ZN(new_n559));
  AOI22_X1  g358(.A1(KEYINPUT8), .A2(new_n558), .B1(new_n559), .B2(new_n359), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n556), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G99gat), .B(G106gat), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n562), .B2(new_n563), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n554), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT10), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n567), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n564), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n552), .A2(new_n573), .A3(new_n553), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n552), .B2(new_n553), .ZN(new_n575));
  OAI211_X1 g374(.A(KEYINPUT10), .B(new_n565), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT98), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n578), .B1(new_n568), .B2(new_n571), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT100), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(KEYINPUT98), .ZN(new_n585));
  XNOR2_X1  g384(.A(G176gat), .B(G204gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(G148gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT99), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n206), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n577), .B2(new_n578), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n585), .B(new_n589), .C1(new_n592), .C2(new_n581), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT100), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n589), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n578), .B(KEYINPUT101), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n598), .B1(new_n572), .B2(new_n576), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n596), .B1(new_n599), .B2(new_n581), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n544), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n554), .A2(KEYINPUT21), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(new_n295), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n604), .B(new_n606), .Z(new_n607));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT21), .B1(new_n574), .B2(new_n575), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n307), .B1(new_n536), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n536), .A2(new_n307), .A3(new_n610), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n612), .A2(G231gat), .A3(G233gat), .A4(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n612), .A2(new_n613), .B1(G231gat), .B2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  INV_X1    g418(.A(new_n616), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(new_n620), .B2(new_n614), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n609), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n617), .B1(new_n615), .B2(new_n616), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n620), .A2(new_n614), .A3(new_n619), .ZN(new_n624));
  INV_X1    g423(.A(new_n609), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(G232gat), .A2(G233gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(KEYINPUT41), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n565), .B1(new_n524), .B2(new_n526), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(KEYINPUT41), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n537), .A2(new_n564), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n630), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NOR4_X1   g436(.A1(new_n631), .A2(new_n635), .A3(KEYINPUT96), .A4(new_n633), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n629), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n524), .A2(new_n526), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n564), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n632), .A3(new_n636), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT96), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n630), .A3(new_n636), .ZN(new_n644));
  INV_X1    g443(.A(new_n629), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n639), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n639), .B2(new_n646), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n603), .A2(new_n627), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n482), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n294), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G1gat), .ZN(G1324gat));
  INV_X1    g455(.A(new_n654), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n446), .ZN(new_n658));
  NAND2_X1  g457(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n494), .A2(new_n501), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT42), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n501), .B2(new_n658), .ZN(G1325gat));
  AOI21_X1  g462(.A(G15gat), .B1(new_n654), .B2(new_n450), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n479), .A2(new_n480), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n666), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g466(.A1(new_n654), .A2(new_n399), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT43), .B(G22gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  INV_X1    g469(.A(new_n652), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n455), .B2(new_n481), .ZN(new_n672));
  INV_X1    g471(.A(new_n627), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n603), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n675), .A2(G29gat), .A3(new_n372), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT45), .Z(new_n677));
  AND3_X1   g476(.A1(new_n438), .A2(KEYINPUT85), .A3(KEYINPUT35), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT85), .B1(new_n438), .B2(KEYINPUT35), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n446), .A2(new_n452), .A3(new_n453), .A4(new_n450), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n294), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n481), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n652), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n482), .A2(KEYINPUT102), .A3(KEYINPUT44), .A4(new_n652), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n688), .A2(KEYINPUT103), .A3(new_n294), .A4(new_n674), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n686), .A2(new_n674), .A3(new_n687), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n691), .B2(new_n372), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(G29gat), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n693), .ZN(G1328gat));
  NOR3_X1   g493(.A1(new_n675), .A2(G36gat), .A3(new_n446), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT46), .ZN(new_n696));
  OAI21_X1  g495(.A(G36gat), .B1(new_n691), .B2(new_n446), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1329gat));
  OR3_X1    g497(.A1(new_n691), .A2(KEYINPUT106), .A3(new_n665), .ZN(new_n699));
  INV_X1    g498(.A(new_n511), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT106), .B1(new_n691), .B2(new_n665), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n672), .A2(new_n450), .A3(new_n511), .A4(new_n674), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(KEYINPUT47), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n703), .B(KEYINPUT104), .Z(new_n705));
  OAI21_X1  g504(.A(new_n700), .B1(new_n691), .B2(new_n665), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT47), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI211_X1 g508(.A(KEYINPUT105), .B(KEYINPUT47), .C1(new_n705), .C2(new_n706), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n704), .B1(new_n709), .B2(new_n710), .ZN(G1330gat));
  NOR2_X1   g510(.A1(new_n453), .A2(new_n389), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n686), .A2(new_n687), .A3(new_n674), .A4(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n389), .B1(new_n675), .B2(new_n453), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(KEYINPUT107), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT48), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n713), .A2(KEYINPUT48), .A3(new_n714), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n717), .ZN(G1331gat));
  INV_X1    g519(.A(new_n601), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n455), .B2(new_n481), .ZN(new_n722));
  INV_X1    g521(.A(new_n544), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n627), .A2(new_n723), .A3(new_n652), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n294), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G57gat), .ZN(G1332gat));
  INV_X1    g527(.A(new_n446), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT49), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(new_n357), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT109), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n357), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n725), .B2(new_n665), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n726), .A2(new_n450), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(G71gat), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g538(.A1(new_n726), .A2(new_n399), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n673), .A2(new_n723), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n672), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(new_n601), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n559), .A3(new_n294), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n686), .A2(new_n687), .A3(new_n601), .A4(new_n742), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n748), .A2(new_n749), .A3(new_n372), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n748), .B2(new_n372), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(G85gat), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n747), .A2(new_n752), .ZN(G1336gat));
  NOR2_X1   g552(.A1(new_n446), .A2(G92gat), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT52), .B1(new_n746), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G92gat), .B1(new_n748), .B2(new_n446), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OR2_X1    g556(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n758));
  AND4_X1   g557(.A1(new_n482), .A2(new_n652), .A3(new_n742), .A4(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n672), .B2(new_n742), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n601), .B(new_n754), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(new_n756), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT52), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n757), .A2(new_n766), .ZN(G1337gat));
  INV_X1    g566(.A(G99gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n746), .A2(new_n768), .A3(new_n450), .ZN(new_n769));
  OAI21_X1  g568(.A(G99gat), .B1(new_n748), .B2(new_n665), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1338gat));
  OR3_X1    g570(.A1(new_n748), .A2(KEYINPUT116), .A3(new_n453), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT116), .B1(new_n748), .B2(new_n453), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(G106gat), .A3(new_n773), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n721), .A2(G106gat), .A3(new_n453), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT113), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT53), .B1(new_n745), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G106gat), .B1(new_n748), .B2(new_n453), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n776), .B1(new_n759), .B2(new_n760), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT114), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n782), .B(new_n776), .C1(new_n759), .C2(new_n760), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n784), .A2(new_n785), .A3(KEYINPUT53), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n784), .B2(KEYINPUT53), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n778), .B1(new_n786), .B2(new_n787), .ZN(G1339gat));
  NAND3_X1  g587(.A1(new_n572), .A2(new_n576), .A3(new_n598), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n579), .A2(KEYINPUT54), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n589), .B1(new_n599), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n790), .A2(KEYINPUT55), .A3(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n595), .B(new_n798), .C1(new_n542), .C2(new_n543), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n532), .B1(new_n527), .B2(new_n528), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n538), .A2(new_n539), .A3(new_n535), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n486), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n543), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n601), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n671), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n797), .B1(new_n594), .B2(new_n590), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n639), .A2(new_n646), .ZN(new_n808));
  INV_X1    g607(.A(new_n649), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n639), .A2(new_n646), .A3(new_n649), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n807), .A2(new_n810), .A3(new_n811), .A4(new_n803), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n652), .A2(KEYINPUT117), .A3(new_n803), .A4(new_n807), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n806), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n627), .ZN(new_n817));
  NOR4_X1   g616(.A1(new_n627), .A2(new_n723), .A3(new_n652), .A4(new_n601), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n450), .A2(new_n453), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n729), .A2(new_n372), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n544), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT118), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n818), .B1(new_n816), .B2(new_n627), .ZN(new_n827));
  INV_X1    g626(.A(new_n437), .ZN(new_n828));
  NOR4_X1   g627(.A1(new_n827), .A2(new_n372), .A3(new_n729), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n204), .A3(new_n723), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n830), .ZN(G1340gat));
  NAND2_X1  g630(.A1(new_n214), .A2(new_n216), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n832), .A3(new_n601), .ZN(new_n833));
  OAI21_X1  g632(.A(G120gat), .B1(new_n824), .B2(new_n721), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1341gat));
  AOI21_X1  g634(.A(G127gat), .B1(new_n829), .B2(new_n673), .ZN(new_n836));
  INV_X1    g635(.A(new_n824), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n673), .A2(G127gat), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(G1342gat));
  INV_X1    g638(.A(G134gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n829), .A2(new_n840), .A3(new_n652), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n837), .B2(new_n652), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n841), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n844), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT120), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n844), .A2(new_n851), .A3(new_n847), .A4(new_n848), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1343gat));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n827), .B2(new_n453), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT121), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n652), .B1(new_n805), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n857), .B2(new_n805), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n814), .A2(new_n815), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n673), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT57), .B(new_n399), .C1(new_n861), .C2(new_n818), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n863), .B(new_n854), .C1(new_n827), .C2(new_n453), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n856), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n665), .A2(new_n823), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n723), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G141gat), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n827), .A2(new_n453), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n870), .A2(new_n231), .A3(new_n723), .A4(new_n866), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n871), .B(KEYINPUT123), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT58), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n868), .A2(KEYINPUT124), .A3(new_n869), .A4(new_n871), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n874), .A2(new_n877), .A3(new_n878), .ZN(G1344gat));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n866), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n880), .B(G148gat), .C1(new_n881), .C2(new_n721), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n673), .B1(new_n859), .B2(new_n812), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n854), .B(new_n399), .C1(new_n883), .C2(new_n818), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT57), .B1(new_n827), .B2(new_n453), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(new_n601), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n229), .B1(new_n887), .B2(new_n866), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n882), .B1(new_n888), .B2(new_n880), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n870), .A2(new_n866), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n229), .A3(new_n601), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1345gat));
  AOI21_X1  g691(.A(G155gat), .B1(new_n890), .B2(new_n673), .ZN(new_n893));
  INV_X1    g692(.A(new_n881), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n627), .A2(new_n225), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(G1346gat));
  AOI21_X1  g695(.A(G162gat), .B1(new_n890), .B2(new_n652), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n671), .A2(new_n226), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n894), .B2(new_n898), .ZN(G1347gat));
  NOR4_X1   g698(.A1(new_n827), .A2(new_n294), .A3(new_n446), .A4(new_n828), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n314), .A3(new_n723), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT125), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n446), .A2(new_n294), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n820), .A2(new_n822), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n544), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n905), .ZN(G1348gat));
  AOI21_X1  g705(.A(G176gat), .B1(new_n900), .B2(new_n601), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n904), .A2(new_n315), .A3(new_n721), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(G1349gat));
  NAND3_X1  g708(.A1(new_n900), .A2(new_n339), .A3(new_n673), .ZN(new_n910));
  OAI21_X1  g709(.A(G183gat), .B1(new_n904), .B2(new_n627), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT126), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n904), .B2(new_n671), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT61), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n308), .A3(new_n652), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1351gat));
  AND2_X1   g718(.A1(new_n665), .A2(new_n903), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n886), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G197gat), .B1(new_n921), .B2(new_n544), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n870), .A2(new_n920), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n298), .A3(new_n723), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1352gat));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n299), .A3(new_n601), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT62), .Z(new_n927));
  AND2_X1   g726(.A1(new_n887), .A2(new_n920), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n299), .ZN(G1353gat));
  NAND3_X1  g728(.A1(new_n886), .A2(new_n673), .A3(new_n920), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(G211gat), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT63), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n923), .A2(new_n295), .A3(new_n673), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(KEYINPUT63), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n932), .A2(KEYINPUT63), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n930), .A2(G211gat), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n934), .A3(new_n937), .ZN(G1354gat));
  OAI21_X1  g737(.A(G218gat), .B1(new_n921), .B2(new_n671), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n296), .A3(new_n652), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1355gat));
endmodule


