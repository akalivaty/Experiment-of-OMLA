//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT69), .Z(G261));
  AOI22_X1  g031(.A1(new_n451), .A2(G567), .B1(new_n454), .B2(G2106), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT71), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT70), .B(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(KEYINPUT70), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND4_X1   g041(.A1(KEYINPUT71), .A2(new_n464), .A3(new_n466), .A4(KEYINPUT3), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n458), .C1(new_n463), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n462), .A2(G2105), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(G2105), .B1(new_n476), .B2(G101), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n468), .A2(new_n477), .ZN(G160));
  NAND3_X1  g053(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(new_n461), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT71), .A4(KEYINPUT3), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n458), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G136), .B2(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n483), .B2(G126), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n488), .B2(G138), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n494), .A2(KEYINPUT72), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(KEYINPUT72), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n496), .A2(new_n497), .A3(G138), .A4(new_n458), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(new_n473), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n493), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G50), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT73), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(new_n502), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  OAI221_X1 g092(.A(new_n505), .B1(new_n514), .B2(new_n515), .C1(new_n516), .C2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  INV_X1    g094(.A(new_n514), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G89), .B1(G51), .B2(new_n504), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT75), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n511), .A2(new_n512), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT74), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n511), .A2(new_n528), .A3(new_n512), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n525), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(new_n504), .A2(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n514), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n527), .A2(new_n529), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  INV_X1    g112(.A(G77), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(new_n506), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n535), .B1(new_n539), .B2(G651), .ZN(G171));
  NAND2_X1  g115(.A1(new_n504), .A2(G43), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n514), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n536), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n543), .B1(new_n546), .B2(G651), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n548), .B(KEYINPUT76), .Z(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n503), .A2(KEYINPUT9), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n503), .B2(new_n554), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n520), .A2(G91), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n517), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  INV_X1    g136(.A(G168), .ZN(G286));
  NAND2_X1  g137(.A1(new_n504), .A2(G49), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n511), .A2(G87), .A3(new_n512), .A4(new_n502), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(G74), .B1(new_n527), .B2(new_n529), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n566), .B2(new_n517), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT77), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n565), .B(new_n569), .C1(new_n566), .C2(new_n517), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G288));
  NAND3_X1  g147(.A1(new_n511), .A2(G61), .A3(new_n512), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(KEYINPUT78), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n573), .A2(KEYINPUT78), .B1(G73), .B2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n517), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n504), .A2(G48), .ZN(new_n577));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n514), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  XNOR2_X1  g156(.A(KEYINPUT80), .B(G85), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n513), .A2(new_n502), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g158(.A(KEYINPUT79), .B(G47), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n504), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT81), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n517), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n587), .B(KEYINPUT82), .C1(new_n517), .C2(new_n588), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G171), .A2(G868), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n513), .A2(G92), .A3(new_n502), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n526), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(G54), .B2(new_n504), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(KEYINPUT83), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(KEYINPUT83), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n594), .B1(new_n605), .B2(G868), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT84), .ZN(G284));
  XOR2_X1   g182(.A(new_n606), .B(KEYINPUT85), .Z(G321));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G299), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G168), .B2(new_n609), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(G168), .B2(new_n609), .ZN(G280));
  INV_X1    g187(.A(G860), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n605), .B1(G559), .B2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT86), .Z(G148));
  INV_X1    g190(.A(new_n547), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n609), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n605), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g195(.A(new_n473), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n476), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n488), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n483), .A2(G123), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(KEYINPUT87), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(KEYINPUT87), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G111), .B2(new_n458), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n626), .B(new_n627), .C1(new_n629), .C2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT88), .B(G2096), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n625), .A2(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT91), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT90), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT14), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(G14), .B1(new_n644), .B2(new_n650), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n657), .B2(new_n654), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n660), .B(new_n662), .Z(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n670), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  AOI211_X1 g250(.A(new_n672), .B(new_n675), .C1(new_n667), .C2(new_n671), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G229));
  INV_X1    g257(.A(G290), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G16), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G16), .B2(G24), .ZN(new_n685));
  INV_X1    g260(.A(G1986), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n688), .ZN(new_n690));
  INV_X1    g265(.A(G1971), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G23), .B(new_n567), .S(G16), .Z(new_n693));
  XOR2_X1   g268(.A(KEYINPUT33), .B(G1976), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NOR2_X1   g271(.A1(G6), .A2(G16), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n580), .B2(G16), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n692), .A2(new_n695), .A3(new_n696), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT34), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n685), .A2(new_n686), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n488), .A2(G131), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n483), .A2(G119), .ZN(new_n705));
  OR2_X1    g280(.A1(G95), .A2(G2105), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n706), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT94), .B(G29), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G25), .B(new_n708), .S(new_n710), .Z(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT35), .B(G1991), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR4_X1   g288(.A1(new_n687), .A2(new_n702), .A3(new_n703), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT36), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT98), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT26), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(KEYINPUT26), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n718), .A2(new_n719), .B1(G105), .B2(new_n476), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n488), .A2(G141), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n483), .A2(G129), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n725), .B2(G32), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT27), .B(G1996), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT99), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n725), .A2(G33), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT25), .Z(new_n733));
  AOI22_X1  g308(.A1(new_n621), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n458), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G139), .B2(new_n488), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(new_n725), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(G2072), .Z(new_n738));
  INV_X1    g313(.A(G2084), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT24), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(G34), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(G34), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n709), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G160), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n725), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n730), .B(new_n738), .C1(new_n739), .C2(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT100), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(KEYINPUT100), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n709), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n488), .A2(G140), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT96), .Z(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n753));
  INV_X1    g328(.A(G116), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(G2105), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n483), .B2(G128), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n750), .B1(new_n758), .B2(new_n725), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT97), .B(G2067), .Z(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n688), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n688), .ZN(new_n763));
  INV_X1    g338(.A(G1961), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n747), .A2(new_n748), .A3(new_n761), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n710), .A2(G35), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n710), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT29), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G2090), .ZN(new_n770));
  INV_X1    g345(.A(new_n605), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(new_n688), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G4), .B2(new_n688), .ZN(new_n773));
  INV_X1    g348(.A(G1348), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n688), .A2(G20), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT23), .Z(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G299), .B2(G16), .ZN(new_n779));
  INV_X1    g354(.A(G1956), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n632), .A2(new_n709), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT102), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n688), .A2(G21), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G168), .B2(new_n688), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT101), .B(G1966), .Z(new_n786));
  OAI21_X1  g361(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n781), .B(new_n787), .C1(new_n785), .C2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n745), .A2(new_n739), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT31), .B(G11), .Z(new_n790));
  INV_X1    g365(.A(G28), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(KEYINPUT30), .ZN(new_n792));
  AOI21_X1  g367(.A(G29), .B1(new_n791), .B2(KEYINPUT30), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n789), .B(new_n794), .C1(new_n727), .C2(new_n729), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n760), .B2(new_n759), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n710), .A2(G27), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G164), .B2(new_n710), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT103), .B(G2078), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT104), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n776), .A2(new_n788), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n688), .A2(G19), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT95), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n547), .B2(new_n688), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(G1341), .Z(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n769), .B2(G2090), .ZN(new_n807));
  OR4_X1    g382(.A1(new_n766), .A2(new_n775), .A3(new_n802), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n715), .A2(new_n808), .ZN(G311));
  INV_X1    g384(.A(G311), .ZN(G150));
  NAND2_X1  g385(.A1(new_n771), .A2(G559), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT38), .Z(new_n812));
  NAND3_X1  g387(.A1(new_n527), .A2(G67), .A3(new_n529), .ZN(new_n813));
  AND2_X1   g388(.A1(G80), .A2(G543), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT105), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n813), .A2(KEYINPUT105), .A3(new_n815), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n818), .A2(G651), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G93), .ZN(new_n821));
  INV_X1    g396(.A(G55), .ZN(new_n822));
  OAI22_X1  g397(.A1(new_n514), .A2(new_n821), .B1(new_n822), .B2(new_n503), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT106), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI221_X1 g400(.A(KEYINPUT106), .B1(new_n822), .B2(new_n503), .C1(new_n514), .C2(new_n821), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n820), .A2(new_n547), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n547), .B1(new_n820), .B2(new_n827), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n812), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n832));
  AOI21_X1  g407(.A(G860), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n832), .B2(new_n831), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n818), .A2(G651), .A3(new_n819), .ZN(new_n835));
  INV_X1    g410(.A(new_n827), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n837), .A2(new_n613), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n834), .A2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(new_n757), .B(new_n500), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n483), .A2(G130), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n458), .A2(G118), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G142), .B2(new_n488), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n841), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n708), .B(KEYINPUT107), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n623), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n723), .B(new_n736), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n847), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n632), .B(G160), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G162), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n852), .A2(new_n854), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n855), .A2(new_n856), .A3(G37), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g433(.A(new_n618), .B(new_n830), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n602), .A2(G299), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n597), .A2(new_n559), .A3(new_n557), .A4(new_n601), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT41), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n860), .A2(new_n864), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n859), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n862), .B(KEYINPUT108), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n859), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT109), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT109), .B1(new_n868), .B2(new_n870), .ZN(new_n873));
  XNOR2_X1  g448(.A(G303), .B(new_n567), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n591), .A2(G305), .A3(new_n592), .ZN(new_n876));
  AOI21_X1  g451(.A(G305), .B1(new_n591), .B2(new_n592), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(G290), .A2(new_n580), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n591), .A2(G305), .A3(new_n592), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n874), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT42), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n872), .B1(new_n873), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n871), .A2(KEYINPUT109), .A3(new_n883), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(G868), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(G868), .B2(new_n837), .ZN(G295));
  OAI21_X1  g464(.A(new_n888), .B1(G868), .B2(new_n837), .ZN(G331));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n878), .A2(new_n881), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n616), .B1(new_n835), .B2(new_n836), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n820), .A2(new_n547), .A3(new_n827), .ZN(new_n894));
  NOR2_X1   g469(.A1(G171), .A2(KEYINPUT111), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n828), .B2(new_n829), .ZN(new_n898));
  AOI21_X1  g473(.A(G286), .B1(KEYINPUT111), .B2(G171), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n900), .A2(new_n901), .A3(new_n862), .ZN(new_n902));
  INV_X1    g477(.A(new_n899), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n896), .B1(new_n893), .B2(new_n894), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n828), .A2(new_n829), .A3(new_n895), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n867), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n892), .A2(new_n902), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(G37), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n865), .A2(KEYINPUT113), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n863), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n862), .A2(KEYINPUT113), .A3(KEYINPUT41), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n906), .A2(new_n907), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT114), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n882), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n913), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n900), .B2(new_n901), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n906), .A2(new_n869), .A3(new_n907), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT114), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n916), .A2(KEYINPUT115), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT115), .B1(new_n916), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n910), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n906), .A2(new_n860), .A3(new_n861), .A4(new_n907), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n866), .B1(new_n900), .B2(new_n901), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n882), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT112), .B1(new_n927), .B2(G37), .ZN(new_n928));
  INV_X1    g503(.A(new_n909), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n892), .B1(new_n902), .B2(new_n908), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n931));
  INV_X1    g506(.A(G37), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n928), .A2(new_n929), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n891), .B1(new_n924), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n928), .A2(new_n929), .A3(new_n933), .ZN(new_n937));
  INV_X1    g512(.A(new_n934), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n910), .B(new_n934), .C1(new_n921), .C2(new_n922), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n939), .A2(new_n891), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n936), .A2(new_n941), .ZN(G397));
  INV_X1    g517(.A(KEYINPUT127), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT53), .ZN(new_n944));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  OAI211_X1 g520(.A(G138), .B(new_n458), .C1(new_n463), .C2(new_n467), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n499), .B1(new_n946), .B2(KEYINPUT4), .ZN(new_n947));
  OAI211_X1 g522(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n467), .ZN(new_n948));
  INV_X1    g523(.A(new_n492), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n945), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n468), .A2(new_n477), .A3(G40), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n944), .B1(new_n956), .B2(G2078), .ZN(new_n957));
  INV_X1    g532(.A(new_n955), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n951), .B2(KEYINPUT50), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n500), .A2(new_n960), .A3(new_n945), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n764), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n958), .A2(new_n944), .A3(G2078), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n954), .A3(new_n953), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n957), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  OR2_X1    g541(.A1(G171), .A2(KEYINPUT54), .ZN(new_n967));
  NAND2_X1  g542(.A1(G171), .A2(KEYINPUT54), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n964), .A2(new_n954), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n946), .A2(KEYINPUT4), .ZN(new_n972));
  INV_X1    g547(.A(new_n499), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(G1384), .B1(new_n974), .B2(new_n493), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT45), .B1(new_n951), .B2(KEYINPUT116), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n971), .A2(new_n979), .B1(new_n967), .B2(new_n968), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(new_n957), .A3(new_n963), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n970), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n983));
  INV_X1    g558(.A(G8), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n951), .A2(KEYINPUT50), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n985), .A2(new_n961), .A3(new_n955), .ZN(new_n986));
  INV_X1    g561(.A(G1966), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n986), .A2(new_n739), .B1(new_n956), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n984), .B1(new_n988), .B2(G168), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n959), .A2(new_n739), .A3(new_n961), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n958), .B1(new_n951), .B2(new_n952), .ZN(new_n991));
  AOI21_X1  g566(.A(G1966), .B1(new_n991), .B2(new_n954), .ZN(new_n992));
  OAI21_X1  g567(.A(G286), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n983), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n956), .A2(new_n987), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n995), .B(G168), .C1(G2084), .C2(new_n962), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n996), .A2(new_n983), .A3(G8), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n982), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n516), .A2(new_n517), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n505), .B1(new_n514), .B2(new_n515), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT55), .B(G8), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT119), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n1003));
  NAND4_X1  g578(.A1(G303), .A2(new_n1003), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT120), .ZN(new_n1006));
  INV_X1    g581(.A(new_n999), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1000), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n984), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1006), .B1(new_n1009), .B2(KEYINPUT55), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT120), .B(new_n1011), .C1(G166), .C2(new_n984), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1005), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT122), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n960), .B1(new_n500), .B2(new_n945), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n958), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT118), .B(G2090), .Z(new_n1018));
  NAND3_X1  g593(.A1(new_n985), .A2(KEYINPUT122), .A3(new_n955), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n961), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1971), .B1(new_n991), .B2(new_n954), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(KEYINPUT123), .B(new_n1014), .C1(new_n1023), .C2(new_n984), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n959), .A2(new_n1018), .A3(new_n961), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1013), .B(G8), .C1(new_n1021), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n574), .A2(new_n575), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(G651), .ZN(new_n1028));
  INV_X1    g603(.A(new_n579), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(G1981), .B1(new_n576), .B2(new_n579), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT49), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n984), .B1(new_n975), .B2(new_n955), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n500), .A2(new_n945), .A3(new_n955), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n565), .B(G1976), .C1(new_n566), .C2(new_n517), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(G8), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1035), .A2(new_n1036), .B1(KEYINPUT52), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n568), .A2(new_n1042), .A3(new_n570), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1041), .B1(new_n1045), .B2(new_n1039), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1037), .A2(G8), .A3(new_n1038), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1047), .A2(KEYINPUT121), .A3(new_n1044), .A4(new_n1043), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1026), .A2(new_n1040), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT123), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n984), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n1052), .B2(new_n1013), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1024), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n943), .B1(new_n998), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n970), .A2(new_n981), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n996), .A2(new_n993), .A3(G8), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT51), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n989), .A2(new_n983), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1052), .A2(new_n1051), .A3(new_n1013), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1026), .A2(new_n1049), .A3(new_n1040), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1060), .A2(KEYINPUT127), .A3(new_n1063), .A4(new_n1053), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1055), .A2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT56), .B(G2072), .Z(new_n1066));
  NOR2_X1   g641(.A1(new_n956), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1017), .A2(new_n961), .A3(new_n1019), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n780), .ZN(new_n1069));
  XOR2_X1   g644(.A(G299), .B(KEYINPUT57), .Z(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT125), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1070), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n959), .A2(KEYINPUT122), .B1(new_n960), .B2(new_n975), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1956), .B1(new_n1076), .B2(new_n1017), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1074), .B(new_n1075), .C1(new_n1077), .C2(new_n1067), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1071), .A2(new_n1073), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1077), .A2(new_n1075), .A3(new_n1067), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1072), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1037), .A2(G2067), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n962), .B2(new_n774), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n1085));
  INV_X1    g660(.A(new_n602), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n1088));
  INV_X1    g663(.A(G1996), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n953), .A2(new_n954), .A3(new_n1089), .A4(new_n955), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT58), .B(G1341), .Z(new_n1091));
  NAND2_X1  g666(.A1(new_n1037), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1088), .B1(new_n1093), .B2(new_n547), .ZN(new_n1094));
  AOI211_X1 g669(.A(KEYINPUT59), .B(new_n616), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1087), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1084), .A2(new_n602), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1348), .B1(new_n959), .B2(new_n961), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1086), .B1(new_n1098), .B2(new_n1083), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1085), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1079), .A2(new_n1082), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT126), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1071), .A2(new_n1099), .A3(new_n1078), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1081), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1102), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1103), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1065), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1049), .A2(new_n1040), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(new_n1026), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n571), .A2(new_n1042), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1031), .B1(new_n1035), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1111), .B1(new_n1036), .B2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n988), .A2(new_n984), .A3(G286), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1024), .A2(new_n1050), .A3(new_n1053), .A4(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT63), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1025), .A2(new_n1021), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1014), .B1(new_n1119), .B2(new_n984), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1115), .A2(new_n1120), .A3(KEYINPUT63), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n1062), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT124), .B(new_n1114), .C1(new_n1118), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1122), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1114), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1124), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT62), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n966), .A2(G171), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1128), .A2(KEYINPUT62), .ZN(new_n1132));
  OR3_X1    g707(.A1(new_n1131), .A2(new_n1054), .A3(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1109), .A2(new_n1123), .A3(new_n1127), .A4(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n977), .A2(new_n978), .A3(new_n955), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1089), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n723), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1135), .B(KEYINPUT117), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n757), .B(G2067), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n724), .A2(new_n1089), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1138), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n708), .A2(new_n712), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n708), .A2(new_n712), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1139), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n683), .A2(new_n686), .ZN(new_n1148));
  NAND2_X1  g723(.A1(G290), .A2(G1986), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1135), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1134), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1139), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n757), .A2(G2067), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1137), .B(KEYINPUT46), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1139), .B1(new_n723), .B2(new_n1140), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT47), .Z(new_n1160));
  INV_X1    g735(.A(new_n1147), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1148), .A2(new_n1135), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n1162), .B(KEYINPUT48), .Z(new_n1163));
  AOI211_X1 g738(.A(new_n1156), .B(new_n1160), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1152), .A2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g740(.A(G227), .ZN(new_n1167));
  OAI211_X1 g741(.A(new_n1167), .B(G319), .C1(new_n651), .C2(new_n652), .ZN(new_n1168));
  NOR3_X1   g742(.A1(new_n857), .A2(G229), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n939), .A2(new_n940), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1170), .ZN(G225));
  INV_X1    g745(.A(G225), .ZN(G308));
endmodule


