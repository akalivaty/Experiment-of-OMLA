//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND3_X1  g0012(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT64), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n212), .B1(new_n214), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT2), .B(G226), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XOR2_X1   g0034(.A(G50), .B(G58), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  INV_X1    g0040(.A(KEYINPUT67), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  INV_X1    g0042(.A(KEYINPUT3), .ZN(new_n243));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n245), .A2(new_n207), .A3(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT7), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g0049(.A1(new_n245), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n246), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n242), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G58), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(new_n242), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G58), .A2(G68), .ZN(new_n254));
  OAI21_X1  g0054(.A(G20), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G159), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(KEYINPUT16), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n241), .B1(new_n251), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT7), .B1(new_n262), .B2(new_n207), .ZN(new_n263));
  INV_X1    g0063(.A(new_n250), .ZN(new_n264));
  OAI21_X1  g0064(.A(G68), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n258), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT67), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT16), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n255), .A2(new_n257), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n269), .B1(new_n251), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G1), .A2(G13), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n276), .B(new_n269), .C1(new_n251), .C2(new_n270), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n268), .A2(new_n272), .A3(new_n275), .A4(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n279), .A2(new_n207), .A3(G1), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(new_n275), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n206), .A2(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n280), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n282), .A2(new_n286), .B1(new_n287), .B2(new_n284), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT65), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT65), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G1698), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n296), .A3(G223), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G226), .A2(G1698), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n262), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G87), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n244), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n292), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(new_n292), .C1(new_n299), .C2(new_n301), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(new_n291), .A3(G274), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n291), .A2(new_n306), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(new_n226), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(G190), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n303), .A2(new_n305), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n308), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n309), .A2(new_n226), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n302), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n278), .A2(new_n289), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(KEYINPUT17), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n278), .A2(new_n289), .A3(new_n319), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT71), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n278), .A2(KEYINPUT71), .A3(new_n289), .A4(new_n319), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n321), .B1(new_n326), .B2(KEYINPUT17), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n310), .A2(G179), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n303), .A2(new_n305), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n316), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT70), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT70), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n329), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n272), .A2(new_n277), .ZN(new_n337));
  INV_X1    g0137(.A(new_n275), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n259), .B2(new_n267), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n288), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n336), .A2(new_n340), .A3(KEYINPUT18), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT18), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n329), .A2(new_n334), .A3(new_n331), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n334), .B1(new_n329), .B2(new_n331), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n278), .A2(new_n289), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n342), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n327), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n349), .A2(KEYINPUT72), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n244), .A2(G20), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G150), .ZN(new_n353));
  INV_X1    g0153(.A(new_n256), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n283), .A2(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(G50), .A2(G58), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n207), .B1(new_n356), .B2(new_n242), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n275), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n281), .A2(G50), .A3(new_n285), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n358), .B(new_n359), .C1(G50), .C2(new_n287), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT9), .ZN(new_n361));
  INV_X1    g0161(.A(G226), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n308), .B1(new_n309), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n293), .B1(new_n245), .B2(new_n246), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(G223), .B1(new_n262), .B2(G77), .ZN(new_n365));
  INV_X1    g0165(.A(G222), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n294), .B(new_n296), .C1(new_n260), .C2(new_n261), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n363), .B1(new_n368), .B2(new_n292), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(new_n317), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(G190), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n361), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT10), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT10), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n361), .A2(new_n375), .A3(new_n371), .A4(new_n372), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G179), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n369), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n360), .B1(new_n369), .B2(G169), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n280), .A2(new_n242), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT12), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n351), .A2(G77), .B1(G20), .B2(new_n242), .ZN(new_n386));
  INV_X1    g0186(.A(G50), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n354), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(KEYINPUT11), .A3(new_n275), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n281), .A2(G68), .A3(new_n285), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT11), .B1(new_n388), .B2(new_n275), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n245), .A2(new_n246), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n226), .A2(new_n293), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n395), .A2(new_n396), .B1(G33), .B2(G97), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT65), .B(G1698), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n395), .A2(new_n398), .A3(G226), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n291), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G238), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n308), .B1(new_n309), .B2(new_n401), .ZN(new_n402));
  OR3_X1    g0202(.A1(new_n400), .A2(KEYINPUT13), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT13), .B1(new_n400), .B2(new_n402), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(G169), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n404), .A3(G179), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n405), .B2(G169), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n394), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n405), .A2(G200), .ZN(new_n412));
  INV_X1    g0212(.A(G190), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n393), .C1(new_n413), .C2(new_n405), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n401), .B1(new_n245), .B2(new_n246), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n262), .A2(G107), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n226), .C2(new_n367), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT66), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n291), .B1(new_n419), .B2(new_n420), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G244), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n308), .B1(new_n309), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(G179), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  INV_X1    g0229(.A(G77), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n429), .A2(new_n352), .B1(new_n207), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n283), .A2(new_n354), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n275), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n430), .B1(new_n206), .B2(G20), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n281), .A2(new_n434), .B1(new_n430), .B2(new_n280), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n425), .B1(new_n421), .B2(new_n422), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n437), .B2(G169), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n428), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n433), .B(new_n435), .C1(new_n427), .C2(new_n413), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n437), .A2(new_n317), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n383), .A2(new_n415), .A3(new_n440), .A4(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n349), .A2(KEYINPUT72), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n350), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT77), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT5), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(G41), .ZN(new_n449));
  INV_X1    g0249(.A(G41), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n206), .B(G45), .C1(new_n450), .C2(KEYINPUT5), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n452), .B1(KEYINPUT76), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(KEYINPUT76), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n291), .A2(G274), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n450), .A2(KEYINPUT5), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n292), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G257), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n364), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT4), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n367), .B2(new_n424), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n395), .A2(new_n398), .A3(KEYINPUT4), .A4(G244), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n292), .ZN(new_n469));
  AOI21_X1  g0269(.A(G169), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT73), .B(KEYINPUT6), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G97), .A2(G107), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n204), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT6), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(KEYINPUT73), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT73), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(KEYINPUT6), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n475), .A2(new_n477), .B1(new_n202), .B2(G107), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(G20), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n256), .A2(G77), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT74), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT74), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n479), .A2(new_n483), .A3(new_n480), .ZN(new_n484));
  OAI21_X1  g0284(.A(G107), .B1(new_n263), .B2(new_n264), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n482), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n275), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n287), .A2(G97), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n244), .A2(G1), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n280), .A2(new_n275), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n490), .B2(G97), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n470), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n468), .A2(KEYINPUT75), .A3(new_n292), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT75), .B1(new_n468), .B2(new_n292), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n458), .A2(new_n379), .A3(new_n462), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT78), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT75), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n469), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n468), .A2(KEYINPUT75), .A3(new_n292), .ZN(new_n500));
  AND4_X1   g0300(.A1(KEYINPUT78), .A2(new_n499), .A3(new_n496), .A4(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n492), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT79), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT79), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n492), .B(new_n504), .C1(new_n497), .C2(new_n501), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n495), .A2(new_n463), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G200), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n487), .A2(new_n491), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n469), .A2(new_n463), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G190), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n503), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n457), .A2(new_n454), .B1(new_n461), .B2(G264), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n395), .A2(G257), .A3(G1698), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G294), .ZN(new_n515));
  INV_X1    g0315(.A(G250), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n515), .C1(new_n516), .C2(new_n367), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n292), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n330), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n513), .A2(new_n518), .A3(G179), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(KEYINPUT86), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT86), .ZN(new_n523));
  INV_X1    g0323(.A(new_n521), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n519), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n207), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(KEYINPUT85), .B2(KEYINPUT22), .ZN(new_n527));
  NOR2_X1   g0327(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n395), .A2(new_n207), .A3(G87), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT23), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n207), .B2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n535));
  INV_X1    g0335(.A(G116), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n244), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n534), .A2(new_n535), .B1(new_n537), .B2(new_n207), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n532), .B1(new_n531), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n275), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT25), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n287), .A2(new_n542), .A3(G107), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n542), .B1(new_n287), .B2(G107), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n544), .A2(new_n545), .B1(G107), .B2(new_n490), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n522), .A2(new_n525), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n513), .A2(new_n518), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n317), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(G190), .B2(new_n549), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n541), .A3(new_n546), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT84), .ZN(new_n554));
  INV_X1    g0354(.A(G45), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n516), .B1(new_n555), .B2(G1), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n206), .A2(G45), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n556), .B(new_n291), .C1(G274), .C2(new_n557), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n558), .B(KEYINPUT80), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n537), .B1(new_n416), .B2(new_n398), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n364), .A2(G244), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n291), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(G200), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n395), .A2(new_n207), .A3(G68), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n352), .B2(new_n202), .ZN(new_n567));
  NAND3_X1  g0367(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n207), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT82), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n300), .A2(new_n202), .A3(new_n203), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n569), .A2(KEYINPUT82), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n565), .B(new_n567), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n275), .B1(new_n280), .B2(new_n429), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n490), .A2(G87), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n554), .B1(new_n564), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n559), .A2(new_n562), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G190), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n563), .A2(new_n575), .A3(KEYINPUT84), .A4(new_n576), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n379), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT81), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n330), .B1(new_n559), .B2(new_n562), .ZN(new_n586));
  INV_X1    g0386(.A(new_n490), .ZN(new_n587));
  XOR2_X1   g0387(.A(new_n429), .B(KEYINPUT83), .Z(new_n588));
  OAI21_X1  g0388(.A(new_n575), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n579), .A2(KEYINPUT81), .A3(new_n379), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n585), .A2(new_n586), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G283), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n593), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n536), .A2(G20), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n275), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n287), .A2(G116), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n490), .B2(G116), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n395), .A2(new_n398), .A3(G257), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n395), .A2(G264), .A3(G1698), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n262), .A2(G303), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n292), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n461), .A2(G270), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n458), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n601), .B1(new_n608), .B2(G200), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n413), .B2(new_n608), .ZN(new_n610));
  INV_X1    g0410(.A(new_n608), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(G179), .A3(new_n601), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT21), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n330), .B1(new_n598), .B2(new_n600), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n608), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n614), .A2(new_n608), .A3(new_n613), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n610), .B(new_n612), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n553), .A2(new_n592), .A3(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n446), .A2(new_n512), .A3(new_n618), .ZN(G372));
  OAI21_X1  g0419(.A(KEYINPUT18), .B1(new_n336), .B2(new_n340), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n345), .A2(new_n342), .A3(new_n346), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n439), .A2(new_n414), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n411), .ZN(new_n624));
  XOR2_X1   g0424(.A(new_n624), .B(KEYINPUT91), .Z(new_n625));
  AOI21_X1  g0425(.A(new_n622), .B1(new_n625), .B2(new_n327), .ZN(new_n626));
  OAI22_X1  g0426(.A1(new_n626), .A2(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT88), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n577), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n575), .A2(KEYINPUT88), .A3(new_n576), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n559), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT87), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n562), .A2(new_n635), .ZN(new_n636));
  AOI211_X1 g0436(.A(KEYINPUT87), .B(new_n291), .C1(new_n560), .C2(new_n561), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G200), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n633), .A2(new_n580), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n638), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n589), .B(new_n583), .C1(new_n641), .C2(G169), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n629), .B1(new_n643), .B2(new_n502), .ZN(new_n644));
  INV_X1    g0444(.A(new_n592), .ZN(new_n645));
  INV_X1    g0445(.A(new_n505), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n495), .A2(KEYINPUT78), .A3(new_n496), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n499), .A2(new_n500), .A3(new_n496), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT78), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n504), .B1(new_n651), .B2(new_n492), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n645), .B1(new_n646), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g0453(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n644), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n640), .A2(new_n552), .A3(new_n642), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n612), .B1(new_n616), .B2(new_n615), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g0459(.A(KEYINPUT89), .B(new_n612), .C1(new_n616), .C2(new_n615), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n547), .B1(new_n519), .B2(new_n524), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n656), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n512), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n655), .A2(new_n642), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n446), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n628), .A2(new_n666), .ZN(G369));
  INV_X1    g0467(.A(new_n657), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n601), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n668), .A2(new_n610), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n661), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  INV_X1    g0478(.A(new_n553), .ZN(new_n679));
  INV_X1    g0479(.A(new_n547), .ZN(new_n680));
  INV_X1    g0480(.A(new_n674), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n548), .A2(new_n681), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n668), .A2(new_n674), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n662), .A2(new_n674), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(KEYINPUT92), .ZN(new_n692));
  INV_X1    g0492(.A(new_n210), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(G41), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n210), .A2(KEYINPUT92), .A3(new_n450), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n571), .A2(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n215), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT29), .B1(new_n665), .B2(new_n681), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n592), .B1(new_n503), .B2(new_n505), .ZN(new_n702));
  INV_X1    g0502(.A(new_n654), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT93), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n653), .A2(new_n705), .A3(new_n654), .ZN(new_n706));
  INV_X1    g0506(.A(new_n643), .ZN(new_n707));
  INV_X1    g0507(.A(new_n502), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(KEYINPUT26), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n704), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n642), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n656), .B1(new_n668), .B2(new_n548), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(new_n512), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n674), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n701), .B1(KEYINPUT29), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n512), .A2(new_n618), .A3(new_n681), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n579), .A2(new_n607), .A3(new_n606), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(new_n509), .A3(new_n524), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n718), .A2(new_n509), .A3(new_n524), .A4(KEYINPUT30), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n549), .A2(new_n608), .A3(new_n379), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n506), .A2(new_n638), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n725), .B2(new_n674), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n716), .B1(new_n717), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n715), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n700), .B1(new_n730), .B2(G1), .ZN(G364));
  INV_X1    g0531(.A(new_n696), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n279), .A2(G20), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G45), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n206), .B1(new_n734), .B2(KEYINPUT94), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(KEYINPUT94), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n677), .B2(G330), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G330), .B2(new_n677), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n274), .B1(G20), .B2(new_n330), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n210), .A2(new_n262), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n236), .A2(G45), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT95), .ZN(new_n747));
  INV_X1    g0547(.A(new_n215), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n745), .B(new_n747), .C1(new_n555), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n210), .A2(new_n395), .ZN(new_n750));
  INV_X1    g0550(.A(G355), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n750), .A2(new_n751), .B1(G116), .B2(new_n210), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n744), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n207), .A2(new_n379), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G190), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n207), .A2(G179), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n755), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G311), .A2(new_n757), .B1(new_n760), .B2(G329), .ZN(new_n761));
  INV_X1    g0561(.A(G322), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n754), .A2(G190), .A3(new_n317), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n761), .B(new_n262), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n413), .A2(G179), .A3(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n207), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n767), .A2(G294), .B1(new_n769), .B2(G303), .ZN(new_n770));
  INV_X1    g0570(.A(G283), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n758), .A2(new_n413), .A3(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n754), .A2(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT33), .B(G317), .Z(new_n776));
  OAI221_X1 g0576(.A(new_n770), .B1(new_n771), .B2(new_n772), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n773), .A2(new_n413), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT96), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n764), .B(new_n777), .C1(G326), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n769), .A2(G87), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n782), .B1(new_n202), .B2(new_n766), .C1(new_n203), .C2(new_n772), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n760), .A2(G159), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  INV_X1    g0585(.A(new_n778), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n387), .A2(new_n786), .B1(new_n775), .B2(new_n242), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n395), .B1(new_n756), .B2(new_n430), .C1(new_n252), .C2(new_n763), .ZN(new_n788));
  NOR4_X1   g0588(.A1(new_n783), .A2(new_n785), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n743), .B1(new_n781), .B2(new_n789), .ZN(new_n790));
  AND3_X1   g0590(.A1(new_n753), .A2(new_n737), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n742), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n677), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n739), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  NOR3_X1   g0595(.A1(new_n428), .A2(new_n438), .A3(new_n674), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n436), .A2(new_n674), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n441), .B2(new_n442), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(new_n798), .B2(new_n440), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n665), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n801), .B2(new_n674), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n665), .A2(new_n681), .A3(new_n799), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n729), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n737), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n802), .A2(new_n729), .A3(new_n803), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n774), .A2(G150), .B1(new_n778), .B2(G137), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT98), .Z(new_n809));
  INV_X1    g0609(.A(new_n763), .ZN(new_n810));
  XNOR2_X1  g0610(.A(KEYINPUT99), .B(G143), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n810), .A2(new_n812), .B1(new_n757), .B2(G159), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n809), .A2(KEYINPUT34), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n772), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G68), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n262), .B1(new_n760), .B2(G132), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n767), .A2(G58), .B1(new_n769), .B2(G50), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n814), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(KEYINPUT34), .B1(new_n809), .B2(new_n813), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G303), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n771), .A2(new_n775), .B1(new_n786), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G87), .B2(new_n815), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n395), .B1(new_n760), .B2(G311), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n810), .A2(G294), .B1(new_n757), .B2(G116), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n767), .A2(G97), .B1(new_n769), .B2(G107), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT97), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n743), .B1(new_n821), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n743), .A2(new_n740), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n736), .B(new_n732), .C1(new_n430), .C2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n830), .B(new_n832), .C1(new_n799), .C2(new_n741), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n807), .A2(new_n833), .ZN(G384));
  NOR2_X1   g0634(.A1(new_n733), .A2(new_n206), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT17), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n324), .B2(new_n325), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n622), .A2(new_n837), .A3(new_n321), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n288), .B1(new_n339), .B2(new_n271), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n672), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT100), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT100), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n349), .A2(new_n843), .A3(new_n840), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n839), .B1(new_n336), .B2(new_n672), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT37), .B1(new_n326), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n672), .B1(new_n278), .B2(new_n289), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(KEYINPUT37), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n346), .A2(new_n335), .A3(new_n333), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n849), .A2(new_n850), .A3(new_n324), .A4(new_n325), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  INV_X1    g0654(.A(new_n672), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n346), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n850), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n326), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n320), .A2(new_n848), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n854), .B1(new_n859), .B2(new_n850), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT101), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n850), .A2(new_n322), .A3(new_n856), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT101), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(new_n851), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n861), .B(new_n865), .C1(new_n838), .C2(new_n856), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n866), .A2(KEYINPUT102), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT102), .B1(new_n866), .B2(new_n867), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n853), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n838), .A2(KEYINPUT100), .A3(new_n841), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n843), .B1(new_n349), .B2(new_n840), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n852), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n867), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(KEYINPUT39), .A3(new_n853), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n411), .A2(new_n674), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n872), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n876), .A2(new_n853), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n394), .A2(new_n674), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n411), .A2(new_n414), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n411), .B2(new_n414), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n796), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n885), .B1(new_n803), .B2(new_n886), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n881), .A2(new_n887), .B1(new_n622), .B2(new_n672), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n627), .B1(new_n715), .B2(new_n446), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n889), .B(new_n890), .Z(new_n891));
  NAND2_X1  g0691(.A1(new_n725), .A2(new_n674), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT103), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT31), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n725), .A2(new_n893), .A3(new_n894), .A4(new_n674), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n717), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n799), .B1(new_n883), .B2(new_n884), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n899), .A2(KEYINPUT104), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT104), .B1(new_n899), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT40), .B1(new_n881), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n901), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n870), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n446), .A2(new_n899), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n716), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n835), .B1(new_n891), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n891), .B2(new_n911), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n214), .A2(new_n536), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n473), .A2(new_n478), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT35), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n916), .B2(new_n915), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT36), .Z(new_n919));
  NOR3_X1   g0719(.A1(new_n253), .A2(new_n215), .A3(new_n430), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n242), .A2(G50), .ZN(new_n921));
  OAI211_X1 g0721(.A(G1), .B(new_n279), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n913), .A2(new_n919), .A3(new_n922), .ZN(G367));
  OAI21_X1  g0723(.A(new_n512), .B1(new_n508), .B2(new_n681), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n708), .A2(new_n674), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n687), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT42), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n503), .B(new_n505), .C1(new_n927), .C2(new_n548), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n681), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n631), .A2(new_n632), .A3(new_n674), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n707), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n642), .A2(new_n933), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n932), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n929), .A2(new_n938), .A3(new_n937), .A4(new_n931), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n941), .A2(new_n684), .A3(new_n926), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n685), .B2(new_n927), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n696), .B(KEYINPUT41), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT105), .B1(new_n927), .B2(new_n689), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT105), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n926), .A2(new_n948), .A3(new_n690), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT45), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n947), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n926), .A2(new_n690), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT44), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n684), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n682), .A2(new_n683), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n687), .B1(new_n958), .B2(new_n686), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT106), .B1(new_n677), .B2(G330), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n959), .B(new_n960), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n730), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n952), .A2(new_n685), .A3(new_n953), .A4(new_n955), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n957), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n946), .B1(new_n965), .B2(new_n730), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n736), .B(KEYINPUT107), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n943), .B(new_n945), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n744), .B1(new_n210), .B2(new_n429), .C1(new_n232), .C2(new_n745), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT108), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n971), .A2(new_n737), .A3(new_n972), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n780), .A2(G311), .B1(G303), .B2(new_n810), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT109), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(KEYINPUT109), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n769), .A2(G116), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT46), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT110), .ZN(new_n980));
  INV_X1    g0780(.A(G317), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n262), .B1(new_n759), .B2(new_n981), .C1(new_n771), .C2(new_n756), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G107), .A2(new_n767), .B1(new_n774), .B2(G294), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n202), .B2(new_n772), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(new_n978), .C2(new_n977), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n975), .A2(new_n976), .A3(new_n980), .A4(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n766), .A2(new_n242), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G150), .B2(new_n810), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT111), .ZN(new_n989));
  INV_X1    g0789(.A(G137), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n395), .B1(new_n759), .B2(new_n990), .C1(new_n387), .C2(new_n756), .ZN(new_n991));
  INV_X1    g0791(.A(G159), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n775), .A2(new_n992), .B1(new_n772), .B2(new_n430), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(G58), .C2(new_n769), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n779), .B2(new_n811), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n986), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT47), .Z(new_n997));
  INV_X1    g0797(.A(new_n743), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n973), .B1(new_n792), .B2(new_n936), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n968), .A2(new_n999), .ZN(G387));
  NOR2_X1   g0800(.A1(new_n963), .A2(new_n696), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n730), .B2(new_n961), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n750), .A2(new_n697), .B1(G107), .B2(new_n210), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n229), .A2(new_n555), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n697), .ZN(new_n1005));
  AOI211_X1 g0805(.A(G45), .B(new_n1005), .C1(G68), .C2(G77), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n283), .A2(G50), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n745), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1003), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n744), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n737), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n763), .A2(new_n387), .B1(new_n756), .B2(new_n242), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n262), .B(new_n1013), .C1(G150), .C2(new_n760), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n778), .A2(G159), .B1(new_n815), .B2(G97), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n588), .A2(new_n766), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n774), .A2(new_n284), .B1(new_n769), .B2(G77), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n395), .B1(new_n760), .B2(G326), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n810), .A2(G317), .B1(new_n757), .B2(G303), .ZN(new_n1020));
  INV_X1    g0820(.A(G311), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n775), .C1(new_n779), .C2(new_n762), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT112), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT48), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(KEYINPUT48), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n767), .A2(G283), .B1(new_n769), .B2(G294), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1019), .B1(new_n536), .B2(new_n772), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1028), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(KEYINPUT49), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1018), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1012), .B1(new_n1033), .B2(new_n743), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n682), .A2(new_n683), .A3(new_n742), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1034), .A2(new_n1035), .B1(new_n961), .B2(new_n967), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1002), .A2(new_n1036), .ZN(G393));
  OAI221_X1 g0837(.A(new_n744), .B1(new_n202), .B2(new_n210), .C1(new_n239), .C2(new_n745), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n737), .A2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G317), .A2(new_n778), .B1(new_n810), .B2(G311), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT52), .ZN(new_n1041));
  INV_X1    g0841(.A(G294), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n262), .B1(new_n759), .B2(new_n762), .C1(new_n1042), .C2(new_n756), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n766), .A2(new_n536), .B1(new_n772), .B2(new_n203), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n775), .A2(new_n822), .B1(new_n771), .B2(new_n768), .ZN(new_n1045));
  NOR4_X1   g0845(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n786), .A2(new_n353), .B1(new_n992), .B2(new_n763), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT51), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n766), .A2(new_n430), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G68), .B2(new_n769), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n395), .B1(new_n759), .B2(new_n811), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n284), .B2(new_n757), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n774), .A2(G50), .B1(new_n815), .B2(G87), .ZN(new_n1053));
  AND3_X1   g0853(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1046), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1039), .B1(new_n998), .B2(new_n1055), .C1(new_n926), .C2(new_n792), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n957), .A2(new_n964), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n967), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n965), .A2(new_n732), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n962), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(G390));
  NAND2_X1  g0863(.A1(new_n899), .A2(G330), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1064), .A2(new_n900), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n887), .A2(new_n879), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n872), .B2(new_n877), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n710), .A2(new_n713), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n798), .A2(new_n440), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n681), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n885), .B1(new_n1070), .B2(new_n886), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n852), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n867), .B(new_n1072), .C1(new_n842), .C2(new_n844), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT102), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n865), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n856), .B1(new_n327), .B2(new_n348), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n864), .B1(new_n863), .B2(new_n851), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1074), .B1(new_n1078), .B2(KEYINPUT38), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n866), .A2(KEYINPUT102), .A3(new_n867), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1073), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1071), .A2(new_n1081), .A3(new_n879), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1065), .B1(new_n1067), .B2(new_n1082), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n887), .A2(new_n879), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT39), .B1(new_n1085), .B2(new_n853), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n877), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n796), .B1(new_n714), .B2(new_n1069), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n870), .B(new_n878), .C1(new_n1089), .C2(new_n885), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n716), .B(new_n800), .C1(new_n717), .C2(new_n728), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n885), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1088), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n899), .A2(G330), .A3(new_n799), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n885), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1070), .A2(new_n1093), .A3(new_n1096), .A4(new_n886), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1091), .A2(new_n1092), .B1(new_n1064), .B2(new_n900), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n803), .A2(new_n886), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n716), .B1(new_n717), .B2(new_n898), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n446), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n890), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1083), .A2(new_n1094), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(KEYINPUT113), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT113), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1083), .A2(new_n1094), .A3(new_n1108), .A4(new_n1105), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1083), .A2(new_n1094), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n696), .B1(new_n1111), .B2(new_n1104), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1111), .A2(new_n1058), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n740), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n831), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n737), .B1(new_n284), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n786), .A2(new_n1118), .B1(new_n772), .B2(new_n387), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G159), .B2(new_n767), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n768), .A2(new_n353), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT53), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n760), .A2(G125), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n262), .B1(new_n810), .B2(G132), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT54), .B(G143), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n774), .A2(G137), .B1(new_n757), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT114), .Z(new_n1129));
  AOI21_X1  g0929(.A(new_n1049), .B1(G283), .B2(new_n778), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n203), .B2(new_n775), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n756), .A2(new_n202), .B1(new_n759), .B2(new_n1042), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n395), .B(new_n1132), .C1(G116), .C2(new_n810), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(new_n782), .A3(new_n816), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1125), .A2(new_n1129), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1117), .B1(new_n1135), .B2(new_n743), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1114), .B1(new_n1115), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1113), .A2(new_n1137), .ZN(G378));
  AOI21_X1  g0938(.A(new_n716), .B1(new_n870), .B2(new_n907), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT121), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n881), .A2(new_n904), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(new_n1140), .C1(new_n1141), .C2(KEYINPUT40), .ZN(new_n1142));
  OAI21_X1  g0942(.A(G330), .B1(new_n1081), .B2(new_n906), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT121), .B1(new_n1143), .B2(new_n905), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n360), .A2(new_n855), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n383), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n383), .A2(new_n1145), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1146), .A2(new_n1147), .A3(KEYINPUT119), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT119), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1142), .A2(new_n1144), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n889), .ZN(new_n1157));
  OAI211_X1 g0957(.A(KEYINPUT121), .B(new_n1154), .C1(new_n1143), .C2(new_n905), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1157), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OR2_X1    g0961(.A1(KEYINPUT117), .A2(G124), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(KEYINPUT117), .A2(G124), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n760), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(G33), .A2(G41), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n992), .C2(new_n772), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G150), .A2(new_n767), .B1(new_n778), .B2(G125), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT115), .Z(new_n1168));
  OAI22_X1  g0968(.A1(new_n763), .A2(new_n1118), .B1(new_n756), .B2(new_n990), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G132), .B2(new_n774), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(new_n768), .C2(new_n1126), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT116), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1166), .B1(new_n1172), .B2(KEYINPUT59), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(KEYINPUT59), .B2(new_n1172), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n395), .A2(G41), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n771), .B2(new_n759), .C1(new_n203), .C2(new_n763), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n987), .B(new_n1176), .C1(G77), .C2(new_n769), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n775), .A2(new_n202), .B1(new_n772), .B2(new_n252), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G116), .B2(new_n778), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(new_n588), .C2(new_n756), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT58), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n387), .B1(G33), .B2(G41), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1174), .B(new_n1181), .C1(new_n1175), .C2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n998), .B1(new_n1183), .B2(KEYINPUT118), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(KEYINPUT118), .B2(new_n1183), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n736), .B(new_n732), .C1(new_n387), .C2(new_n831), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n1154), .C2(new_n741), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT120), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(KEYINPUT120), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1161), .A2(new_n967), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n701), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n446), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(new_n628), .A3(new_n1103), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1110), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1161), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n889), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(KEYINPUT57), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1194), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n732), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1190), .B1(new_n1197), .B2(new_n1203), .ZN(G375));
  AND3_X1   g1004(.A1(new_n729), .A2(new_n799), .A3(new_n1092), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1092), .B1(new_n1102), .B2(new_n799), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1207), .A2(new_n1089), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1194), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n946), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1104), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n737), .B1(G68), .B2(new_n1116), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n763), .A2(new_n990), .B1(new_n756), .B2(new_n353), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n262), .B(new_n1213), .C1(G128), .C2(new_n760), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n769), .A2(G159), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G132), .A2(new_n778), .B1(new_n774), .B2(new_n1127), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n767), .A2(G50), .B1(new_n815), .B2(G58), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1016), .B1(new_n771), .B2(new_n763), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT122), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n786), .A2(new_n1042), .B1(new_n772), .B2(new_n430), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n775), .A2(new_n536), .B1(new_n202), .B2(new_n768), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n262), .B1(new_n759), .B2(new_n822), .C1(new_n203), .C2(new_n756), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1218), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1212), .B1(new_n1225), .B2(new_n743), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1092), .B2(new_n741), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1208), .B2(new_n1058), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1211), .A2(new_n1229), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT123), .Z(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(G381));
  NAND3_X1  g1032(.A1(new_n1002), .A2(new_n794), .A3(new_n1036), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1233), .A2(G384), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT124), .Z(new_n1235));
  NAND3_X1  g1035(.A1(new_n968), .A2(new_n1062), .A3(new_n999), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1235), .A2(G381), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(G378), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1239), .B1(new_n1240), .B2(new_n1058), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT57), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1159), .A2(new_n1160), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n696), .B1(new_n1196), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1202), .B2(new_n1240), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1241), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1237), .A2(new_n1238), .A3(new_n1246), .ZN(G407));
  NAND2_X1  g1047(.A1(new_n673), .A2(G213), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1246), .A2(new_n1238), .A3(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(G407), .A2(G213), .A3(new_n1250), .ZN(G409));
  AOI21_X1  g1051(.A(new_n1062), .B1(new_n968), .B2(new_n999), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G393), .A2(G396), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1233), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1236), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1255), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1236), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(new_n1252), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT125), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1194), .A2(new_n1208), .A3(KEYINPUT60), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n1104), .A3(new_n732), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT60), .B1(new_n1194), .B2(new_n1208), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1261), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n696), .B1(new_n1195), .B2(new_n1101), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1209), .A2(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1266), .A2(new_n1268), .A3(KEYINPUT125), .A4(new_n1262), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1265), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1229), .ZN(new_n1271));
  INV_X1    g1071(.A(G384), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(G384), .A3(new_n1229), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(KEYINPUT126), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT126), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G384), .B1(new_n1270), .B2(new_n1229), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1272), .B(new_n1228), .C1(new_n1265), .C2(new_n1269), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1249), .A2(G2897), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1275), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(G2897), .A3(new_n1249), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1196), .A2(new_n1210), .A3(new_n1161), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G378), .B1(new_n1285), .B2(new_n1190), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(new_n1246), .B2(G378), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1284), .B1(new_n1287), .B2(new_n1249), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G378), .B(new_n1190), .C1(new_n1197), .C2(new_n1203), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1202), .A2(new_n1240), .A3(new_n946), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1238), .B1(new_n1291), .B2(new_n1241), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1248), .A4(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1288), .A2(new_n1289), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1249), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1294), .B1(new_n1298), .B2(new_n1295), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1260), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1256), .A2(new_n1259), .A3(new_n1289), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1301), .B(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1298), .A2(new_n1295), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1298), .A2(KEYINPUT63), .A3(new_n1295), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1303), .A2(new_n1306), .A3(new_n1288), .A4(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1300), .A2(new_n1308), .ZN(G405));
  NOR2_X1   g1109(.A1(new_n1246), .A2(G378), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1290), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1282), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1295), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1313), .A2(new_n1314), .A3(new_n1260), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1260), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(G402));
endmodule


