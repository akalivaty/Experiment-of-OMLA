

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603;

  XNOR2_X1 U326 ( .A(n373), .B(n372), .ZN(n391) );
  XNOR2_X1 U327 ( .A(n362), .B(n412), .ZN(n363) );
  XOR2_X1 U328 ( .A(n412), .B(n411), .Z(n414) );
  XNOR2_X1 U329 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U330 ( .A(n490), .B(n489), .ZN(n519) );
  XNOR2_X1 U331 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n372) );
  XNOR2_X1 U332 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n397) );
  XNOR2_X1 U333 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U334 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U335 ( .A(n431), .B(n354), .ZN(n357) );
  XNOR2_X1 U336 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n394) );
  XOR2_X1 U337 ( .A(G36GAT), .B(G190GAT), .Z(n411) );
  XNOR2_X1 U338 ( .A(n361), .B(n360), .ZN(n412) );
  XNOR2_X1 U339 ( .A(n395), .B(n394), .ZN(n403) );
  INV_X1 U340 ( .A(KEYINPUT93), .ZN(n416) );
  INV_X1 U341 ( .A(KEYINPUT96), .ZN(n477) );
  INV_X1 U342 ( .A(KEYINPUT54), .ZN(n426) );
  XNOR2_X1 U343 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U344 ( .A(n364), .B(n363), .ZN(n367) );
  XNOR2_X1 U345 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U346 ( .A(n305), .B(n304), .ZN(n311) );
  INV_X1 U347 ( .A(G183GAT), .ZN(n495) );
  INV_X1 U348 ( .A(G43GAT), .ZN(n491) );
  XNOR2_X1 U349 ( .A(n424), .B(n443), .ZN(n542) );
  XNOR2_X1 U350 ( .A(n466), .B(KEYINPUT58), .ZN(n467) );
  XNOR2_X1 U351 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U352 ( .A(n468), .B(n467), .ZN(G1351GAT) );
  XNOR2_X1 U353 ( .A(n494), .B(n493), .ZN(G1330GAT) );
  XOR2_X1 U354 ( .A(G99GAT), .B(G85GAT), .Z(n365) );
  XOR2_X1 U355 ( .A(KEYINPUT79), .B(n365), .Z(n295) );
  XOR2_X1 U356 ( .A(G134GAT), .B(KEYINPUT78), .Z(n318) );
  XNOR2_X1 U357 ( .A(G218GAT), .B(n318), .ZN(n294) );
  XNOR2_X1 U358 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U359 ( .A(G92GAT), .B(n411), .Z(n297) );
  NAND2_X1 U360 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U361 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U362 ( .A(n299), .B(n298), .Z(n305) );
  XOR2_X1 U363 ( .A(G50GAT), .B(G162GAT), .Z(n437) );
  XNOR2_X1 U364 ( .A(G106GAT), .B(n437), .ZN(n303) );
  XOR2_X1 U365 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n301) );
  XNOR2_X1 U366 ( .A(KEYINPUT9), .B(KEYINPUT66), .ZN(n300) );
  XNOR2_X1 U367 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U368 ( .A(G43GAT), .B(KEYINPUT71), .ZN(n306) );
  XNOR2_X1 U369 ( .A(n306), .B(G29GAT), .ZN(n307) );
  XOR2_X1 U370 ( .A(n307), .B(KEYINPUT7), .Z(n309) );
  XNOR2_X1 U371 ( .A(KEYINPUT70), .B(KEYINPUT8), .ZN(n308) );
  XNOR2_X1 U372 ( .A(n309), .B(n308), .ZN(n343) );
  INV_X1 U373 ( .A(n343), .ZN(n310) );
  XOR2_X1 U374 ( .A(n311), .B(n310), .Z(n577) );
  XOR2_X1 U375 ( .A(G85GAT), .B(G162GAT), .Z(n313) );
  XNOR2_X1 U376 ( .A(G127GAT), .B(G148GAT), .ZN(n312) );
  XNOR2_X1 U377 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U378 ( .A(n314), .B(G120GAT), .Z(n316) );
  XOR2_X1 U379 ( .A(G113GAT), .B(KEYINPUT0), .Z(n456) );
  XNOR2_X1 U380 ( .A(G29GAT), .B(n456), .ZN(n315) );
  XNOR2_X1 U381 ( .A(n316), .B(n315), .ZN(n322) );
  XNOR2_X1 U382 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n317) );
  XNOR2_X1 U383 ( .A(n317), .B(KEYINPUT2), .ZN(n436) );
  XOR2_X1 U384 ( .A(n318), .B(n436), .Z(n320) );
  NAND2_X1 U385 ( .A1(G225GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U386 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U387 ( .A(n322), .B(n321), .Z(n330) );
  XOR2_X1 U388 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n324) );
  XNOR2_X1 U389 ( .A(G1GAT), .B(G155GAT), .ZN(n323) );
  XNOR2_X1 U390 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U391 ( .A(G57GAT), .B(KEYINPUT4), .Z(n326) );
  XNOR2_X1 U392 ( .A(KEYINPUT6), .B(KEYINPUT92), .ZN(n325) );
  XNOR2_X1 U393 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U394 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n330), .B(n329), .ZN(n540) );
  XOR2_X1 U396 ( .A(G15GAT), .B(G113GAT), .Z(n332) );
  XOR2_X1 U397 ( .A(G1GAT), .B(KEYINPUT72), .Z(n375) );
  XOR2_X1 U398 ( .A(G169GAT), .B(G8GAT), .Z(n415) );
  XNOR2_X1 U399 ( .A(n375), .B(n415), .ZN(n331) );
  XNOR2_X1 U400 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U401 ( .A(n333), .B(G50GAT), .Z(n338) );
  XOR2_X1 U402 ( .A(KEYINPUT30), .B(G22GAT), .Z(n335) );
  XNOR2_X1 U403 ( .A(G197GAT), .B(G141GAT), .ZN(n334) );
  XNOR2_X1 U404 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U405 ( .A(n336), .B(G36GAT), .ZN(n337) );
  XNOR2_X1 U406 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U407 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n340) );
  NAND2_X1 U408 ( .A1(G229GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U409 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U410 ( .A(n342), .B(n341), .Z(n345) );
  XNOR2_X1 U411 ( .A(n343), .B(KEYINPUT68), .ZN(n344) );
  XNOR2_X1 U412 ( .A(n345), .B(n344), .ZN(n587) );
  INV_X1 U413 ( .A(G148GAT), .ZN(n346) );
  NAND2_X1 U414 ( .A1(n346), .A2(G78GAT), .ZN(n349) );
  INV_X1 U415 ( .A(G78GAT), .ZN(n347) );
  NAND2_X1 U416 ( .A1(n347), .A2(G148GAT), .ZN(n348) );
  NAND2_X1 U417 ( .A1(n349), .A2(n348), .ZN(n351) );
  XNOR2_X1 U418 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n431) );
  NAND2_X1 U420 ( .A1(G230GAT), .A2(G233GAT), .ZN(n353) );
  INV_X1 U421 ( .A(KEYINPUT31), .ZN(n352) );
  INV_X1 U422 ( .A(n357), .ZN(n355) );
  NAND2_X1 U423 ( .A1(n355), .A2(KEYINPUT74), .ZN(n359) );
  INV_X1 U424 ( .A(KEYINPUT74), .ZN(n356) );
  NAND2_X1 U425 ( .A1(n357), .A2(n356), .ZN(n358) );
  NAND2_X1 U426 ( .A1(n359), .A2(n358), .ZN(n364) );
  XOR2_X1 U427 ( .A(G57GAT), .B(KEYINPUT13), .Z(n374) );
  XNOR2_X1 U428 ( .A(n374), .B(KEYINPUT76), .ZN(n362) );
  XOR2_X1 U429 ( .A(G64GAT), .B(G92GAT), .Z(n361) );
  XNOR2_X1 U430 ( .A(G176GAT), .B(G204GAT), .ZN(n360) );
  XOR2_X1 U431 ( .A(G120GAT), .B(G71GAT), .Z(n452) );
  XOR2_X1 U432 ( .A(n452), .B(n365), .Z(n366) );
  XNOR2_X1 U433 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U434 ( .A(KEYINPUT77), .B(KEYINPUT73), .Z(n369) );
  XNOR2_X1 U435 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n368) );
  XOR2_X1 U436 ( .A(n369), .B(n368), .Z(n370) );
  XNOR2_X1 U437 ( .A(n371), .B(n370), .ZN(n592) );
  XOR2_X1 U438 ( .A(KEYINPUT41), .B(n592), .Z(n522) );
  NOR2_X1 U439 ( .A1(n587), .A2(n522), .ZN(n373) );
  XOR2_X1 U440 ( .A(G22GAT), .B(G155GAT), .Z(n438) );
  XOR2_X1 U441 ( .A(n374), .B(n438), .Z(n377) );
  XOR2_X1 U442 ( .A(G15GAT), .B(G127GAT), .Z(n451) );
  XNOR2_X1 U443 ( .A(n375), .B(n451), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n390) );
  XOR2_X1 U445 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n379) );
  NAND2_X1 U446 ( .A1(G231GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U448 ( .A(n380), .B(KEYINPUT12), .Z(n388) );
  XOR2_X1 U449 ( .A(G78GAT), .B(G211GAT), .Z(n382) );
  XNOR2_X1 U450 ( .A(G183GAT), .B(G71GAT), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U452 ( .A(G64GAT), .B(KEYINPUT80), .Z(n384) );
  XNOR2_X1 U453 ( .A(G8GAT), .B(KEYINPUT81), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U456 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U457 ( .A(n390), .B(n389), .Z(n498) );
  NOR2_X1 U458 ( .A1(n391), .A2(n498), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n392), .B(KEYINPUT113), .ZN(n393) );
  INV_X1 U460 ( .A(n577), .ZN(n396) );
  NOR2_X1 U461 ( .A1(n393), .A2(n396), .ZN(n395) );
  XNOR2_X1 U462 ( .A(KEYINPUT36), .B(n396), .ZN(n598) );
  NAND2_X1 U463 ( .A1(n498), .A2(n598), .ZN(n398) );
  NAND2_X1 U464 ( .A1(n399), .A2(n592), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n400), .B(KEYINPUT115), .ZN(n401) );
  NAND2_X1 U466 ( .A1(n401), .A2(n587), .ZN(n402) );
  NAND2_X1 U467 ( .A1(n403), .A2(n402), .ZN(n405) );
  INV_X1 U468 ( .A(KEYINPUT48), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n551) );
  XOR2_X1 U470 ( .A(KEYINPUT17), .B(G183GAT), .Z(n407) );
  XNOR2_X1 U471 ( .A(KEYINPUT87), .B(KEYINPUT19), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U473 ( .A(n408), .B(KEYINPUT18), .Z(n410) );
  XNOR2_X1 U474 ( .A(KEYINPUT86), .B(KEYINPUT88), .ZN(n409) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n462) );
  NAND2_X1 U476 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n415), .B(KEYINPUT80), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n462), .B(n420), .ZN(n424) );
  XOR2_X1 U480 ( .A(KEYINPUT91), .B(G218GAT), .Z(n422) );
  XNOR2_X1 U481 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U483 ( .A(G197GAT), .B(n423), .Z(n443) );
  INV_X1 U484 ( .A(n542), .ZN(n425) );
  NOR2_X1 U485 ( .A1(n551), .A2(n425), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n428) );
  NOR2_X1 U487 ( .A1(n540), .A2(n428), .ZN(n586) );
  XOR2_X1 U488 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n430) );
  XNOR2_X1 U489 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n435) );
  XOR2_X1 U491 ( .A(n431), .B(G204GAT), .Z(n433) );
  NAND2_X1 U492 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n480) );
  NAND2_X1 U499 ( .A1(n586), .A2(n480), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n444), .B(KEYINPUT55), .ZN(n465) );
  XOR2_X1 U501 ( .A(G99GAT), .B(G134GAT), .Z(n446) );
  XNOR2_X1 U502 ( .A(G43GAT), .B(G190GAT), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U504 ( .A(KEYINPUT89), .B(KEYINPUT64), .Z(n448) );
  XNOR2_X1 U505 ( .A(G169GAT), .B(KEYINPUT85), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U507 ( .A(n450), .B(n449), .Z(n458) );
  XOR2_X1 U508 ( .A(n452), .B(n451), .Z(n454) );
  NAND2_X1 U509 ( .A1(G227GAT), .A2(G233GAT), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U511 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n458), .B(n457), .ZN(n464) );
  XOR2_X1 U513 ( .A(G176GAT), .B(KEYINPUT84), .Z(n460) );
  XNOR2_X1 U514 ( .A(KEYINPUT20), .B(KEYINPUT83), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U516 ( .A(n462), .B(n461), .Z(n463) );
  XNOR2_X1 U517 ( .A(n464), .B(n463), .ZN(n552) );
  NAND2_X1 U518 ( .A1(n465), .A2(n552), .ZN(n580) );
  NOR2_X1 U519 ( .A1(n577), .A2(n580), .ZN(n468) );
  INV_X1 U520 ( .A(G190GAT), .ZN(n466) );
  INV_X1 U521 ( .A(n498), .ZN(n595) );
  NAND2_X1 U522 ( .A1(n552), .A2(n542), .ZN(n469) );
  NAND2_X1 U523 ( .A1(n469), .A2(n480), .ZN(n470) );
  XNOR2_X1 U524 ( .A(n470), .B(KEYINPUT95), .ZN(n471) );
  XOR2_X1 U525 ( .A(KEYINPUT25), .B(n471), .Z(n475) );
  XNOR2_X1 U526 ( .A(KEYINPUT27), .B(n542), .ZN(n481) );
  NOR2_X1 U527 ( .A1(n552), .A2(n480), .ZN(n472) );
  XNOR2_X1 U528 ( .A(KEYINPUT26), .B(n472), .ZN(n585) );
  AND2_X1 U529 ( .A1(n481), .A2(n585), .ZN(n473) );
  XNOR2_X1 U530 ( .A(KEYINPUT94), .B(n473), .ZN(n474) );
  NOR2_X1 U531 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U532 ( .A1(n540), .A2(n476), .ZN(n478) );
  XNOR2_X1 U533 ( .A(n478), .B(n477), .ZN(n484) );
  XOR2_X1 U534 ( .A(KEYINPUT28), .B(KEYINPUT67), .Z(n479) );
  XNOR2_X1 U535 ( .A(n480), .B(n479), .ZN(n555) );
  NAND2_X1 U536 ( .A1(n540), .A2(n481), .ZN(n550) );
  NOR2_X1 U537 ( .A1(n552), .A2(n550), .ZN(n482) );
  NAND2_X1 U538 ( .A1(n555), .A2(n482), .ZN(n483) );
  NAND2_X1 U539 ( .A1(n484), .A2(n483), .ZN(n501) );
  NAND2_X1 U540 ( .A1(n595), .A2(n501), .ZN(n485) );
  XOR2_X1 U541 ( .A(KEYINPUT100), .B(n485), .Z(n486) );
  NAND2_X1 U542 ( .A1(n598), .A2(n486), .ZN(n487) );
  XNOR2_X1 U543 ( .A(KEYINPUT37), .B(n487), .ZN(n539) );
  INV_X1 U544 ( .A(n587), .ZN(n523) );
  NAND2_X1 U545 ( .A1(n523), .A2(n592), .ZN(n503) );
  INV_X1 U546 ( .A(n503), .ZN(n488) );
  NAND2_X1 U547 ( .A1(n539), .A2(n488), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT101), .B(KEYINPUT38), .ZN(n489) );
  NAND2_X1 U549 ( .A1(n519), .A2(n552), .ZN(n494) );
  XOR2_X1 U550 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n492) );
  NOR2_X1 U551 ( .A1(n595), .A2(n580), .ZN(n497) );
  XNOR2_X1 U552 ( .A(n495), .B(KEYINPUT124), .ZN(n496) );
  XNOR2_X1 U553 ( .A(n497), .B(n496), .ZN(G1350GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT97), .B(KEYINPUT34), .Z(n505) );
  XOR2_X1 U555 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n500) );
  NAND2_X1 U556 ( .A1(n498), .A2(n577), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n500), .B(n499), .ZN(n502) );
  NAND2_X1 U558 ( .A1(n502), .A2(n501), .ZN(n524) );
  NOR2_X1 U559 ( .A1(n503), .A2(n524), .ZN(n511) );
  NAND2_X1 U560 ( .A1(n511), .A2(n540), .ZN(n504) );
  XNOR2_X1 U561 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U562 ( .A(G1GAT), .B(n506), .ZN(G1324GAT) );
  NAND2_X1 U563 ( .A1(n511), .A2(n542), .ZN(n507) );
  XNOR2_X1 U564 ( .A(n507), .B(KEYINPUT98), .ZN(n508) );
  XNOR2_X1 U565 ( .A(G8GAT), .B(n508), .ZN(G1325GAT) );
  XOR2_X1 U566 ( .A(G15GAT), .B(KEYINPUT35), .Z(n510) );
  NAND2_X1 U567 ( .A1(n511), .A2(n552), .ZN(n509) );
  XNOR2_X1 U568 ( .A(n510), .B(n509), .ZN(G1326GAT) );
  INV_X1 U569 ( .A(n555), .ZN(n545) );
  NAND2_X1 U570 ( .A1(n545), .A2(n511), .ZN(n512) );
  XNOR2_X1 U571 ( .A(n512), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U572 ( .A1(n519), .A2(n540), .ZN(n517) );
  XOR2_X1 U573 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n514) );
  XNOR2_X1 U574 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n513) );
  XNOR2_X1 U575 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U576 ( .A(KEYINPUT99), .B(n515), .ZN(n516) );
  XNOR2_X1 U577 ( .A(n517), .B(n516), .ZN(G1328GAT) );
  NAND2_X1 U578 ( .A1(n519), .A2(n542), .ZN(n518) );
  XNOR2_X1 U579 ( .A(n518), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U580 ( .A(G50GAT), .B(KEYINPUT105), .Z(n521) );
  NAND2_X1 U581 ( .A1(n519), .A2(n545), .ZN(n520) );
  XNOR2_X1 U582 ( .A(n521), .B(n520), .ZN(G1331GAT) );
  NOR2_X1 U583 ( .A1(n522), .A2(n523), .ZN(n538) );
  INV_X1 U584 ( .A(n538), .ZN(n525) );
  NOR2_X1 U585 ( .A1(n525), .A2(n524), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n534), .A2(n540), .ZN(n528) );
  XNOR2_X1 U587 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n526) );
  XNOR2_X1 U588 ( .A(n526), .B(KEYINPUT42), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n528), .B(n527), .ZN(G1332GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n530) );
  NAND2_X1 U591 ( .A1(n534), .A2(n542), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U593 ( .A(G64GAT), .B(n531), .ZN(G1333GAT) );
  XOR2_X1 U594 ( .A(G71GAT), .B(KEYINPUT109), .Z(n533) );
  NAND2_X1 U595 ( .A1(n534), .A2(n552), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1334GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n536) );
  NAND2_X1 U598 ( .A1(n534), .A2(n545), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U600 ( .A(G78GAT), .B(n537), .ZN(G1335GAT) );
  AND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n546), .A2(n540), .ZN(n541) );
  XNOR2_X1 U603 ( .A(n541), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U604 ( .A1(n546), .A2(n542), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U606 ( .A1(n552), .A2(n546), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n544), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n548) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U611 ( .A(G106GAT), .B(n549), .ZN(G1339GAT) );
  NOR2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n565) );
  NAND2_X1 U613 ( .A1(n565), .A2(n552), .ZN(n553) );
  XOR2_X1 U614 ( .A(KEYINPUT116), .B(n553), .Z(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n562) );
  NOR2_X1 U616 ( .A1(n587), .A2(n562), .ZN(n556) );
  XOR2_X1 U617 ( .A(G113GAT), .B(n556), .Z(G1340GAT) );
  NOR2_X1 U618 ( .A1(n522), .A2(n562), .ZN(n558) );
  XNOR2_X1 U619 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n558), .B(n557), .ZN(G1341GAT) );
  NOR2_X1 U621 ( .A1(n595), .A2(n562), .ZN(n560) );
  XNOR2_X1 U622 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U624 ( .A(G127GAT), .B(n561), .ZN(G1342GAT) );
  NOR2_X1 U625 ( .A1(n577), .A2(n562), .ZN(n564) );
  XNOR2_X1 U626 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n564), .B(n563), .ZN(G1343GAT) );
  NAND2_X1 U628 ( .A1(n565), .A2(n585), .ZN(n576) );
  NOR2_X1 U629 ( .A1(n587), .A2(n576), .ZN(n567) );
  XNOR2_X1 U630 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U632 ( .A(G141GAT), .B(n568), .ZN(G1344GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n570) );
  XNOR2_X1 U634 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n572) );
  NOR2_X1 U636 ( .A1(n522), .A2(n576), .ZN(n571) );
  XOR2_X1 U637 ( .A(n572), .B(n571), .Z(G1345GAT) );
  NOR2_X1 U638 ( .A1(n595), .A2(n576), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G155GAT), .B(n575), .ZN(G1346GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(G162GAT), .B(n578), .Z(G1347GAT) );
  NOR2_X1 U644 ( .A1(n587), .A2(n580), .ZN(n579) );
  XOR2_X1 U645 ( .A(G169GAT), .B(n579), .Z(G1348GAT) );
  NOR2_X1 U646 ( .A1(n580), .A2(n522), .ZN(n584) );
  XOR2_X1 U647 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n582) );
  XNOR2_X1 U648 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1349GAT) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n597) );
  NOR2_X1 U652 ( .A1(n587), .A2(n597), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1352GAT) );
  NOR2_X1 U657 ( .A1(n592), .A2(n597), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n594), .B(n593), .ZN(G1353GAT) );
  NOR2_X1 U660 ( .A1(n595), .A2(n597), .ZN(n596) );
  XOR2_X1 U661 ( .A(G211GAT), .B(n596), .Z(G1354GAT) );
  INV_X1 U662 ( .A(n597), .ZN(n599) );
  NAND2_X1 U663 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U664 ( .A(n600), .B(KEYINPUT127), .ZN(n601) );
  XOR2_X1 U665 ( .A(n601), .B(KEYINPUT126), .Z(n603) );
  XNOR2_X1 U666 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n602) );
  XNOR2_X1 U667 ( .A(n603), .B(n602), .ZN(G1355GAT) );
endmodule

