//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n574, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(KEYINPUT67), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n473), .A2(G137), .A3(new_n474), .A4(new_n463), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT67), .B(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n469), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n482));
  INV_X1    g057(.A(new_n463), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(new_n476), .B2(KEYINPUT3), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n473), .A2(new_n474), .A3(new_n463), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n487), .B1(G136), .B2(new_n489), .ZN(G162));
  NAND4_X1  g065(.A1(new_n473), .A2(G126), .A3(G2105), .A4(new_n463), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n474), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(new_n474), .A3(G138), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n466), .A2(KEYINPUT68), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT3), .B(G2104), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n500), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n500), .A2(G2105), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n473), .A2(new_n463), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n494), .B1(new_n503), .B2(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n508), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n511), .A2(new_n515), .ZN(G166));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  INV_X1    g092(.A(G51), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n513), .A2(KEYINPUT69), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n520), .B1(new_n513), .B2(KEYINPUT69), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n519), .A2(new_n521), .A3(KEYINPUT70), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n518), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT71), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(G63), .A2(G651), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n514), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(new_n508), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n517), .B1(new_n526), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n529), .A2(new_n530), .B1(new_n508), .B2(new_n534), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n519), .A2(new_n521), .A3(KEYINPUT70), .ZN(new_n539));
  AOI21_X1  g114(.A(KEYINPUT70), .B1(new_n519), .B2(new_n521), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g116(.A(KEYINPUT72), .B(new_n538), .C1(new_n541), .C2(new_n518), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n537), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(new_n524), .A2(new_n525), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT73), .B(G52), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n508), .A2(new_n513), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n547), .A2(new_n510), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(G171));
  AOI22_X1  g128(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n554), .A2(new_n510), .B1(new_n548), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G43), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n541), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND3_X1  g140(.A1(new_n519), .A2(new_n521), .A3(G53), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR3_X1    g143(.A1(new_n568), .A2(KEYINPUT74), .A3(new_n510), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT74), .B1(new_n568), .B2(new_n510), .ZN(new_n570));
  INV_X1    g145(.A(new_n548), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n569), .A2(new_n570), .B1(G91), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n567), .A2(new_n572), .ZN(G299));
  XNOR2_X1  g148(.A(new_n552), .B(KEYINPUT75), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND3_X1  g152(.A1(new_n519), .A2(new_n521), .A3(G49), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n571), .A2(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  AND2_X1   g156(.A1(G48), .A2(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n513), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n510), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n548), .A2(new_n586), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n585), .A2(new_n587), .ZN(G305));
  AND2_X1   g163(.A1(new_n544), .A2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n590), .A2(new_n510), .B1(new_n548), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n589), .A2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(new_n544), .A2(G54), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n571), .A2(KEYINPUT10), .A3(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n548), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  XOR2_X1   g174(.A(KEYINPUT5), .B(G543), .Z(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n595), .A2(new_n598), .B1(G651), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n574), .B2(G868), .ZN(G284));
  AOI21_X1  g181(.A(new_n605), .B1(new_n574), .B2(G868), .ZN(G321));
  NOR2_X1   g182(.A1(G299), .A2(G868), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g184(.A(new_n608), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(new_n604), .ZN(new_n611));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G860), .ZN(G148));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n559), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n604), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n477), .A2(new_n499), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n489), .A2(G135), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n473), .A2(G2105), .A3(new_n463), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G123), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n474), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n623), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n622), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT76), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2430), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT77), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  NOR2_X1   g222(.A1(G2072), .A2(G2078), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n442), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT78), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT80), .Z(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(KEYINPUT79), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n649), .A2(KEYINPUT79), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n653), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n658), .B(new_n659), .C1(new_n652), .C2(new_n650), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n652), .A2(new_n659), .A3(new_n649), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT18), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  MUX2_X1   g250(.A(new_n675), .B(new_n674), .S(new_n667), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT81), .ZN(new_n678));
  INV_X1    g253(.A(G1981), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT82), .B(KEYINPUT83), .Z(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT84), .ZN(new_n686));
  INV_X1    g261(.A(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n684), .B(new_n688), .ZN(G229));
  XOR2_X1   g264(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n690));
  NAND3_X1  g265(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G139), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n488), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT89), .Z(new_n695));
  AOI22_X1  g270(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(new_n474), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G33), .B(new_n698), .S(G29), .Z(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(G2072), .Z(new_n700));
  INV_X1    g275(.A(G2084), .ZN(new_n701));
  INV_X1    g276(.A(G34), .ZN(new_n702));
  AOI21_X1  g277(.A(G29), .B1(new_n702), .B2(KEYINPUT24), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(KEYINPUT24), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n479), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT27), .B(G1996), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n489), .A2(G141), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n624), .A2(G129), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT26), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n477), .A2(G105), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n708), .A2(new_n709), .A3(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(new_n705), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n716), .B(KEYINPUT90), .C1(G29), .C2(G32), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(KEYINPUT90), .B2(new_n716), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n700), .B1(new_n701), .B2(new_n706), .C1(new_n707), .C2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT91), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G5), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G171), .B2(new_n721), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(G1961), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n718), .A2(new_n707), .ZN(new_n725));
  NOR2_X1   g300(.A1(G16), .A2(G19), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n560), .B2(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G1341), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n706), .A2(new_n701), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT94), .Z(new_n730));
  NAND4_X1  g305(.A1(new_n724), .A2(new_n725), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n723), .A2(G1961), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT93), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n721), .A2(G21), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G168), .B2(new_n721), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n733), .B1(G1966), .B2(new_n735), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n731), .B(new_n736), .C1(G1966), .C2(new_n735), .ZN(new_n737));
  NOR2_X1   g312(.A1(G29), .A2(G35), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G162), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2090), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT96), .B(KEYINPUT23), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n721), .A2(G20), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G299), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT97), .B(G1956), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n742), .A2(new_n748), .A3(KEYINPUT98), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n727), .A2(G1341), .ZN(new_n750));
  NAND2_X1  g325(.A1(G164), .A2(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G27), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT31), .B(G11), .Z(new_n755));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n705), .B1(new_n756), .B2(G28), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(KEYINPUT92), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n757), .A2(KEYINPUT92), .B1(new_n756), .B2(G28), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n754), .B(new_n760), .C1(new_n705), .C2(new_n628), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n489), .A2(G140), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n624), .A2(G128), .ZN(new_n763));
  OR2_X1    g338(.A1(G104), .A2(G2105), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n764), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G29), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n705), .A2(G26), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT28), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n752), .A2(new_n753), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n750), .A2(new_n761), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n721), .A2(G4), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n611), .B2(new_n721), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(G1348), .Z(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n776), .C1(G2090), .C2(new_n741), .ZN(new_n777));
  AOI21_X1  g352(.A(KEYINPUT98), .B1(new_n742), .B2(new_n748), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n720), .A2(new_n737), .A3(new_n749), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n721), .A2(G6), .ZN(new_n781));
  INV_X1    g356(.A(G305), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n721), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT86), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT32), .B(G1981), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n721), .A2(G22), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G166), .B2(new_n721), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1971), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n721), .A2(G23), .ZN(new_n790));
  INV_X1    g365(.A(G288), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n721), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT33), .B(G1976), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT87), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n789), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n786), .B(new_n796), .C1(new_n795), .C2(new_n794), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT34), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(KEYINPUT34), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n589), .A2(new_n592), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(new_n721), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n721), .B2(G24), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(new_n687), .ZN(new_n803));
  OR2_X1    g378(.A1(G95), .A2(G2105), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n804), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT85), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n489), .A2(G131), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n624), .A2(G119), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G25), .B(new_n809), .S(G29), .Z(new_n810));
  XOR2_X1   g385(.A(KEYINPUT35), .B(G1991), .Z(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n810), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n802), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G1986), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n798), .A2(new_n799), .A3(new_n803), .A4(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT36), .Z(new_n817));
  NOR2_X1   g392(.A1(new_n780), .A2(new_n817), .ZN(G311));
  INV_X1    g393(.A(G311), .ZN(G150));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n524), .B2(new_n525), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n571), .A2(G93), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n820), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  OAI211_X1 g400(.A(KEYINPUT99), .B(new_n823), .C1(new_n541), .C2(new_n821), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n510), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT101), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT37), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n611), .A2(G559), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n831), .A2(new_n559), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n827), .A2(new_n560), .A3(new_n830), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n836), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT100), .ZN(new_n843));
  INV_X1    g418(.A(G860), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n840), .B2(new_n841), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n834), .B1(new_n843), .B2(new_n845), .ZN(G145));
  XOR2_X1   g421(.A(new_n715), .B(new_n766), .Z(new_n847));
  AOI21_X1  g422(.A(new_n495), .B1(new_n484), .B2(new_n504), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT68), .B1(new_n466), .B2(new_n496), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n499), .A2(new_n498), .A3(new_n501), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n491), .B(new_n493), .C1(new_n848), .C2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(G164), .A2(KEYINPUT102), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n847), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT103), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n698), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n847), .A2(new_n856), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n695), .A2(KEYINPUT103), .A3(new_n697), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n809), .B(new_n620), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n624), .A2(G130), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n474), .A2(G118), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(G142), .B2(new_n489), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n864), .B(new_n869), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n863), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n628), .B(G160), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G162), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n873), .B2(new_n871), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g451(.A1(G290), .A2(new_n782), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n800), .A2(G305), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(G288), .B(G166), .Z(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n880), .A3(new_n878), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(KEYINPUT42), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n882), .A2(KEYINPUT104), .A3(new_n883), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT104), .B1(new_n882), .B2(new_n883), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n885), .B1(new_n888), .B2(KEYINPUT42), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n839), .B(new_n616), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n604), .A2(G299), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n604), .A2(G299), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n894), .A2(KEYINPUT41), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(KEYINPUT41), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n894), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(new_n891), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n890), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n889), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G868), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n831), .A2(new_n614), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(G295));
  NAND2_X1  g482(.A1(G295), .A2(KEYINPUT105), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n909), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(G331));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n837), .A2(new_n912), .A3(new_n838), .ZN(new_n913));
  AOI211_X1 g488(.A(new_n829), .B(new_n559), .C1(new_n825), .C2(new_n826), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n560), .B1(new_n827), .B2(new_n830), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT106), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(G168), .A2(G171), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n574), .B2(G168), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n913), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n913), .B2(new_n916), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n920), .A2(new_n921), .A3(new_n894), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n913), .A2(new_n916), .ZN(new_n923));
  INV_X1    g498(.A(new_n918), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n897), .B1(new_n925), .B2(new_n919), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n886), .A2(new_n887), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n922), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n922), .B2(new_n926), .ZN(new_n929));
  INV_X1    g504(.A(G37), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n931), .B2(KEYINPUT107), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT43), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n928), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n895), .A2(KEYINPUT108), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT108), .ZN(new_n938));
  AOI211_X1 g513(.A(new_n937), .B(new_n938), .C1(new_n919), .C2(new_n925), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n927), .B1(new_n939), .B2(new_n922), .ZN(new_n940));
  AND4_X1   g515(.A1(KEYINPUT43), .A2(new_n936), .A3(new_n940), .A4(new_n930), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT44), .B1(new_n935), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(new_n932), .B2(new_n934), .ZN(new_n945));
  AND4_X1   g520(.A1(new_n944), .A2(new_n936), .A3(new_n940), .A4(new_n930), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n947), .ZN(G397));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n854), .A2(new_n855), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n469), .A2(G40), .A3(new_n478), .A4(new_n475), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n687), .A3(new_n800), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT48), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n809), .B(new_n812), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT109), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n959), .A2(KEYINPUT109), .ZN(new_n962));
  INV_X1    g537(.A(G1996), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n715), .B(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G2067), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n766), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n961), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(new_n954), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT127), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n958), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n956), .A2(new_n957), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n971), .B(new_n972), .C1(new_n970), .C2(new_n969), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n967), .A2(new_n812), .A3(new_n809), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n766), .A2(G2067), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n955), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n966), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n955), .B1(new_n715), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n954), .A2(G1996), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n978), .B1(KEYINPUT46), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(KEYINPUT46), .B2(new_n979), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT47), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT126), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n973), .B(new_n976), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n983), .B2(new_n982), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n951), .A2(G1384), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n854), .A2(new_n855), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n951), .B1(G164), .B2(G1384), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n753), .A3(new_n953), .A4(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n952), .B1(new_n852), .B2(new_n986), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(new_n988), .A3(KEYINPUT53), .A4(new_n753), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n852), .B2(new_n949), .ZN(new_n995));
  NOR2_X1   g570(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n953), .B1(G164), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT118), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1961), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n952), .B1(new_n852), .B2(new_n996), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n999), .A2(new_n1000), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n991), .A2(new_n993), .A3(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1006), .A2(new_n574), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n953), .A2(new_n852), .A3(new_n949), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1008), .A2(G8), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G73), .A2(G543), .ZN(new_n1011));
  INV_X1    g586(.A(G61), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(new_n600), .B2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1013), .A2(G651), .B1(new_n513), .B2(new_n582), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT112), .B(G86), .Z(new_n1015));
  NAND2_X1  g590(.A1(new_n571), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n679), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n585), .A2(G1981), .A3(new_n587), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1010), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT49), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1010), .B(new_n1021), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1009), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n791), .A2(G1976), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1008), .A2(new_n1024), .A3(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1009), .A2(new_n1024), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1009), .A2(KEYINPUT111), .A3(new_n1024), .A4(new_n1029), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1027), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT45), .B1(new_n852), .B2(new_n949), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(new_n952), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1971), .B1(new_n1036), .B2(new_n987), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(G2090), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G303), .A2(G8), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT55), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1036), .A2(new_n987), .ZN(new_n1045));
  INV_X1    g620(.A(G1971), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1039), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1042), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1007), .A2(new_n1034), .A3(new_n1043), .A4(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n537), .A2(new_n542), .A3(G8), .ZN(new_n1053));
  INV_X1    g628(.A(G1966), .ZN(new_n1054));
  INV_X1    g629(.A(new_n986), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n953), .B1(G164), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1054), .B1(new_n1035), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1001), .A2(new_n1002), .A3(new_n701), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1053), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1001), .A2(new_n1002), .A3(new_n701), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1966), .B1(new_n992), .B2(new_n988), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1061), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1044), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT122), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1069));
  OAI211_X1 g644(.A(KEYINPUT51), .B(G8), .C1(new_n1069), .C2(G286), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1066), .A2(new_n1068), .B1(new_n1070), .B2(KEYINPUT121), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1053), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1072), .B(KEYINPUT51), .C1(new_n1067), .C2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1059), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1052), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1061), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n1068), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1070), .A2(KEYINPUT121), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n1074), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1059), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1078), .B1(new_n1085), .B2(KEYINPUT62), .ZN(new_n1086));
  AOI211_X1 g661(.A(KEYINPUT123), .B(new_n1076), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1077), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(KEYINPUT124), .B(new_n1077), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n791), .A2(new_n1028), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(KEYINPUT115), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1009), .B1(new_n1094), .B2(new_n1018), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1034), .A2(KEYINPUT114), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1034), .A2(KEYINPUT114), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1095), .B1(new_n1098), .B2(new_n1051), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n1100));
  INV_X1    g675(.A(G1956), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n995), .B2(new_n998), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1038), .A2(KEYINPUT117), .A3(new_n1101), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n506), .A2(new_n849), .A3(new_n850), .ZN(new_n1106));
  INV_X1    g681(.A(new_n494), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1106), .A2(KEYINPUT102), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT102), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n1055), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n988), .A2(new_n953), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1104), .A2(new_n1105), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n567), .B2(new_n572), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1100), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1008), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n965), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n999), .A2(new_n1004), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(G1348), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n611), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1036), .A2(new_n987), .A3(new_n1113), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1105), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT117), .B1(new_n1038), .B2(new_n1101), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1118), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(KEYINPUT119), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1119), .A2(new_n1124), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(new_n1118), .A3(new_n1125), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1119), .A2(new_n1136), .A3(new_n1130), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1133), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1118), .B1(new_n1132), .B2(new_n1125), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1135), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT60), .B(new_n1121), .C1(new_n1122), .C2(G1348), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1141), .A2(new_n611), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1137), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1045), .B2(G1996), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1112), .A2(KEYINPUT120), .A3(new_n963), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT58), .B(G1341), .Z(new_n1147));
  NAND2_X1  g722(.A1(new_n1008), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n560), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1149), .A2(KEYINPUT59), .A3(new_n560), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1123), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(new_n611), .A3(new_n1141), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1152), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1134), .B1(new_n1143), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n950), .A2(new_n951), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n952), .A2(new_n990), .A3(G2078), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(new_n987), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n991), .A2(new_n1005), .A3(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1163), .A2(new_n574), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1159), .B1(new_n1007), .B2(new_n1164), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1051), .A2(new_n1034), .A3(new_n1043), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(G171), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1167), .B(KEYINPUT54), .C1(new_n574), .C2(new_n1006), .ZN(new_n1168));
  AND4_X1   g743(.A1(new_n1085), .A2(new_n1165), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1099), .B1(new_n1158), .B2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1040), .B(new_n1050), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1171), .A2(G168), .A3(new_n1067), .A4(new_n1034), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT116), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1172), .A2(KEYINPUT116), .A3(new_n1173), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1064), .A2(new_n1173), .A3(G286), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1171), .B(new_n1178), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1090), .A2(new_n1091), .A3(new_n1170), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n800), .B(new_n687), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n969), .B1(new_n955), .B2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT110), .Z(new_n1185));
  AND3_X1   g760(.A1(new_n1181), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1182), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n985), .B1(new_n1186), .B2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g763(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1190));
  OAI211_X1 g764(.A(new_n1190), .B(new_n875), .C1(new_n945), .C2(new_n946), .ZN(G225));
  INV_X1    g765(.A(G225), .ZN(G308));
endmodule


