//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n449, new_n451, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n562, new_n563, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1104, new_n1105, new_n1106,
    new_n1107;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n465), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  AND3_X1   g048(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(KEYINPUT3), .B1(KEYINPUT68), .B2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n463), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  INV_X1    g056(.A(new_n476), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OAI21_X1  g058(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OR2_X1    g065(.A1(new_n466), .A2(new_n467), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n463), .C1(new_n474), .C2(new_n475), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  OAI21_X1  g075(.A(G2105), .B1(new_n500), .B2(G114), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n500), .A2(G114), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(G2105), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT70), .A3(new_n499), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g086(.A(G126), .B(G2105), .C1(new_n474), .C2(new_n475), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n497), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT71), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n515), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n525), .A2(KEYINPUT72), .A3(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n518), .A2(new_n520), .B1(KEYINPUT5), .B2(new_n517), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT6), .B(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n531), .A2(G543), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n533), .A2(G88), .B1(G50), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n528), .A2(new_n529), .A3(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  NAND2_X1  g112(.A1(new_n533), .A2(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT73), .B(G51), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n538), .A2(new_n539), .A3(new_n541), .A4(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  AOI22_X1  g120(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G651), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  INV_X1    g124(.A(G52), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n531), .A2(G543), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n532), .A2(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n548), .A2(new_n552), .ZN(G171));
  AOI22_X1  g128(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n547), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT74), .B(G43), .Z(new_n557));
  OAI22_X1  g132(.A1(new_n532), .A2(new_n556), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT75), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT76), .ZN(G188));
  XNOR2_X1  g141(.A(new_n530), .B(KEYINPUT78), .ZN(new_n567));
  XOR2_X1   g142(.A(KEYINPUT79), .B(G65), .Z(new_n568));
  AND2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g144(.A1(G78), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n533), .A2(KEYINPUT77), .A3(G91), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n532), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT9), .B1(new_n551), .B2(new_n576), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n551), .A2(KEYINPUT9), .A3(new_n576), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n572), .A2(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n571), .A2(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  OAI21_X1  g156(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n534), .A2(G49), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n530), .A2(G87), .A3(new_n531), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  INV_X1    g161(.A(G48), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n532), .A2(new_n586), .B1(new_n587), .B2(new_n551), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n530), .A2(G61), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n547), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n533), .A2(G85), .B1(G47), .B2(new_n534), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n547), .B2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT80), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n567), .B2(G66), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(new_n547), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n533), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n532), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n603), .A2(new_n606), .B1(G54), .B2(new_n534), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  INV_X1    g192(.A(new_n559), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n612), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n608), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g196(.A(KEYINPUT81), .B(KEYINPUT11), .ZN(new_n622));
  XNOR2_X1  g197(.A(G323), .B(new_n622), .ZN(G282));
  NAND2_X1  g198(.A1(new_n491), .A2(new_n472), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT82), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT83), .ZN(new_n631));
  AOI22_X1  g206(.A1(G135), .A2(new_n482), .B1(new_n485), .B2(G123), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(G111), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n633), .A2(KEYINPUT84), .B1(new_n634), .B2(G2105), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(KEYINPUT84), .B2(new_n633), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G2096), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n629), .A2(new_n631), .A3(new_n639), .ZN(G156));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n627), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n638), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n669), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G229));
  MUX2_X1   g260(.A(G6), .B(G305), .S(G16), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT32), .ZN(new_n687));
  INV_X1    g262(.A(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G22), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G166), .B2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT88), .ZN(new_n693));
  INV_X1    g268(.A(G1971), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(G23), .ZN(new_n697));
  INV_X1    g272(.A(G288), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n690), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT87), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT33), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n689), .A2(new_n695), .A3(new_n696), .A4(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(KEYINPUT34), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n482), .A2(G131), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n485), .A2(G119), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT85), .B1(G95), .B2(G2105), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g284(.A1(KEYINPUT85), .A2(G95), .A3(G2105), .ZN(new_n710));
  OAI221_X1 g285(.A(G2104), .B1(G107), .B2(new_n463), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n706), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G25), .B(new_n712), .S(G29), .Z(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n717), .A2(KEYINPUT86), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(KEYINPUT86), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n690), .A2(G24), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G290), .B2(G16), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(G1986), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n722), .A2(G1986), .ZN(new_n724));
  NOR4_X1   g299(.A1(new_n718), .A2(new_n719), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n704), .A2(new_n705), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT89), .B(KEYINPUT36), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT98), .B1(G29), .B2(G32), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT97), .B(KEYINPUT26), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n472), .A2(G105), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT96), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n732), .B(new_n734), .C1(G129), .C2(new_n485), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n482), .A2(G141), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(new_n729), .B(KEYINPUT98), .S(new_n739), .Z(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G16), .A2(G19), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n559), .B2(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G1341), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n690), .A2(G21), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G168), .B2(new_n690), .ZN(new_n747));
  INV_X1    g322(.A(G2072), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n738), .A2(G33), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n482), .A2(G139), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT25), .Z(new_n752));
  AOI22_X1  g327(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n750), .B(new_n752), .C1(new_n753), .C2(new_n463), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n749), .B1(new_n754), .B2(G29), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n747), .A2(G1966), .B1(new_n748), .B2(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n744), .A2(G1341), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n742), .A2(new_n745), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT30), .B(G28), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n759), .A2(new_n738), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n637), .B2(new_n738), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT99), .Z(new_n764));
  INV_X1    g339(.A(G2078), .ZN(new_n765));
  NAND2_X1  g340(.A1(G164), .A2(G29), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G27), .B2(G29), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n764), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n768), .B1(new_n765), .B2(new_n767), .C1(new_n740), .C2(new_n741), .ZN(new_n769));
  INV_X1    g344(.A(new_n747), .ZN(new_n770));
  INV_X1    g345(.A(G1966), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n738), .A2(G26), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT28), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n482), .A2(G140), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n485), .A2(G128), .ZN(new_n775));
  OR2_X1    g350(.A1(G104), .A2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n776), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n773), .B1(new_n778), .B2(G29), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT91), .B(G2067), .Z(new_n780));
  AOI22_X1  g355(.A1(new_n770), .A2(new_n771), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n690), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n690), .ZN(new_n783));
  INV_X1    g358(.A(G1961), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n781), .B(new_n785), .C1(new_n779), .C2(new_n780), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n758), .A2(new_n769), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G4), .A2(G16), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n609), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT90), .Z(new_n790));
  INV_X1    g365(.A(G1348), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n787), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n738), .A2(G35), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G162), .B2(new_n738), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT29), .Z(new_n797));
  INV_X1    g372(.A(G2090), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT100), .Z(new_n800));
  NOR2_X1   g375(.A1(new_n755), .A2(new_n748), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT95), .ZN(new_n802));
  AND2_X1   g377(.A1(KEYINPUT24), .A2(G34), .ZN(new_n803));
  NOR2_X1   g378(.A1(KEYINPUT24), .A2(G34), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n738), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT92), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n480), .B2(new_n738), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT93), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(G2084), .ZN(new_n810));
  AOI211_X1 g385(.A(new_n802), .B(new_n810), .C1(new_n798), .C2(new_n797), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n800), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n690), .A2(G20), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT23), .Z(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G299), .B2(G16), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1956), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n809), .A2(G2084), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT94), .Z(new_n818));
  NAND4_X1  g393(.A1(new_n794), .A2(new_n812), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n728), .A2(new_n819), .ZN(G311));
  INV_X1    g395(.A(G311), .ZN(G150));
  XOR2_X1   g396(.A(KEYINPUT102), .B(G93), .Z(new_n822));
  AOI22_X1  g397(.A1(new_n533), .A2(new_n822), .B1(G55), .B2(new_n534), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT101), .ZN(new_n825));
  OAI21_X1  g400(.A(G651), .B1(new_n824), .B2(KEYINPUT101), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G860), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  AOI21_X1  g404(.A(new_n559), .B1(new_n827), .B2(KEYINPUT103), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(KEYINPUT103), .B2(new_n827), .ZN(new_n831));
  OR3_X1    g406(.A1(new_n827), .A2(new_n618), .A3(KEYINPUT103), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n609), .A2(G559), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n833), .B(new_n834), .Z(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n838), .B2(KEYINPUT39), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n829), .B1(new_n839), .B2(new_n841), .ZN(G145));
  XNOR2_X1  g417(.A(new_n737), .B(new_n754), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n625), .B(new_n712), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n778), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n513), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n482), .A2(G142), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT105), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n485), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n463), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n847), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n845), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n637), .B(new_n480), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n489), .ZN(new_n857));
  AOI21_X1  g432(.A(G37), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n855), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(G395));
  NAND2_X1  g436(.A1(new_n827), .A2(new_n612), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n608), .B(G299), .Z(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(KEYINPUT41), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(KEYINPUT41), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n833), .B(new_n620), .ZN(new_n867));
  INV_X1    g442(.A(new_n863), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT107), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n866), .A2(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  XNOR2_X1  g447(.A(G303), .B(G290), .ZN(new_n873));
  XNOR2_X1  g448(.A(G305), .B(new_n698), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT42), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n872), .B(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n862), .B1(new_n877), .B2(new_n612), .ZN(G295));
  OAI21_X1  g453(.A(new_n862), .B1(new_n877), .B2(new_n612), .ZN(G331));
  XNOR2_X1  g454(.A(G286), .B(G171), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n833), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(new_n864), .A3(new_n865), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n863), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n875), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  INV_X1    g462(.A(new_n875), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n888), .A3(new_n884), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT43), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(KEYINPUT43), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT108), .B1(new_n890), .B2(KEYINPUT43), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  OAI22_X1  g470(.A1(new_n892), .A2(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n890), .A2(KEYINPUT43), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n897), .A2(KEYINPUT108), .A3(KEYINPUT44), .A4(new_n891), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(G397));
  INV_X1    g474(.A(G1384), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n463), .B1(KEYINPUT69), .B2(new_n502), .ZN(new_n901));
  AOI211_X1 g476(.A(new_n505), .B(new_n498), .C1(new_n901), .C2(new_n507), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT70), .B1(new_n509), .B2(new_n499), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n512), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n491), .A2(new_n493), .B1(new_n495), .B2(KEYINPUT4), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(KEYINPUT109), .B(G40), .Z(new_n910));
  NOR3_X1   g485(.A1(new_n470), .A2(new_n478), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT110), .ZN(new_n913));
  INV_X1    g488(.A(G2067), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n778), .B(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n737), .ZN(new_n916));
  INV_X1    g491(.A(G1996), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n912), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n917), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n919), .B1(new_n737), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n712), .B(new_n715), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n922), .B1(new_n923), .B2(new_n913), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(G290), .B(G1986), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n911), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n506), .A2(new_n510), .B1(new_n485), .B2(G126), .ZN(new_n929));
  AOI21_X1  g504(.A(G1384), .B1(new_n929), .B2(new_n497), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT50), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT118), .B(G2084), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n906), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT111), .B1(new_n906), .B2(KEYINPUT50), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n932), .B(new_n933), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n900), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n908), .A2(new_n911), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n771), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(G168), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(G8), .ZN(new_n941));
  AOI21_X1  g516(.A(G168), .B1(new_n936), .B2(new_n939), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT51), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT124), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n940), .A2(new_n945), .A3(G8), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n944), .B1(new_n943), .B2(new_n946), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT62), .ZN(new_n949));
  OR3_X1    g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n938), .A2(new_n694), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n952));
  XNOR2_X1  g527(.A(KEYINPUT112), .B(G2090), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(G303), .A2(G8), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n958), .A3(G8), .ZN(new_n959));
  INV_X1    g534(.A(new_n957), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n956), .B(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n911), .B1(new_n906), .B2(KEYINPUT50), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n931), .B1(new_n513), .B2(new_n900), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n964), .A2(new_n953), .B1(new_n938), .B2(new_n694), .ZN(new_n965));
  INV_X1    g540(.A(G8), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n961), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n513), .A2(new_n911), .A3(new_n900), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  AND2_X1   g544(.A1(G288), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n582), .A2(new_n583), .A3(G1976), .A4(new_n584), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n968), .A2(new_n970), .A3(G8), .A4(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n968), .A2(G8), .A3(new_n973), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n971), .B2(new_n972), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n974), .B(new_n975), .C1(new_n977), .C2(new_n979), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n968), .A2(G8), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n688), .B1(new_n589), .B2(new_n593), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n588), .A2(new_n592), .A3(G1981), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT116), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n983), .B1(new_n986), .B2(KEYINPUT49), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT116), .B(new_n988), .C1(new_n984), .C2(new_n985), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n981), .A2(new_n982), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n959), .A2(new_n967), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n908), .A2(new_n765), .A3(new_n911), .A4(new_n937), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n952), .A2(new_n784), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n993), .A2(new_n992), .ZN(new_n995));
  AOI21_X1  g570(.A(G301), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n949), .B1(new_n947), .B2(new_n948), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n950), .A2(new_n991), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n987), .A2(new_n989), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(new_n969), .A3(new_n698), .ZN(new_n1000));
  INV_X1    g575(.A(new_n985), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n983), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n981), .A2(new_n982), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n999), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT117), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n990), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n959), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1002), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n990), .B(KEYINPUT117), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n955), .A2(G8), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n961), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n966), .B(G286), .C1(new_n936), .C2(new_n939), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1013), .A2(KEYINPUT63), .A3(new_n959), .A4(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT63), .B1(new_n991), .B2(new_n1014), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1010), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(G299), .B(KEYINPUT57), .ZN(new_n1019));
  INV_X1    g594(.A(G1956), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT119), .B(new_n1020), .C1(new_n962), .C2(new_n963), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n906), .A2(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n513), .A2(new_n931), .A3(new_n900), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n911), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT119), .B1(new_n1025), .B2(new_n1020), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT56), .B(G2072), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n908), .A2(new_n911), .A3(new_n937), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1019), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n1033));
  XNOR2_X1  g608(.A(G299), .B(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1029), .B(KEYINPUT120), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1020), .B1(new_n962), .B2(new_n963), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1021), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1034), .A2(new_n1035), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1032), .A2(KEYINPUT61), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT122), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1032), .A2(KEYINPUT122), .A3(new_n1040), .A4(KEYINPUT61), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT61), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1040), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1034), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT58), .B(G1341), .Z(new_n1049));
  NAND2_X1  g624(.A1(new_n968), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT121), .B(G1996), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n938), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1052), .A2(new_n1053), .A3(new_n559), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1052), .B2(new_n559), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT60), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n608), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n930), .A2(new_n914), .A3(new_n911), .ZN(new_n1058));
  INV_X1    g633(.A(new_n935), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n963), .A2(KEYINPUT111), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n962), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1057), .B(new_n1058), .C1(new_n1061), .C2(G1348), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n607), .B(KEYINPUT60), .C1(new_n547), .C2(new_n601), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1054), .A2(new_n1055), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1043), .A2(new_n1044), .A3(new_n1048), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n952), .A2(new_n791), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n608), .B1(new_n1070), .B2(new_n1058), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1047), .B1(new_n1040), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n765), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n908), .A2(G160), .A3(new_n937), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n993), .A2(new_n992), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1075), .B(new_n1076), .C1(new_n1061), .C2(G1961), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n994), .A2(G301), .A3(new_n995), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(KEYINPUT54), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1077), .A2(G171), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(new_n996), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n991), .B(new_n1080), .C1(new_n1082), .C2(KEYINPUT54), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1083), .A2(new_n947), .A3(new_n948), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1018), .B1(new_n1073), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT125), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n998), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g662(.A(KEYINPUT125), .B(new_n1018), .C1(new_n1073), .C2(new_n1084), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n927), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n913), .ZN(new_n1090));
  OR3_X1    g665(.A1(new_n922), .A2(new_n715), .A3(new_n712), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n846), .A2(new_n914), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1090), .B1(new_n916), .B2(new_n915), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n921), .B(KEYINPUT46), .Z(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1096), .B(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n912), .A2(G1986), .A3(G290), .ZN(new_n1099));
  XOR2_X1   g674(.A(new_n1099), .B(KEYINPUT48), .Z(new_n1100));
  AOI211_X1 g675(.A(new_n1093), .B(new_n1098), .C1(new_n924), .C2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1089), .A2(new_n1101), .ZN(G329));
  assign    G231 = 1'b0;
  XNOR2_X1  g677(.A(new_n890), .B(KEYINPUT43), .ZN(new_n1104));
  NOR3_X1   g678(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1105));
  NAND2_X1  g679(.A1(new_n684), .A2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g680(.A(new_n1106), .B(KEYINPUT127), .ZN(new_n1107));
  AND3_X1   g681(.A1(new_n1104), .A2(new_n859), .A3(new_n1107), .ZN(G308));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n859), .A3(new_n1107), .ZN(G225));
endmodule


