

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n640, n641, n642, n643,
         n644, n645, n648, n649, n650, n651, n653, n654, n655, n656, n657,
         n658, n659, n660, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762;

  NAND2_X1 U367 ( .A1(n360), .A2(n359), .ZN(n358) );
  XNOR2_X1 U368 ( .A(n659), .B(n660), .ZN(n360) );
  INV_X1 U369 ( .A(n732), .ZN(n359) );
  INV_X1 U370 ( .A(n732), .ZN(n346) );
  INV_X1 U371 ( .A(n732), .ZN(n350) );
  INV_X1 U372 ( .A(n732), .ZN(n354) );
  NAND2_X1 U373 ( .A1(n572), .A2(n393), .ZN(n576) );
  XNOR2_X1 U374 ( .A(n560), .B(n559), .ZN(n577) );
  NAND2_X1 U375 ( .A1(n344), .A2(n435), .ZN(n434) );
  OR2_X2 U376 ( .A1(n573), .A2(n574), .ZN(n344) );
  XNOR2_X1 U377 ( .A(n645), .B(n348), .ZN(n347) );
  XNOR2_X1 U378 ( .A(n637), .B(n352), .ZN(n351) );
  XNOR2_X1 U379 ( .A(n651), .B(n356), .ZN(n355) );
  INV_X1 U380 ( .A(n345), .ZN(n357) );
  NAND2_X1 U381 ( .A1(n347), .A2(n346), .ZN(n345) );
  INV_X1 U382 ( .A(n644), .ZN(n348) );
  INV_X1 U383 ( .A(n349), .ZN(n640) );
  NAND2_X1 U384 ( .A1(n351), .A2(n350), .ZN(n349) );
  INV_X1 U385 ( .A(n636), .ZN(n352) );
  XNOR2_X2 U386 ( .A(n587), .B(n365), .ZN(n396) );
  INV_X1 U387 ( .A(n353), .ZN(n653) );
  NAND2_X1 U388 ( .A1(n355), .A2(n354), .ZN(n353) );
  INV_X1 U389 ( .A(n650), .ZN(n356) );
  INV_X2 U390 ( .A(KEYINPUT71), .ZN(n374) );
  XNOR2_X2 U391 ( .A(n750), .B(n445), .ZN(n468) );
  NAND2_X2 U392 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U393 ( .A(n357), .B(n648), .ZN(G57) );
  INV_X1 U394 ( .A(n358), .ZN(G66) );
  INV_X1 U395 ( .A(G146), .ZN(n445) );
  INV_X1 U396 ( .A(G953), .ZN(n755) );
  XNOR2_X1 U397 ( .A(n527), .B(n742), .ZN(n633) );
  NOR2_X2 U398 ( .A1(n409), .A2(n534), .ZN(n404) );
  AND2_X2 U399 ( .A1(n411), .A2(n410), .ZN(n409) );
  XNOR2_X2 U400 ( .A(n374), .B(G131), .ZN(n495) );
  NOR2_X1 U401 ( .A1(n398), .A2(n654), .ZN(n431) );
  XNOR2_X1 U402 ( .A(n376), .B(n375), .ZN(n570) );
  NAND2_X1 U403 ( .A1(n432), .A2(n430), .ZN(n429) );
  XNOR2_X1 U404 ( .A(n431), .B(KEYINPUT88), .ZN(n430) );
  OR2_X1 U405 ( .A1(n655), .A2(n578), .ZN(n433) );
  XNOR2_X1 U406 ( .A(n547), .B(KEYINPUT31), .ZN(n582) );
  XNOR2_X1 U407 ( .A(n592), .B(n593), .ZN(n760) );
  XNOR2_X1 U408 ( .A(KEYINPUT18), .B(KEYINPUT92), .ZN(n427) );
  OR2_X2 U409 ( .A1(n608), .A2(n540), .ZN(n380) );
  NOR2_X1 U410 ( .A1(n760), .A2(n762), .ZN(n417) );
  OR2_X1 U411 ( .A1(n531), .A2(n632), .ZN(n408) );
  XOR2_X1 U412 ( .A(G104), .B(G110), .Z(n740) );
  INV_X1 U413 ( .A(n598), .ZN(n395) );
  XNOR2_X1 U414 ( .A(n444), .B(n511), .ZN(n750) );
  XNOR2_X1 U415 ( .A(n443), .B(G143), .ZN(n517) );
  INV_X1 U416 ( .A(G128), .ZN(n443) );
  XNOR2_X1 U417 ( .A(n386), .B(n385), .ZN(n628) );
  INV_X1 U418 ( .A(KEYINPUT48), .ZN(n385) );
  XNOR2_X1 U419 ( .A(n420), .B(KEYINPUT113), .ZN(n686) );
  XNOR2_X1 U420 ( .A(n384), .B(n382), .ZN(n552) );
  XNOR2_X1 U421 ( .A(n504), .B(n383), .ZN(n382) );
  OR2_X1 U422 ( .A1(n649), .A2(G902), .ZN(n384) );
  INV_X1 U423 ( .A(G475), .ZN(n383) );
  XOR2_X1 U424 ( .A(G134), .B(n517), .Z(n511) );
  XNOR2_X1 U425 ( .A(G113), .B(G104), .ZN(n496) );
  XOR2_X1 U426 ( .A(KEYINPUT10), .B(G140), .Z(n480) );
  XNOR2_X1 U427 ( .A(G143), .B(G122), .ZN(n381) );
  XNOR2_X1 U428 ( .A(G107), .B(G140), .ZN(n462) );
  INV_X1 U429 ( .A(KEYINPUT80), .ZN(n463) );
  XNOR2_X1 U430 ( .A(G101), .B(KEYINPUT69), .ZN(n460) );
  XNOR2_X1 U431 ( .A(n390), .B(n595), .ZN(n625) );
  NAND2_X1 U432 ( .A1(n594), .A2(n688), .ZN(n390) );
  NOR2_X1 U433 ( .A1(n405), .A2(n404), .ZN(n403) );
  AND2_X1 U434 ( .A1(n407), .A2(n363), .ZN(n402) );
  INV_X1 U435 ( .A(KEYINPUT1), .ZN(n373) );
  INV_X1 U436 ( .A(KEYINPUT22), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n377) );
  NAND2_X1 U438 ( .A1(n369), .A2(n687), .ZN(n368) );
  NAND2_X1 U439 ( .A1(n582), .A2(KEYINPUT99), .ZN(n369) );
  XNOR2_X1 U440 ( .A(n612), .B(KEYINPUT76), .ZN(n415) );
  XOR2_X1 U441 ( .A(KEYINPUT69), .B(G101), .Z(n446) );
  XNOR2_X1 U442 ( .A(KEYINPUT3), .B(G119), .ZN(n448) );
  NAND2_X1 U443 ( .A1(n399), .A2(n361), .ZN(n405) );
  OR2_X1 U444 ( .A1(n408), .A2(n534), .ZN(n400) );
  INV_X1 U445 ( .A(KEYINPUT108), .ZN(n378) );
  NAND2_X1 U446 ( .A1(n531), .A2(n632), .ZN(n410) );
  XNOR2_X1 U447 ( .A(G119), .B(G128), .ZN(n472) );
  XNOR2_X1 U448 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n519) );
  AND2_X1 U449 ( .A1(n628), .A2(n364), .ZN(n422) );
  INV_X1 U450 ( .A(KEYINPUT2), .ZN(n423) );
  XNOR2_X1 U451 ( .A(n419), .B(n418), .ZN(n704) );
  INV_X1 U452 ( .A(KEYINPUT41), .ZN(n418) );
  NOR2_X1 U453 ( .A1(n546), .A2(n676), .ZN(n682) );
  AND2_X1 U454 ( .A1(n494), .A2(n541), .ZN(n594) );
  NOR2_X1 U455 ( .A1(n458), .A2(n584), .ZN(n494) );
  XNOR2_X1 U456 ( .A(n387), .B(KEYINPUT30), .ZN(n458) );
  NAND2_X1 U457 ( .A1(n587), .A2(n406), .ZN(n387) );
  XNOR2_X1 U458 ( .A(n513), .B(n512), .ZN(n728) );
  XNOR2_X1 U459 ( .A(n503), .B(n502), .ZN(n649) );
  XNOR2_X1 U460 ( .A(n466), .B(n465), .ZN(n467) );
  AND2_X1 U461 ( .A1(n638), .A2(G953), .ZN(n732) );
  XNOR2_X1 U462 ( .A(n389), .B(n596), .ZN(n762) );
  NOR2_X1 U463 ( .A1(n604), .A2(n603), .ZN(n724) );
  XNOR2_X1 U464 ( .A(n544), .B(KEYINPUT104), .ZN(n721) );
  NOR2_X1 U465 ( .A1(n553), .A2(n548), .ZN(n544) );
  XNOR2_X1 U466 ( .A(n397), .B(KEYINPUT109), .ZN(n654) );
  INV_X1 U467 ( .A(n604), .ZN(n561) );
  OR2_X1 U468 ( .A1(n406), .A2(n534), .ZN(n361) );
  AND2_X1 U469 ( .A1(n713), .A2(KEYINPUT99), .ZN(n362) );
  XNOR2_X1 U470 ( .A(n489), .B(n488), .ZN(n673) );
  INV_X1 U471 ( .A(n677), .ZN(n394) );
  NOR2_X1 U472 ( .A1(n689), .A2(KEYINPUT90), .ZN(n363) );
  AND2_X1 U473 ( .A1(n631), .A2(n630), .ZN(n364) );
  XOR2_X1 U474 ( .A(n556), .B(KEYINPUT6), .Z(n365) );
  XOR2_X1 U475 ( .A(KEYINPUT68), .B(KEYINPUT0), .Z(n366) );
  INV_X1 U476 ( .A(KEYINPUT90), .ZN(n534) );
  NAND2_X1 U477 ( .A1(n370), .A2(n367), .ZN(n391) );
  NOR2_X1 U478 ( .A1(n368), .A2(n362), .ZN(n367) );
  NAND2_X1 U479 ( .A1(n372), .A2(n371), .ZN(n370) );
  INV_X1 U480 ( .A(n713), .ZN(n371) );
  NOR2_X1 U481 ( .A1(n582), .A2(KEYINPUT99), .ZN(n372) );
  XNOR2_X2 U482 ( .A(n590), .B(n373), .ZN(n604) );
  XNOR2_X2 U483 ( .A(n469), .B(G469), .ZN(n590) );
  NAND2_X1 U484 ( .A1(n426), .A2(n377), .ZN(n376) );
  NAND2_X1 U485 ( .A1(n692), .A2(n672), .ZN(n379) );
  XNOR2_X2 U486 ( .A(n380), .B(n366), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n495), .B(n381), .ZN(n499) );
  NAND2_X1 U488 ( .A1(n412), .A2(n416), .ZN(n386) );
  XNOR2_X2 U489 ( .A(n388), .B(G472), .ZN(n587) );
  NAND2_X1 U490 ( .A1(n643), .A2(n484), .ZN(n388) );
  NAND2_X1 U491 ( .A1(n625), .A2(n721), .ZN(n389) );
  NAND2_X1 U492 ( .A1(n392), .A2(n391), .ZN(n398) );
  NAND2_X1 U493 ( .A1(n657), .A2(KEYINPUT44), .ZN(n392) );
  XNOR2_X2 U494 ( .A(n569), .B(KEYINPUT35), .ZN(n657) );
  AND2_X1 U495 ( .A1(n396), .A2(n393), .ZN(n557) );
  INV_X1 U496 ( .A(n673), .ZN(n393) );
  NOR2_X1 U497 ( .A1(n396), .A2(n394), .ZN(n562) );
  NOR2_X1 U498 ( .A1(n396), .A2(n395), .ZN(n599) );
  AND2_X1 U499 ( .A1(n396), .A2(n673), .ZN(n580) );
  XNOR2_X1 U500 ( .A(n555), .B(n554), .ZN(n692) );
  NAND2_X1 U501 ( .A1(n670), .A2(n632), .ZN(n421) );
  NAND2_X1 U502 ( .A1(n581), .A2(n580), .ZN(n397) );
  OR2_X1 U503 ( .A1(n633), .A2(n408), .ZN(n407) );
  OR2_X1 U504 ( .A1(n633), .A2(n400), .ZN(n399) );
  NAND2_X1 U505 ( .A1(n409), .A2(n407), .ZN(n533) );
  NAND2_X1 U506 ( .A1(n403), .A2(n401), .ZN(n600) );
  NAND2_X1 U507 ( .A1(n409), .A2(n402), .ZN(n401) );
  INV_X1 U508 ( .A(n689), .ZN(n406) );
  NAND2_X1 U509 ( .A1(n633), .A2(n531), .ZN(n411) );
  NOR2_X1 U510 ( .A1(n415), .A2(n413), .ZN(n412) );
  NAND2_X1 U511 ( .A1(n414), .A2(n438), .ZN(n413) );
  XNOR2_X1 U512 ( .A(n724), .B(KEYINPUT87), .ZN(n414) );
  XNOR2_X1 U513 ( .A(n417), .B(n597), .ZN(n416) );
  NAND2_X1 U514 ( .A1(n686), .A2(n692), .ZN(n419) );
  NAND2_X1 U515 ( .A1(n688), .A2(n406), .ZN(n420) );
  NOR2_X4 U516 ( .A1(n669), .A2(n421), .ZN(n658) );
  NAND2_X1 U517 ( .A1(n733), .A2(n422), .ZN(n670) );
  AND2_X2 U518 ( .A1(n424), .A2(n423), .ZN(n669) );
  NAND2_X1 U519 ( .A1(n733), .A2(n425), .ZN(n424) );
  INV_X1 U520 ( .A(n753), .ZN(n425) );
  XNOR2_X2 U521 ( .A(n429), .B(KEYINPUT45), .ZN(n733) );
  INV_X1 U522 ( .A(n426), .ZN(n543) );
  NAND2_X1 U523 ( .A1(n426), .A2(n682), .ZN(n547) );
  NAND2_X1 U524 ( .A1(n426), .A2(n702), .ZN(n565) );
  XNOR2_X1 U525 ( .A(n516), .B(n427), .ZN(n428) );
  XNOR2_X2 U526 ( .A(G146), .B(G125), .ZN(n516) );
  XNOR2_X1 U527 ( .A(n428), .B(n517), .ZN(n521) );
  NAND2_X1 U528 ( .A1(n434), .A2(n433), .ZN(n432) );
  INV_X1 U529 ( .A(KEYINPUT44), .ZN(n435) );
  AND2_X1 U530 ( .A1(KEYINPUT44), .A2(KEYINPUT70), .ZN(n437) );
  AND2_X1 U531 ( .A1(n616), .A2(n615), .ZN(n438) );
  INV_X1 U532 ( .A(KEYINPUT74), .ZN(n459) );
  XNOR2_X1 U533 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U534 ( .A(KEYINPUT107), .ZN(n554) );
  XNOR2_X1 U535 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U536 ( .A(KEYINPUT34), .ZN(n564) );
  XNOR2_X1 U537 ( .A(n479), .B(n478), .ZN(n481) );
  XNOR2_X1 U538 ( .A(n565), .B(n564), .ZN(n568) );
  XNOR2_X1 U539 ( .A(n481), .B(n749), .ZN(n482) );
  INV_X1 U540 ( .A(G902), .ZN(n484) );
  INV_X1 U541 ( .A(G237), .ZN(n439) );
  NAND2_X1 U542 ( .A1(n484), .A2(n439), .ZN(n529) );
  NAND2_X1 U543 ( .A1(n529), .A2(G214), .ZN(n440) );
  XNOR2_X1 U544 ( .A(n440), .B(KEYINPUT93), .ZN(n689) );
  XNOR2_X1 U545 ( .A(n495), .B(KEYINPUT72), .ZN(n442) );
  XOR2_X1 U546 ( .A(G137), .B(KEYINPUT4), .Z(n441) );
  XNOR2_X1 U547 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U548 ( .A(KEYINPUT5), .B(n446), .Z(n451) );
  NOR2_X1 U549 ( .A1(G953), .A2(G237), .ZN(n500) );
  NAND2_X1 U550 ( .A1(G210), .A2(n500), .ZN(n447) );
  XNOR2_X1 U551 ( .A(n447), .B(G116), .ZN(n449) );
  XNOR2_X1 U552 ( .A(n448), .B(G113), .ZN(n524) );
  XNOR2_X1 U553 ( .A(n449), .B(n524), .ZN(n450) );
  XNOR2_X1 U554 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U555 ( .A(n468), .B(n452), .ZN(n643) );
  NAND2_X1 U556 ( .A1(G234), .A2(G237), .ZN(n453) );
  XNOR2_X1 U557 ( .A(n453), .B(KEYINPUT14), .ZN(n454) );
  XNOR2_X1 U558 ( .A(KEYINPUT78), .B(n454), .ZN(n455) );
  NAND2_X1 U559 ( .A1(G952), .A2(n455), .ZN(n700) );
  NOR2_X1 U560 ( .A1(n700), .A2(G953), .ZN(n539) );
  NAND2_X1 U561 ( .A1(n455), .A2(G902), .ZN(n537) );
  OR2_X1 U562 ( .A1(n755), .A2(n537), .ZN(n456) );
  NOR2_X1 U563 ( .A1(G900), .A2(n456), .ZN(n457) );
  NOR2_X1 U564 ( .A1(n539), .A2(n457), .ZN(n584) );
  XNOR2_X1 U565 ( .A(n461), .B(n740), .ZN(n522) );
  XNOR2_X1 U566 ( .A(n522), .B(n462), .ZN(n466) );
  NAND2_X1 U567 ( .A1(G227), .A2(n755), .ZN(n464) );
  XNOR2_X1 U568 ( .A(n468), .B(n467), .ZN(n665) );
  NAND2_X1 U569 ( .A1(n665), .A2(n484), .ZN(n469) );
  XOR2_X1 U570 ( .A(KEYINPUT86), .B(KEYINPUT8), .Z(n471) );
  NAND2_X1 U571 ( .A1(G234), .A2(n755), .ZN(n470) );
  XNOR2_X1 U572 ( .A(n471), .B(n470), .ZN(n507) );
  NAND2_X1 U573 ( .A1(n507), .A2(G221), .ZN(n475) );
  XOR2_X1 U574 ( .A(G110), .B(G137), .Z(n473) );
  XNOR2_X1 U575 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U576 ( .A(n475), .B(n474), .ZN(n483) );
  XOR2_X1 U577 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n477) );
  XNOR2_X1 U578 ( .A(KEYINPUT24), .B(KEYINPUT85), .ZN(n476) );
  XNOR2_X1 U579 ( .A(n477), .B(n476), .ZN(n479) );
  XOR2_X1 U580 ( .A(KEYINPUT97), .B(KEYINPUT23), .Z(n478) );
  XNOR2_X1 U581 ( .A(n516), .B(n480), .ZN(n749) );
  XNOR2_X1 U582 ( .A(n483), .B(n482), .ZN(n660) );
  NAND2_X1 U583 ( .A1(n660), .A2(n484), .ZN(n489) );
  XNOR2_X1 U584 ( .A(G902), .B(KEYINPUT15), .ZN(n528) );
  NAND2_X1 U585 ( .A1(G234), .A2(n528), .ZN(n485) );
  XNOR2_X1 U586 ( .A(KEYINPUT20), .B(n485), .ZN(n490) );
  NAND2_X1 U587 ( .A1(G217), .A2(n490), .ZN(n487) );
  XNOR2_X1 U588 ( .A(KEYINPUT25), .B(KEYINPUT79), .ZN(n486) );
  XNOR2_X1 U589 ( .A(n487), .B(n486), .ZN(n488) );
  NAND2_X1 U590 ( .A1(G221), .A2(n490), .ZN(n491) );
  XOR2_X1 U591 ( .A(n491), .B(KEYINPUT21), .Z(n672) );
  AND2_X1 U592 ( .A1(n673), .A2(n672), .ZN(n677) );
  NAND2_X1 U593 ( .A1(n590), .A2(n677), .ZN(n493) );
  INV_X1 U594 ( .A(KEYINPUT98), .ZN(n492) );
  XNOR2_X1 U595 ( .A(n493), .B(n492), .ZN(n541) );
  XOR2_X1 U596 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n497) );
  XNOR2_X1 U597 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U598 ( .A(n499), .B(n498), .Z(n503) );
  NAND2_X1 U599 ( .A1(G214), .A2(n500), .ZN(n501) );
  XNOR2_X1 U600 ( .A(n749), .B(n501), .ZN(n502) );
  XNOR2_X1 U601 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n504) );
  XNOR2_X1 U602 ( .A(KEYINPUT103), .B(G478), .ZN(n515) );
  XOR2_X1 U603 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n506) );
  XNOR2_X1 U604 ( .A(KEYINPUT7), .B(KEYINPUT101), .ZN(n505) );
  XNOR2_X1 U605 ( .A(n506), .B(n505), .ZN(n509) );
  NAND2_X1 U606 ( .A1(G217), .A2(n507), .ZN(n508) );
  XNOR2_X1 U607 ( .A(n509), .B(n508), .ZN(n513) );
  XNOR2_X1 U608 ( .A(G122), .B(G116), .ZN(n510) );
  XNOR2_X1 U609 ( .A(n510), .B(G107), .ZN(n525) );
  XNOR2_X1 U610 ( .A(n511), .B(n525), .ZN(n512) );
  NOR2_X1 U611 ( .A1(G902), .A2(n728), .ZN(n514) );
  XNOR2_X1 U612 ( .A(n515), .B(n514), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n552), .A2(n553), .ZN(n566) );
  NAND2_X1 U614 ( .A1(n755), .A2(G224), .ZN(n518) );
  XNOR2_X1 U615 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U616 ( .A(n521), .B(n520), .ZN(n523) );
  XNOR2_X1 U617 ( .A(n523), .B(n522), .ZN(n527) );
  XNOR2_X1 U618 ( .A(n524), .B(KEYINPUT16), .ZN(n526) );
  XNOR2_X1 U619 ( .A(n526), .B(n525), .ZN(n742) );
  INV_X1 U620 ( .A(n528), .ZN(n632) );
  NAND2_X1 U621 ( .A1(n529), .A2(G210), .ZN(n530) );
  XNOR2_X1 U622 ( .A(n530), .B(KEYINPUT82), .ZN(n531) );
  NOR2_X1 U623 ( .A1(n566), .A2(n533), .ZN(n532) );
  NAND2_X1 U624 ( .A1(n594), .A2(n532), .ZN(n615) );
  XNOR2_X1 U625 ( .A(n615), .B(G143), .ZN(G45) );
  XNOR2_X1 U626 ( .A(KEYINPUT67), .B(KEYINPUT19), .ZN(n535) );
  XNOR2_X1 U627 ( .A(n600), .B(n535), .ZN(n608) );
  NOR2_X1 U628 ( .A1(G898), .A2(n755), .ZN(n536) );
  XOR2_X1 U629 ( .A(KEYINPUT94), .B(n536), .Z(n746) );
  NOR2_X1 U630 ( .A1(n746), .A2(n537), .ZN(n538) );
  NOR2_X1 U631 ( .A1(n539), .A2(n538), .ZN(n540) );
  INV_X1 U632 ( .A(n587), .ZN(n676) );
  NAND2_X1 U633 ( .A1(n541), .A2(n676), .ZN(n542) );
  NOR2_X1 U634 ( .A1(n543), .A2(n542), .ZN(n713) );
  INV_X1 U635 ( .A(n552), .ZN(n548) );
  NAND2_X1 U636 ( .A1(n713), .A2(n721), .ZN(n545) );
  XNOR2_X1 U637 ( .A(n545), .B(G104), .ZN(G6) );
  OR2_X1 U638 ( .A1(n604), .A2(n394), .ZN(n546) );
  NAND2_X1 U639 ( .A1(n548), .A2(n553), .ZN(n549) );
  XNOR2_X1 U640 ( .A(n549), .B(KEYINPUT105), .ZN(n717) );
  NAND2_X1 U641 ( .A1(n582), .A2(n717), .ZN(n550) );
  XNOR2_X1 U642 ( .A(n550), .B(G116), .ZN(G18) );
  NAND2_X1 U643 ( .A1(n582), .A2(n721), .ZN(n551) );
  XNOR2_X1 U644 ( .A(n551), .B(G113), .ZN(G15) );
  NOR2_X1 U645 ( .A1(n553), .A2(n552), .ZN(n555) );
  INV_X1 U646 ( .A(KEYINPUT106), .ZN(n556) );
  AND2_X1 U647 ( .A1(n561), .A2(n557), .ZN(n558) );
  AND2_X1 U648 ( .A1(n570), .A2(n558), .ZN(n560) );
  XNOR2_X1 U649 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n559) );
  XNOR2_X1 U650 ( .A(n577), .B(G119), .ZN(G21) );
  XNOR2_X2 U651 ( .A(n563), .B(KEYINPUT33), .ZN(n702) );
  XNOR2_X1 U652 ( .A(n566), .B(KEYINPUT81), .ZN(n567) );
  NAND2_X1 U653 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U654 ( .A(n657), .B(KEYINPUT70), .ZN(n574) );
  NAND2_X1 U655 ( .A1(n570), .A2(n604), .ZN(n579) );
  NOR2_X1 U656 ( .A1(n579), .A2(n587), .ZN(n571) );
  XNOR2_X1 U657 ( .A(n571), .B(KEYINPUT66), .ZN(n572) );
  NAND2_X1 U658 ( .A1(n576), .A2(n577), .ZN(n573) );
  INV_X1 U659 ( .A(n576), .ZN(n655) );
  NAND2_X1 U660 ( .A1(n577), .A2(n437), .ZN(n578) );
  INV_X1 U661 ( .A(n579), .ZN(n581) );
  OR2_X1 U662 ( .A1(n721), .A2(n717), .ZN(n687) );
  XOR2_X1 U663 ( .A(KEYINPUT114), .B(KEYINPUT42), .Z(n593) );
  XOR2_X1 U664 ( .A(KEYINPUT112), .B(KEYINPUT28), .Z(n589) );
  INV_X1 U665 ( .A(n672), .ZN(n583) );
  NOR2_X1 U666 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U667 ( .A(n585), .B(KEYINPUT73), .ZN(n586) );
  NOR2_X1 U668 ( .A1(n673), .A2(n586), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n598), .A2(n587), .ZN(n588) );
  XNOR2_X1 U670 ( .A(n589), .B(n588), .ZN(n591) );
  NAND2_X1 U671 ( .A1(n591), .A2(n590), .ZN(n607) );
  XNOR2_X1 U672 ( .A(n533), .B(KEYINPUT38), .ZN(n688) );
  OR2_X1 U673 ( .A1(n607), .A2(n704), .ZN(n592) );
  INV_X1 U674 ( .A(KEYINPUT40), .ZN(n596) );
  XOR2_X1 U675 ( .A(KEYINPUT75), .B(KEYINPUT39), .Z(n595) );
  XNOR2_X1 U676 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n721), .A2(n599), .ZN(n617) );
  NOR2_X1 U678 ( .A1(n617), .A2(n600), .ZN(n602) );
  XNOR2_X1 U679 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n601) );
  XNOR2_X1 U680 ( .A(n602), .B(n601), .ZN(n603) );
  INV_X1 U681 ( .A(n687), .ZN(n605) );
  NOR2_X1 U682 ( .A1(n605), .A2(KEYINPUT47), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n606), .B(KEYINPUT77), .ZN(n611) );
  INV_X1 U684 ( .A(n607), .ZN(n610) );
  INV_X1 U685 ( .A(n608), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n613) );
  NOR2_X1 U687 ( .A1(n611), .A2(n613), .ZN(n612) );
  INV_X1 U688 ( .A(n613), .ZN(n722) );
  NAND2_X1 U689 ( .A1(n722), .A2(n687), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n614), .A2(KEYINPUT47), .ZN(n616) );
  INV_X1 U691 ( .A(n617), .ZN(n619) );
  NOR2_X1 U692 ( .A1(n561), .A2(n689), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U694 ( .A(KEYINPUT43), .B(n620), .ZN(n621) );
  XNOR2_X1 U695 ( .A(KEYINPUT110), .B(n621), .ZN(n622) );
  AND2_X1 U696 ( .A1(n622), .A2(n533), .ZN(n624) );
  INV_X1 U697 ( .A(KEYINPUT111), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n624), .B(n623), .ZN(n759) );
  NAND2_X1 U699 ( .A1(n625), .A2(n717), .ZN(n726) );
  INV_X1 U700 ( .A(n726), .ZN(n626) );
  NOR2_X1 U701 ( .A1(n759), .A2(n626), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n753) );
  INV_X1 U703 ( .A(n759), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n726), .A2(KEYINPUT2), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n629), .B(KEYINPUT83), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n658), .A2(G210), .ZN(n637) );
  XNOR2_X1 U707 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n634) );
  XNOR2_X1 U708 ( .A(n634), .B(KEYINPUT55), .ZN(n635) );
  XNOR2_X1 U709 ( .A(n633), .B(n635), .ZN(n636) );
  INV_X1 U710 ( .A(G952), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n640), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U712 ( .A(KEYINPUT63), .ZN(n648) );
  NAND2_X1 U713 ( .A1(n658), .A2(G472), .ZN(n645) );
  XNOR2_X1 U714 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n641), .B(KEYINPUT62), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n643), .B(n642), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n658), .A2(G475), .ZN(n651) );
  XOR2_X1 U718 ( .A(KEYINPUT59), .B(n649), .Z(n650) );
  XNOR2_X1 U719 ( .A(n653), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U720 ( .A(G101), .B(n654), .Z(G3) );
  INV_X1 U721 ( .A(n655), .ZN(n656) );
  XNOR2_X1 U722 ( .A(n656), .B(G110), .ZN(G12) );
  XOR2_X1 U723 ( .A(n657), .B(G122), .Z(G24) );
  BUF_X2 U724 ( .A(n658), .Z(n727) );
  NAND2_X1 U725 ( .A1(n727), .A2(G217), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n727), .A2(G469), .ZN(n667) );
  XOR2_X1 U727 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n663) );
  XNOR2_X1 U728 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n662) );
  XNOR2_X1 U729 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U731 ( .A(n667), .B(n666), .ZN(n668) );
  NOR2_X1 U732 ( .A1(n668), .A2(n732), .ZN(G54) );
  XOR2_X1 U733 ( .A(KEYINPUT84), .B(n669), .Z(n671) );
  NAND2_X1 U734 ( .A1(n671), .A2(n670), .ZN(n710) );
  NOR2_X1 U735 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U736 ( .A(n674), .B(KEYINPUT49), .ZN(n675) );
  NAND2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n680) );
  NOR2_X1 U738 ( .A1(n677), .A2(n561), .ZN(n678) );
  XNOR2_X1 U739 ( .A(n678), .B(KEYINPUT50), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U741 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U742 ( .A(n683), .B(KEYINPUT51), .ZN(n685) );
  INV_X1 U743 ( .A(n704), .ZN(n684) );
  NAND2_X1 U744 ( .A1(n685), .A2(n684), .ZN(n698) );
  NAND2_X1 U745 ( .A1(n687), .A2(n686), .ZN(n695) );
  INV_X1 U746 ( .A(n688), .ZN(n690) );
  NAND2_X1 U747 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U748 ( .A(KEYINPUT118), .B(n691), .ZN(n693) );
  NAND2_X1 U749 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U750 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U751 ( .A1(n696), .A2(n702), .ZN(n697) );
  NAND2_X1 U752 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U753 ( .A(KEYINPUT52), .B(n699), .Z(n701) );
  NOR2_X1 U754 ( .A1(n701), .A2(n700), .ZN(n708) );
  INV_X1 U755 ( .A(n702), .ZN(n703) );
  NOR2_X1 U756 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U757 ( .A(n705), .B(KEYINPUT119), .ZN(n706) );
  NAND2_X1 U758 ( .A1(n706), .A2(n755), .ZN(n707) );
  NOR2_X1 U759 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U760 ( .A1(n710), .A2(n709), .ZN(n712) );
  XOR2_X1 U761 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n711) );
  XNOR2_X1 U762 ( .A(n712), .B(n711), .ZN(G75) );
  NAND2_X1 U763 ( .A1(n713), .A2(n717), .ZN(n715) );
  XOR2_X1 U764 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n714) );
  XNOR2_X1 U765 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U766 ( .A(G107), .B(n716), .ZN(G9) );
  XOR2_X1 U767 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n719) );
  NAND2_X1 U768 ( .A1(n722), .A2(n717), .ZN(n718) );
  XNOR2_X1 U769 ( .A(n719), .B(n718), .ZN(n720) );
  XOR2_X1 U770 ( .A(G128), .B(n720), .Z(G30) );
  NAND2_X1 U771 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U772 ( .A(n723), .B(G146), .ZN(G48) );
  XNOR2_X1 U773 ( .A(G125), .B(n724), .ZN(n725) );
  XNOR2_X1 U774 ( .A(n725), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U775 ( .A(G134), .B(n726), .ZN(G36) );
  NAND2_X1 U776 ( .A1(n727), .A2(G478), .ZN(n730) );
  XOR2_X1 U777 ( .A(n728), .B(KEYINPUT123), .Z(n729) );
  XNOR2_X1 U778 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U779 ( .A1(n732), .A2(n731), .ZN(G63) );
  BUF_X1 U780 ( .A(n733), .Z(n734) );
  NAND2_X1 U781 ( .A1(n734), .A2(n755), .ZN(n739) );
  NAND2_X1 U782 ( .A1(G224), .A2(G953), .ZN(n735) );
  XNOR2_X1 U783 ( .A(n735), .B(KEYINPUT124), .ZN(n736) );
  XNOR2_X1 U784 ( .A(KEYINPUT61), .B(n736), .ZN(n737) );
  NAND2_X1 U785 ( .A1(G898), .A2(n737), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n739), .A2(n738), .ZN(n748) );
  XOR2_X1 U787 ( .A(G101), .B(KEYINPUT126), .Z(n744) );
  XNOR2_X1 U788 ( .A(KEYINPUT125), .B(n740), .ZN(n741) );
  XNOR2_X1 U789 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U790 ( .A(n744), .B(n743), .ZN(n745) );
  NAND2_X1 U791 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U792 ( .A(n748), .B(n747), .Z(G69) );
  XOR2_X1 U793 ( .A(n750), .B(n749), .Z(n754) );
  XNOR2_X1 U794 ( .A(G227), .B(n754), .ZN(n751) );
  NAND2_X1 U795 ( .A1(G900), .A2(n751), .ZN(n752) );
  NAND2_X1 U796 ( .A1(n752), .A2(G953), .ZN(n758) );
  XNOR2_X1 U797 ( .A(n754), .B(n753), .ZN(n756) );
  NAND2_X1 U798 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U799 ( .A1(n758), .A2(n757), .ZN(G72) );
  XOR2_X1 U800 ( .A(G140), .B(n759), .Z(G42) );
  XNOR2_X1 U801 ( .A(G137), .B(n760), .ZN(n761) );
  XNOR2_X1 U802 ( .A(n761), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U803 ( .A(G131), .B(n762), .Z(G33) );
endmodule

