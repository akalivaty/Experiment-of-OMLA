//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(G58), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n203), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  INV_X1    g0026(.A(G116), .ZN(new_n227));
  INV_X1    g0027(.A(G270), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n206), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n209), .B(new_n218), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT67), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g0050(.A1(KEYINPUT67), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n250), .A2(new_n215), .A3(new_n251), .A4(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(G20), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G50), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n250), .A2(new_n215), .A3(new_n251), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n216), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n216), .A2(new_n262), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G50), .A2(G58), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n216), .B1(new_n265), .B2(new_n211), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n258), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n257), .B(new_n267), .C1(G50), .C2(new_n253), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT9), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT66), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(G222), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(G223), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n280), .B1(new_n220), .B2(new_n278), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT64), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n215), .B1(KEYINPUT65), .B2(new_n289), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n289), .A2(KEYINPUT65), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n288), .A2(G274), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n286), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n290), .B2(new_n291), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n294), .B1(G226), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n285), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n269), .B(new_n270), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(G200), .B2(new_n298), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n305), .B(new_n268), .C1(G179), .C2(new_n298), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n296), .A2(G238), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n293), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n275), .A2(KEYINPUT66), .A3(new_n276), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n273), .B1(new_n271), .B2(new_n272), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(G232), .A4(G1698), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(G226), .A4(new_n279), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G97), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n284), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT13), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(KEYINPUT70), .ZN(new_n320));
  XOR2_X1   g0120(.A(new_n318), .B(new_n320), .Z(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G179), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n319), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n310), .A2(KEYINPUT13), .A3(new_n317), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(G169), .A3(new_n324), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(KEYINPUT14), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(KEYINPUT14), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n322), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n211), .A2(G20), .ZN(new_n329));
  INV_X1    g0129(.A(G50), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n329), .B1(new_n260), .B2(new_n220), .C1(new_n330), .C2(new_n263), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT11), .B1(new_n331), .B2(new_n258), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n253), .A2(G68), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT12), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n255), .A2(G68), .A3(new_n256), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n321), .A2(G190), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n323), .A2(G200), .A3(new_n324), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n255), .A2(G77), .A3(new_n256), .ZN(new_n344));
  XOR2_X1   g0144(.A(new_n344), .B(KEYINPUT68), .Z(new_n345));
  NAND2_X1  g0145(.A1(G20), .A2(G77), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT15), .B(G87), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n346), .B1(new_n259), .B2(new_n263), .C1(new_n260), .C2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n253), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n348), .A2(new_n258), .B1(new_n220), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n278), .A2(G232), .A3(new_n279), .ZN(new_n352));
  INV_X1    g0152(.A(G238), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n352), .B1(new_n203), .B2(new_n278), .C1(new_n281), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n284), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n294), .B1(G244), .B2(new_n296), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n351), .B1(new_n358), .B2(G169), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n357), .A2(G179), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G200), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n345), .B(new_n350), .C1(new_n357), .C2(new_n299), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n308), .A2(new_n340), .A3(new_n343), .A4(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n258), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT72), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n210), .B2(new_n211), .ZN(new_n370));
  NAND3_X1  g0170(.A1(KEYINPUT72), .A2(G58), .A3(G68), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n370), .A2(new_n212), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G159), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n372), .A2(new_n216), .B1(new_n373), .B2(new_n263), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n271), .A2(new_n272), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n275), .A2(new_n216), .A3(new_n276), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT71), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n378), .B1(new_n377), .B2(new_n379), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n376), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n374), .B1(new_n382), .B2(G68), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n368), .B1(new_n383), .B2(KEYINPUT16), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n216), .B1(new_n274), .B2(new_n277), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(KEYINPUT73), .A3(new_n379), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT73), .ZN(new_n387));
  AOI21_X1  g0187(.A(G20), .B1(new_n311), .B2(new_n312), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n387), .B1(new_n388), .B2(KEYINPUT7), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n389), .A3(new_n376), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n374), .B1(new_n390), .B2(G68), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n384), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n296), .A2(G232), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n293), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n282), .A2(G1698), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n271), .B2(new_n272), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G87), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(G226), .A2(G1698), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n271), .B2(new_n272), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT74), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(KEYINPUT74), .B(new_n399), .C1(new_n271), .C2(new_n272), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n398), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT75), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n284), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n275), .A2(new_n276), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n395), .B1(G33), .B2(G87), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT74), .B1(new_n407), .B2(new_n399), .ZN(new_n409));
  INV_X1    g0209(.A(new_n403), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n408), .B(new_n405), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n299), .B(new_n394), .C1(new_n406), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n293), .A2(new_n393), .ZN(new_n414));
  INV_X1    g0214(.A(new_n284), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(KEYINPUT75), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n414), .B1(new_n417), .B2(new_n411), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n413), .B1(G200), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n259), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n256), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n421), .A2(new_n254), .B1(new_n253), .B2(new_n420), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n392), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT76), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT76), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n392), .A2(new_n419), .A3(new_n426), .A4(new_n423), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(KEYINPUT17), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n392), .A2(new_n419), .A3(new_n429), .A4(new_n423), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n430), .A2(KEYINPUT77), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n392), .A2(new_n423), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n418), .A2(G179), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n304), .B2(new_n418), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(KEYINPUT18), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT18), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n433), .B2(new_n435), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT77), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n425), .A2(new_n441), .A3(KEYINPUT17), .A4(new_n427), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n432), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n367), .A2(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(KEYINPUT78), .A2(G97), .ZN(new_n445));
  NAND2_X1  g0245(.A1(KEYINPUT78), .A2(G97), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n262), .ZN(new_n448));
  AOI21_X1  g0248(.A(G20), .B1(G33), .B2(G283), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n227), .A2(G20), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n450), .A2(KEYINPUT20), .A3(new_n258), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT86), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT20), .ZN(new_n455));
  AOI21_X1  g0255(.A(G33), .B1(new_n445), .B2(new_n446), .ZN(new_n456));
  INV_X1    g0256(.A(new_n449), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n451), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n455), .B1(new_n458), .B2(new_n368), .ZN(new_n459));
  INV_X1    g0259(.A(new_n458), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n460), .A2(KEYINPUT86), .A3(KEYINPUT20), .A4(new_n258), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n454), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n253), .A2(G116), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n463), .B(KEYINPUT85), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n254), .B1(new_n252), .B2(G33), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(G116), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT87), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n462), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n467), .B1(new_n462), .B2(new_n466), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n222), .A2(G1698), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n407), .B(new_n472), .C1(G257), .C2(G1698), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G303), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n311), .B2(new_n312), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT83), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT83), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n478), .B(new_n473), .C1(new_n278), .C2(new_n475), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n284), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G45), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G1), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n292), .A2(G274), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n482), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n292), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n486), .B2(new_n228), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT82), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT82), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n484), .B(new_n489), .C1(new_n486), .C2(new_n228), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n480), .A2(KEYINPUT84), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT84), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n477), .A2(new_n479), .A3(new_n492), .A4(new_n284), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(G179), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n480), .A2(KEYINPUT84), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n488), .A2(new_n490), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(KEYINPUT21), .A3(G169), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n471), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n462), .A2(new_n466), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n468), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n497), .A2(new_n299), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n362), .B1(new_n491), .B2(new_n493), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  XOR2_X1   g0305(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n304), .B1(new_n491), .B2(new_n493), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n502), .B2(new_n508), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n499), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n407), .A2(new_n216), .A3(G87), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT22), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT89), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(KEYINPUT89), .A3(KEYINPUT22), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n225), .A2(KEYINPUT22), .A3(G20), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n514), .A2(new_n515), .B1(new_n278), .B2(new_n516), .ZN(new_n517));
  OR3_X1    g0317(.A1(new_n216), .A2(KEYINPUT23), .A3(G107), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n216), .A2(G33), .A3(G116), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT90), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT23), .B1(new_n216), .B2(G107), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n520), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT24), .B1(new_n517), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n278), .A2(new_n516), .ZN(new_n527));
  INV_X1    g0327(.A(new_n515), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT89), .B1(new_n511), .B2(KEYINPUT22), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n524), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n258), .ZN(new_n534));
  NOR2_X1   g0334(.A1(G250), .A2(G1698), .ZN(new_n535));
  INV_X1    g0335(.A(G257), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n536), .B2(G1698), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(new_n407), .B1(G33), .B2(G294), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n486), .A2(new_n222), .B1(new_n538), .B2(new_n415), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n362), .B1(new_n540), .B2(new_n484), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n484), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n541), .B1(new_n543), .B2(G190), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n349), .A2(new_n203), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n545), .B(KEYINPUT25), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n465), .B2(G107), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n534), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n253), .A2(G97), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n465), .B2(G97), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n447), .A2(KEYINPUT6), .A3(new_n203), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT6), .B1(new_n204), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n554), .A2(new_n216), .B1(new_n220), .B2(new_n263), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n390), .B2(G107), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n550), .B1(new_n556), .B2(new_n368), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n484), .B1(new_n486), .B2(new_n536), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT4), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n560), .A2(new_n221), .A3(G1698), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n278), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n407), .A2(G244), .A3(new_n279), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n563), .A2(new_n560), .B1(G33), .B2(G283), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n559), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n558), .B1(new_n565), .B2(new_n284), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(G169), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n284), .ZN(new_n569));
  INV_X1    g0369(.A(new_n558), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n557), .B(new_n568), .C1(G179), .C2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(KEYINPUT79), .A3(G200), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT79), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n566), .B2(new_n362), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n566), .A2(G190), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n548), .B(new_n572), .C1(new_n557), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n542), .A2(new_n304), .ZN(new_n579));
  INV_X1    g0379(.A(G179), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n543), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n368), .B1(new_n526), .B2(new_n532), .ZN(new_n582));
  INV_X1    g0382(.A(new_n547), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n579), .B(new_n581), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n292), .A2(G274), .A3(new_n482), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT80), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n292), .A2(KEYINPUT80), .A3(G274), .A4(new_n482), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n292), .B(G250), .C1(G1), .C2(new_n481), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n221), .A2(G1698), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(G238), .B2(G1698), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n591), .A2(new_n375), .B1(new_n262), .B2(new_n227), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n284), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G169), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n580), .B2(new_n594), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT81), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n445), .A2(new_n446), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(new_n225), .A3(new_n203), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT19), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n216), .B1(new_n315), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n375), .A2(G20), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n600), .A2(new_n602), .B1(new_n603), .B2(G68), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n601), .B1(new_n599), .B2(new_n260), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n368), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n349), .B2(new_n347), .ZN(new_n607));
  INV_X1    g0407(.A(new_n465), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n607), .B1(new_n347), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n595), .B(KEYINPUT81), .C1(new_n580), .C2(new_n594), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n598), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n594), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G190), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n594), .A2(G200), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n465), .A2(G87), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n607), .A2(new_n613), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n584), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n578), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n444), .A2(new_n510), .A3(new_n618), .ZN(G372));
  NAND2_X1  g0419(.A1(new_n609), .A2(new_n596), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n616), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n578), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n502), .A2(new_n508), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n506), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n498), .A2(new_n494), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n624), .B(new_n584), .C1(new_n625), .C2(new_n471), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n622), .A2(new_n626), .B1(new_n596), .B2(new_n609), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n611), .A2(new_n616), .ZN(new_n628));
  INV_X1    g0428(.A(new_n572), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT26), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n572), .A2(KEYINPUT91), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT91), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n567), .B1(new_n580), .B2(new_n566), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(new_n634), .B2(new_n557), .ZN(new_n635));
  OR3_X1    g0435(.A1(new_n632), .A2(new_n635), .A3(new_n621), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n627), .B(new_n631), .C1(KEYINPUT26), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n444), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n341), .A2(new_n338), .A3(new_n342), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n359), .A2(new_n360), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n340), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n641), .A2(new_n432), .A3(new_n442), .ZN(new_n642));
  INV_X1    g0442(.A(new_n440), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n303), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n306), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT92), .ZN(G369));
  INV_X1    g0447(.A(new_n499), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n624), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n252), .A2(new_n216), .A3(G13), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT93), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g0454(.A(KEYINPUT94), .B(G343), .Z(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n471), .A2(new_n657), .ZN(new_n658));
  MUX2_X1   g0458(.A(new_n510), .B(new_n649), .S(new_n658), .Z(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n581), .A2(new_n579), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n534), .B2(new_n547), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n656), .B1(new_n582), .B2(new_n583), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n548), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n584), .A2(new_n656), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n665), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n656), .B1(new_n648), .B2(new_n624), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(G399));
  NOR2_X1   g0471(.A1(new_n600), .A2(G116), .ZN(new_n672));
  INV_X1    g0472(.A(new_n207), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(G1), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n213), .B2(new_n675), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n637), .A2(new_n657), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(KEYINPUT29), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n499), .A2(new_n509), .A3(new_n662), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n577), .A2(new_n557), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n620), .A2(new_n616), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n572), .A4(new_n548), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n620), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n628), .A2(new_n686), .A3(new_n629), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n632), .A2(new_n635), .A3(new_n621), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n657), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(KEYINPUT29), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n680), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT96), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT95), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n612), .A2(new_n695), .A3(new_n540), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT95), .B1(new_n594), .B2(new_n539), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n566), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n693), .B(new_n694), .C1(new_n699), .C2(new_n494), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n543), .A2(new_n566), .A3(G179), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n497), .A3(new_n594), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n497), .A2(new_n580), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n693), .A2(new_n694), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n566), .A3(new_n704), .A4(new_n698), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n700), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n656), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT98), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(KEYINPUT98), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT97), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n711), .A2(KEYINPUT97), .A3(new_n714), .A4(new_n712), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n510), .A2(new_n618), .A3(new_n657), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n692), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n678), .B1(new_n721), .B2(G1), .ZN(G364));
  AND2_X1   g0522(.A1(new_n216), .A2(G13), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n252), .B1(new_n723), .B2(G45), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n674), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n660), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(G330), .B2(new_n659), .ZN(new_n728));
  INV_X1    g0528(.A(new_n726), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n216), .A2(new_n580), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n731), .A2(new_n299), .A3(G200), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n362), .A2(G190), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT33), .B(G317), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n732), .A2(G322), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT102), .Z(new_n738));
  NOR2_X1   g0538(.A1(new_n299), .A2(new_n362), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n730), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n216), .A2(G179), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G190), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n741), .A2(G326), .B1(new_n745), .B2(G329), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n730), .A2(new_n743), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G311), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n739), .A2(new_n742), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT101), .Z(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G303), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n733), .A2(new_n742), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT100), .Z(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G283), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n299), .A2(G179), .A3(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n216), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n278), .B1(G294), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n750), .A2(new_n753), .A3(new_n756), .A4(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n732), .A2(G58), .B1(G68), .B2(new_n735), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n762), .B(new_n278), .C1(new_n202), .C2(new_n758), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n755), .A2(G107), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n744), .A2(new_n373), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT32), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n740), .A2(new_n330), .B1(new_n751), .B2(new_n225), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(G77), .B2(new_n748), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n764), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n738), .A2(new_n761), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n215), .B1(G20), .B2(new_n304), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n729), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n771), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n278), .A2(new_n207), .ZN(new_n778));
  INV_X1    g0578(.A(G355), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n778), .A2(new_n779), .B1(G116), .B2(new_n207), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT99), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n214), .A2(new_n481), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n673), .A2(new_n407), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n783), .B(new_n784), .C1(new_n243), .C2(new_n481), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n780), .A2(new_n781), .ZN(new_n786));
  AND3_X1   g0586(.A1(new_n782), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n772), .B1(new_n777), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT103), .ZN(new_n789));
  INV_X1    g0589(.A(new_n775), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n659), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n728), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  NAND2_X1  g0593(.A1(new_n351), .A2(new_n656), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT106), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n351), .A2(KEYINPUT106), .A3(new_n656), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n365), .A2(new_n798), .B1(new_n360), .B2(new_n359), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n361), .A2(new_n657), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n679), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n801), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n631), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n657), .B(new_n803), .C1(new_n804), .C2(new_n685), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n726), .B1(new_n720), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n720), .B2(new_n806), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G150), .A2(new_n735), .B1(new_n748), .B2(G159), .ZN(new_n809));
  INV_X1    g0609(.A(G137), .ZN(new_n810));
  INV_X1    g0610(.A(G143), .ZN(new_n811));
  INV_X1    g0611(.A(new_n732), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n809), .B1(new_n810), .B2(new_n740), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT105), .B(KEYINPUT34), .Z(new_n814));
  XNOR2_X1  g0614(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n752), .A2(G50), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n755), .A2(G68), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n759), .A2(G58), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n375), .B1(new_n745), .B2(G132), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G283), .A2(new_n735), .B1(new_n745), .B2(G311), .ZN(new_n821));
  INV_X1    g0621(.A(new_n278), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n821), .B(new_n822), .C1(new_n202), .C2(new_n758), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n812), .A2(new_n824), .B1(new_n740), .B2(new_n475), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G116), .B2(new_n748), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n752), .A2(G107), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n755), .A2(G87), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n815), .A2(new_n820), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n771), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n771), .A2(new_n773), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT104), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n729), .B1(new_n834), .B2(new_n220), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n831), .B(new_n835), .C1(new_n803), .C2(new_n774), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n808), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G384));
  INV_X1    g0638(.A(new_n554), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n839), .A2(KEYINPUT35), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(KEYINPUT35), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n840), .A2(G116), .A3(new_n217), .A4(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT36), .Z(new_n843));
  NAND4_X1  g0643(.A1(new_n214), .A2(G77), .A3(new_n370), .A4(new_n371), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n330), .A2(G68), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n252), .B(G13), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n384), .B1(KEYINPUT16), .B2(new_n383), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n654), .B1(new_n848), .B2(new_n423), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n443), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n423), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n434), .B(new_n654), .C1(new_n304), .C2(new_n418), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n425), .A2(new_n427), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT107), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT107), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n854), .A2(new_n857), .A3(KEYINPUT37), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n425), .A2(new_n427), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT16), .ZN(new_n860));
  INV_X1    g0660(.A(new_n376), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n385), .A2(new_n379), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n862), .B2(new_n387), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n211), .B1(new_n863), .B2(new_n386), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n860), .B1(new_n864), .B2(new_n374), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n422), .B1(new_n865), .B2(new_n384), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n418), .A2(new_n304), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(G179), .B2(new_n418), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT108), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT108), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n433), .A2(new_n435), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n866), .A2(new_n654), .ZN(new_n873));
  XOR2_X1   g0673(.A(KEYINPUT109), .B(KEYINPUT37), .Z(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n859), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n856), .A2(new_n858), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n850), .A2(new_n878), .A3(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n436), .A2(new_n424), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n875), .B1(new_n880), .B2(new_n873), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n443), .A2(new_n873), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n879), .B1(KEYINPUT38), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n850), .A2(new_n878), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n340), .A2(new_n656), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n805), .A2(new_n800), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n339), .B(new_n656), .C1(new_n639), .C2(new_n328), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n339), .A2(new_n656), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n340), .A2(new_n343), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n850), .A2(new_n878), .A3(KEYINPUT38), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n850), .B2(new_n878), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n654), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n898), .A2(new_n901), .B1(new_n440), .B2(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n891), .A2(new_n892), .B1(new_n903), .B2(KEYINPUT110), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n903), .A2(KEYINPUT110), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n444), .B1(new_n680), .B2(new_n691), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n645), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n906), .B(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n718), .A2(new_n709), .A3(new_n714), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n444), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT111), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n801), .B1(new_n894), .B2(new_n896), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n443), .A2(new_n873), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n877), .A2(new_n881), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT38), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n914), .B1(new_n899), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n888), .A2(new_n879), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n910), .A2(new_n920), .A3(new_n913), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n918), .A2(KEYINPUT40), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n912), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n912), .A2(new_n922), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(G330), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n909), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n252), .B2(new_n723), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n909), .A2(new_n925), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n847), .B1(new_n927), .B2(new_n928), .ZN(G367));
  NAND2_X1  g0729(.A1(new_n239), .A2(new_n784), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(new_n776), .C1(new_n207), .C2(new_n347), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT116), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n729), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n931), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n812), .A2(new_n261), .B1(new_n740), .B2(new_n811), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n734), .A2(new_n373), .B1(new_n744), .B2(new_n810), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n278), .B1(new_n211), .B2(new_n758), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n754), .ZN(new_n939));
  AOI22_X1  g0739(.A1(G50), .A2(new_n748), .B1(new_n939), .B2(G77), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n938), .B(new_n940), .C1(new_n210), .C2(new_n751), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n734), .A2(new_n824), .ZN(new_n942));
  INV_X1    g0742(.A(G283), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n375), .B1(new_n747), .B2(new_n943), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n942), .B(new_n944), .C1(G311), .C2(new_n741), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n751), .A2(new_n227), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n945), .B1(KEYINPUT46), .B2(new_n946), .C1(new_n203), .C2(new_n758), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n752), .A2(KEYINPUT46), .A3(G116), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n732), .A2(G303), .B1(G317), .B2(new_n745), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(new_n599), .C2(new_n754), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n941), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT47), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n934), .B1(new_n952), .B2(new_n771), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n607), .A2(new_n615), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n656), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n683), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n620), .A2(new_n955), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n953), .B1(new_n959), .B2(new_n790), .ZN(new_n960));
  XOR2_X1   g0760(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT113), .Z(new_n964));
  NAND2_X1  g0764(.A1(new_n557), .A2(new_n656), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n682), .A2(new_n572), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n572), .B2(new_n657), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(new_n666), .A3(new_n669), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n572), .B1(new_n966), .B2(new_n584), .ZN(new_n969));
  AOI22_X1  g0769(.A1(KEYINPUT42), .A2(new_n968), .B1(new_n969), .B2(new_n657), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(KEYINPUT42), .B2(new_n968), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n964), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n962), .B1(new_n973), .B2(KEYINPUT114), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT114), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n972), .A2(new_n975), .A3(new_n962), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n660), .A2(new_n666), .A3(new_n967), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT115), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n977), .A2(new_n978), .B1(KEYINPUT115), .B2(new_n979), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n666), .B(new_n669), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n660), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n721), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n670), .A2(new_n668), .A3(new_n967), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT45), .Z(new_n988));
  AOI21_X1  g0788(.A(new_n967), .B1(new_n670), .B2(new_n668), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n660), .A3(new_n666), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(new_n667), .A3(new_n990), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n721), .B1(new_n986), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n674), .B(KEYINPUT41), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n725), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n960), .B1(new_n983), .B2(new_n998), .ZN(G387));
  OAI21_X1  g0799(.A(new_n784), .B1(new_n236), .B2(new_n481), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n672), .B2(new_n778), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n259), .A2(G50), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT50), .ZN(new_n1003));
  AOI21_X1  g0803(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1003), .A2(new_n672), .A3(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1001), .A2(new_n1005), .B1(new_n203), .B2(new_n673), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n726), .B1(new_n1006), .B2(new_n777), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n732), .A2(G50), .B1(new_n420), .B2(new_n735), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n220), .B2(new_n751), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G97), .B2(new_n755), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n740), .A2(new_n373), .B1(new_n744), .B2(new_n261), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n375), .B(new_n1011), .C1(G68), .C2(new_n748), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(new_n347), .C2(new_n758), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n407), .B1(new_n745), .B2(G326), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n758), .A2(new_n943), .B1(new_n751), .B2(new_n824), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n732), .A2(G317), .B1(new_n741), .B2(G322), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G303), .A2(new_n748), .B1(new_n735), .B2(G311), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT48), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1015), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n1019), .B2(new_n1018), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT49), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1014), .B1(new_n227), .B2(new_n754), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1013), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(KEYINPUT117), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n771), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n1025), .B2(KEYINPUT117), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1007), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n666), .B2(new_n790), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT118), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n985), .B2(new_n725), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n986), .A2(new_n674), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n721), .A2(new_n985), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(G393));
  INV_X1    g0835(.A(new_n994), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n721), .A2(new_n985), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n675), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n986), .A2(new_n994), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(KEYINPUT121), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT121), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1039), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n674), .B1(new_n986), .B2(new_n994), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1036), .A2(new_n725), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n732), .A2(G159), .B1(new_n741), .B2(G150), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT119), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1048), .A2(KEYINPUT51), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(KEYINPUT51), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n330), .A2(new_n734), .B1(new_n751), .B2(new_n211), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n407), .B1(new_n747), .B2(new_n259), .C1(new_n758), .C2(new_n220), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(G143), .C2(new_n745), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1049), .A2(new_n828), .A3(new_n1050), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n732), .A2(G311), .B1(new_n741), .B2(G317), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT52), .Z(new_n1056));
  NOR2_X1   g0856(.A1(new_n751), .A2(new_n943), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n824), .A2(new_n747), .B1(new_n734), .B2(new_n475), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(G322), .C2(new_n745), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n278), .B1(G116), .B2(new_n759), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1056), .A2(new_n764), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1027), .B1(new_n1054), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n246), .A2(new_n784), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n777), .B1(new_n673), .B2(new_n447), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n729), .B(new_n1062), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT120), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n967), .B2(new_n790), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1046), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1045), .A2(new_n1069), .ZN(G390));
  NAND4_X1  g0870(.A1(new_n719), .A2(G330), .A3(new_n803), .A4(new_n897), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n657), .B(new_n799), .C1(new_n685), .C2(new_n689), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n800), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n910), .A2(G330), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n803), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n897), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1071), .A2(new_n1078), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1074), .A2(new_n801), .A3(new_n1077), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n719), .A2(G330), .A3(new_n803), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1080), .B1(new_n1081), .B2(new_n1077), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n893), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1079), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n444), .A2(new_n1075), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n907), .A2(new_n645), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT122), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n907), .A2(KEYINPUT122), .A3(new_n645), .A4(new_n1085), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1084), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1073), .A2(new_n897), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n892), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n1092), .A3(new_n883), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n892), .B1(new_n893), .B2(new_n897), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1071), .C1(new_n891), .C2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n885), .A2(new_n889), .B1(new_n898), .B2(new_n1092), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1093), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1080), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n675), .B1(new_n1090), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n1099), .B2(new_n1090), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n890), .A2(new_n773), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n726), .B1(new_n833), .B2(new_n420), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n752), .A2(G87), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n745), .A2(G294), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G283), .A2(new_n741), .B1(new_n748), .B2(new_n447), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1105), .A2(new_n817), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n732), .A2(G116), .B1(G107), .B2(new_n735), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1109), .B(new_n822), .C1(new_n220), .C2(new_n758), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n751), .A2(new_n261), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT53), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G128), .A2(new_n741), .B1(new_n748), .B2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n939), .A2(G50), .B1(new_n745), .B2(G125), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n732), .A2(G132), .B1(G137), .B2(new_n735), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n278), .C1(new_n373), .C2(new_n758), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1108), .A2(new_n1110), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1104), .B1(new_n1120), .B2(new_n771), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1102), .A2(new_n725), .B1(new_n1103), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1101), .A2(new_n1122), .ZN(G378));
  INV_X1    g0923(.A(KEYINPUT125), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n902), .A2(new_n268), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n307), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n307), .A2(new_n1128), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1126), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1131), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(new_n1129), .A3(new_n1125), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(G330), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1136), .B1(new_n922), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n920), .B1(new_n883), .B2(new_n914), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n910), .A2(new_n913), .A3(new_n920), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n888), .B2(new_n879), .ZN(new_n1141));
  OAI211_X1 g0941(.A(G330), .B(new_n1135), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT124), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1124), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(KEYINPUT124), .B(KEYINPUT125), .C1(new_n1138), .C2(new_n1142), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n906), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1142), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n921), .B1(new_n899), .B2(new_n900), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n910), .A2(new_n913), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n915), .A2(new_n916), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n887), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n1152), .B2(new_n879), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1149), .B1(new_n1153), .B2(new_n920), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1135), .B1(new_n1154), .B2(G330), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1144), .B1(new_n1148), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT125), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n906), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1143), .A2(new_n1144), .A3(new_n1124), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1147), .A2(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1084), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n1099), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT57), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(KEYINPUT57), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1148), .A2(new_n1155), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n906), .B(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n674), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1136), .A2(new_n773), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n726), .B1(new_n833), .B2(G50), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n407), .A2(G41), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n740), .A2(new_n227), .B1(new_n751), .B2(new_n220), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(G97), .C2(new_n735), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n744), .A2(new_n943), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n747), .A2(new_n347), .B1(new_n754), .B2(new_n210), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(G107), .C2(new_n732), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1175), .B(new_n1178), .C1(new_n211), .C2(new_n758), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT58), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1173), .B(new_n330), .C1(G33), .C2(G41), .ZN(new_n1181));
  INV_X1    g0981(.A(G125), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n740), .A2(new_n1182), .B1(new_n747), .B2(new_n810), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n732), .A2(G128), .ZN(new_n1184));
  INV_X1    g0984(.A(G132), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1184), .B1(new_n1185), .B2(new_n734), .C1(new_n751), .C2(new_n1113), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1183), .B(new_n1186), .C1(G150), .C2(new_n759), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n939), .A2(G159), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G33), .B(G41), .C1(new_n745), .C2(G124), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1180), .B(new_n1181), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT123), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1027), .B1(new_n1194), .B2(KEYINPUT123), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1172), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1171), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1161), .B2(new_n725), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1170), .A2(new_n1200), .ZN(G375));
  NAND2_X1  g1001(.A1(new_n1077), .A2(new_n773), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n812), .A2(new_n810), .B1(new_n734), .B2(new_n1113), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n375), .B(new_n1203), .C1(G58), .C2(new_n939), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n759), .A2(G50), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n752), .A2(G159), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n740), .A2(new_n1185), .B1(new_n747), .B2(new_n261), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G128), .B2(new_n745), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n740), .A2(new_n824), .B1(new_n734), .B2(new_n227), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G107), .B2(new_n748), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT126), .Z(new_n1212));
  OAI22_X1  g1012(.A1(new_n812), .A2(new_n943), .B1(new_n744), .B2(new_n475), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n758), .A2(new_n347), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1213), .A2(new_n278), .A3(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G97), .A2(new_n752), .B1(new_n755), .B2(G77), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1212), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1027), .B1(new_n1209), .B2(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n729), .B(new_n1218), .C1(new_n211), .C2(new_n834), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1084), .A2(new_n725), .B1(new_n1202), .B2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1162), .A2(new_n1084), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1090), .A2(new_n997), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1220), .B1(new_n1221), .B2(new_n1222), .ZN(G381));
  INV_X1    g1023(.A(new_n960), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n995), .A2(new_n997), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n724), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n981), .A2(new_n982), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1224), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1068), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OR4_X1    g1031(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1231), .ZN(G407));
  AND2_X1   g1032(.A1(new_n1101), .A2(new_n1122), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n655), .A2(G213), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G375), .C2(new_n1236), .ZN(G409));
  OAI211_X1 g1037(.A(G378), .B(new_n1200), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1102), .B2(new_n1084), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n996), .B(new_n1240), .C1(new_n1147), .C2(new_n1160), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1198), .B1(new_n1168), .B2(new_n724), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1233), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1238), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1234), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1235), .A2(G2897), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n675), .B1(new_n1162), .B2(new_n1084), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1162), .A2(KEYINPUT60), .A3(new_n1084), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT60), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1163), .B2(new_n1239), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1248), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1252), .A2(G384), .A3(new_n1220), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G384), .B1(new_n1252), .B2(new_n1220), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1247), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1252), .A2(new_n1220), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n837), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1252), .A2(G384), .A3(new_n1220), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n1246), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT61), .B1(new_n1245), .B2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT127), .B1(G390), .B2(new_n1228), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(G393), .B(G396), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G387), .A2(new_n1229), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G390), .A2(new_n1228), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1262), .A2(new_n1266), .A3(new_n1265), .A4(new_n1263), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1235), .B1(new_n1238), .B2(new_n1243), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1272), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1261), .B(new_n1270), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1271), .A2(new_n1277), .A3(new_n1273), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1271), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1277), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1278), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1276), .B1(new_n1283), .B2(new_n1270), .ZN(G405));
  NAND2_X1  g1084(.A1(G375), .A2(new_n1233), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1270), .A2(new_n1285), .A3(new_n1238), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G378), .B1(new_n1170), .B2(new_n1200), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1238), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1269), .B(new_n1268), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1286), .A2(new_n1273), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1273), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(G402));
endmodule


