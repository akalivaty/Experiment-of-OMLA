//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  INV_X1    g0026(.A(new_n201), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT65), .Z(new_n229));
  AND2_X1   g0029(.A1(KEYINPUT64), .A2(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(KEYINPUT64), .A2(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n212), .A2(new_n226), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT66), .B(G50), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G58), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(KEYINPUT8), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT69), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT67), .B(G58), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT68), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT8), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n260), .B2(KEYINPUT8), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n232), .A2(G33), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n256), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n233), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(new_n206), .B2(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G50), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n270), .B(new_n272), .C1(G50), .C2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  OAI211_X1 g0078(.A(G1), .B(G13), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n279), .A3(G274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n275), .ZN(new_n281));
  INV_X1    g0081(.A(G226), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n277), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G222), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(new_n285), .B2(new_n286), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G223), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n289), .B1(new_n220), .B2(new_n287), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n283), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n274), .B(new_n297), .C1(G169), .C2(new_n295), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(G190), .B2(new_n295), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n274), .A2(KEYINPUT9), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n274), .A2(KEYINPUT9), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n299), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OR2_X1    g0108(.A1(KEYINPUT64), .A2(G20), .ZN(new_n309));
  NAND2_X1  g0109(.A1(KEYINPUT64), .A2(G20), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT7), .B1(new_n311), .B2(new_n287), .ZN(new_n312));
  AND2_X1   g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NOR2_X1   g0113(.A1(KEYINPUT3), .A2(G33), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT7), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n207), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(G68), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n227), .B1(new_n260), .B2(new_n214), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT73), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n207), .A2(new_n277), .ZN(new_n323));
  INV_X1    g0123(.A(G159), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n255), .A2(KEYINPUT73), .A3(G159), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n321), .A2(G20), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n312), .A2(KEYINPUT74), .A3(G68), .A4(new_n317), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n320), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT16), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT7), .B1(new_n287), .B2(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n232), .A2(new_n315), .A3(new_n316), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(G68), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n327), .A2(KEYINPUT16), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n269), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n265), .A2(new_n273), .ZN(new_n338));
  INV_X1    g0138(.A(new_n271), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n264), .A2(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n331), .A2(new_n337), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n292), .A2(new_n288), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n282), .A2(G1698), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n344), .C1(new_n313), .C2(new_n314), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT75), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G87), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n346), .B1(new_n345), .B2(new_n347), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n294), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n280), .B1(new_n281), .B2(new_n239), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n342), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(new_n352), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n353), .B1(new_n355), .B2(G179), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT18), .B1(new_n341), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n356), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT18), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n338), .A2(new_n340), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n325), .A2(new_n326), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT67), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G58), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n201), .B1(new_n365), .B2(G68), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n361), .B1(new_n366), .B2(new_n207), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n319), .B2(new_n318), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT16), .B1(new_n368), .B2(new_n328), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n360), .B1(new_n369), .B2(new_n336), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n358), .A2(new_n359), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n357), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT76), .ZN(new_n373));
  INV_X1    g0173(.A(G190), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n280), .B(new_n374), .C1(new_n281), .C2(new_n239), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n345), .A2(new_n347), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT75), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n375), .B1(new_n379), .B2(new_n294), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n373), .A2(new_n380), .B1(new_n354), .B2(new_n300), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n279), .B1(new_n377), .B2(new_n378), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT76), .B1(new_n382), .B2(new_n375), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT77), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n300), .B1(new_n382), .B2(new_n351), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n350), .A2(new_n373), .A3(new_n374), .A4(new_n352), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n383), .A2(new_n385), .A3(KEYINPUT77), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n341), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT77), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n370), .B1(new_n395), .B2(new_n387), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT17), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(KEYINPUT78), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n372), .B1(new_n392), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n214), .A2(G20), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n402), .B1(new_n202), .B2(new_n323), .C1(new_n266), .C2(new_n220), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n269), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT71), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n405), .A2(KEYINPUT11), .ZN(new_n406));
  INV_X1    g0206(.A(G13), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(G1), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI211_X1 g0209(.A(new_n402), .B(new_n409), .C1(KEYINPUT72), .C2(KEYINPUT12), .ZN(new_n410));
  OR3_X1    g0210(.A1(new_n410), .A2(KEYINPUT72), .A3(KEYINPUT12), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n410), .B1(KEYINPUT72), .B2(KEYINPUT12), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(new_n412), .C1(new_n214), .C2(new_n339), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n405), .B2(KEYINPUT11), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n406), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n287), .A2(G232), .A3(G1698), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n287), .A2(G226), .A3(new_n288), .ZN(new_n417));
  INV_X1    g0217(.A(G97), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n416), .B(new_n417), .C1(new_n277), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n294), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n276), .A2(new_n279), .A3(G274), .ZN(new_n421));
  INV_X1    g0221(.A(new_n281), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(G238), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT13), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(G169), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n296), .B2(new_n425), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n425), .B2(G169), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n415), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n415), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n425), .A2(G200), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n431), .B(new_n432), .C1(new_n374), .C2(new_n425), .ZN(new_n433));
  INV_X1    g0233(.A(new_n269), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT8), .B(G58), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(new_n255), .B1(new_n311), .B2(G77), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT15), .B(G87), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(G33), .A3(new_n232), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n434), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n273), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n220), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n339), .B2(new_n220), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n287), .A2(G232), .A3(new_n288), .ZN(new_n446));
  OAI221_X1 g0246(.A(new_n446), .B1(new_n222), .B2(new_n287), .C1(new_n291), .C2(new_n215), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n294), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n421), .B1(G244), .B2(new_n422), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n445), .B1(new_n451), .B2(new_n342), .ZN(new_n452));
  AND4_X1   g0252(.A1(KEYINPUT70), .A2(new_n448), .A3(new_n296), .A4(new_n449), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT70), .B1(new_n450), .B2(new_n296), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n445), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n451), .B2(G200), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n374), .B2(new_n451), .ZN(new_n458));
  AND4_X1   g0258(.A1(new_n430), .A2(new_n433), .A3(new_n455), .A4(new_n458), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n308), .A2(new_n401), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(G97), .A2(G107), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n216), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT19), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n463), .A2(new_n277), .A3(new_n418), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n464), .B2(new_n311), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n309), .A2(G33), .A3(G97), .A4(new_n310), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n463), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n287), .A2(new_n232), .A3(G68), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n469), .A2(new_n269), .B1(new_n442), .B2(new_n438), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n206), .A2(G33), .ZN(new_n471));
  AND4_X1   g0271(.A1(new_n233), .A2(new_n273), .A3(new_n268), .A4(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n470), .B1(new_n438), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n217), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n279), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n279), .A2(G274), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n206), .A2(G45), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(G238), .B(new_n288), .C1(new_n313), .C2(new_n314), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n287), .A2(KEYINPUT81), .A3(G238), .A4(new_n288), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n287), .A2(G244), .A3(G1698), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G116), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n481), .B1(new_n488), .B2(new_n294), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n296), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n474), .B(new_n490), .C1(G169), .C2(new_n489), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n290), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT80), .ZN(new_n493));
  OAI211_X1 g0293(.A(G244), .B(new_n288), .C1(new_n313), .C2(new_n314), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT4), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n221), .B1(new_n285), .B2(new_n286), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n288), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n494), .A2(new_n495), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n492), .A2(new_n496), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n294), .ZN(new_n501));
  OR2_X1    g0301(.A1(KEYINPUT5), .A2(G41), .ZN(new_n502));
  NAND2_X1  g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n480), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n294), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G257), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n503), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(new_n279), .A3(G274), .A4(new_n476), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n501), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G200), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n316), .B1(new_n232), .B2(new_n315), .ZN(new_n511));
  NOR4_X1   g0311(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT7), .A4(G20), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n511), .A2(new_n512), .A3(new_n222), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n222), .A2(KEYINPUT6), .A3(G97), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT6), .ZN(new_n516));
  XNOR2_X1  g0316(.A(G97), .B(G107), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI22_X1  g0318(.A1(new_n518), .A2(new_n232), .B1(new_n220), .B2(new_n323), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n269), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT79), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n312), .A2(G107), .A3(new_n317), .ZN(new_n523));
  AND2_X1   g0323(.A1(G97), .A2(G107), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n516), .B1(new_n524), .B2(new_n461), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n514), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(new_n311), .B1(G77), .B2(new_n255), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n434), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT79), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n273), .A2(G97), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n472), .B2(G97), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n500), .A2(new_n294), .B1(G257), .B2(new_n505), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(G190), .A3(new_n508), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n510), .A2(new_n530), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n528), .A2(KEYINPUT79), .ZN(new_n536));
  AOI211_X1 g0336(.A(new_n521), .B(new_n434), .C1(new_n523), .C2(new_n527), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n533), .A2(new_n296), .A3(new_n508), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n509), .A2(new_n342), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n488), .A2(new_n294), .ZN(new_n542));
  INV_X1    g0342(.A(new_n481), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(G190), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n472), .A2(G87), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n470), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n542), .A2(new_n543), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n489), .A2(KEYINPUT82), .A3(G190), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n546), .A2(new_n548), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  AND4_X1   g0352(.A1(new_n491), .A2(new_n535), .A3(new_n541), .A4(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT21), .ZN(new_n554));
  OAI211_X1 g0354(.A(G257), .B(new_n288), .C1(new_n313), .C2(new_n314), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT83), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n287), .A2(KEYINPUT83), .A3(G257), .A4(new_n288), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(G264), .B(G1698), .C1(new_n313), .C2(new_n314), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n285), .A2(G303), .A3(new_n286), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n279), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n503), .ZN(new_n565));
  NOR2_X1   g0365(.A1(KEYINPUT5), .A2(G41), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n476), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n279), .ZN(new_n568));
  INV_X1    g0368(.A(G270), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n508), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(G116), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n442), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n472), .A2(G116), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n277), .A2(G97), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G283), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n309), .A2(new_n575), .A3(new_n310), .A4(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n268), .A2(new_n233), .B1(G20), .B2(new_n572), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n577), .A2(KEYINPUT20), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT20), .B1(new_n577), .B2(new_n578), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n573), .B(new_n574), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G169), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n554), .B1(new_n571), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n570), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n562), .B1(new_n557), .B2(new_n558), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n585), .B2(new_n279), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n586), .A2(KEYINPUT21), .A3(G169), .A4(new_n581), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n571), .A2(G179), .A3(new_n581), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n217), .A2(new_n288), .ZN(new_n590));
  INV_X1    g0390(.A(G257), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G1698), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n590), .B(new_n592), .C1(new_n313), .C2(new_n314), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G33), .A2(G294), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT84), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(KEYINPUT84), .A3(new_n594), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n294), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n508), .B1(new_n568), .B2(new_n223), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(G169), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n279), .B1(new_n595), .B2(new_n596), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n600), .B1(new_n603), .B2(new_n598), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(new_n296), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n287), .A2(new_n232), .A3(G87), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT22), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT22), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n287), .A2(new_n232), .A3(new_n608), .A4(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(KEYINPUT23), .A2(G107), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(G20), .ZN(new_n613));
  NOR2_X1   g0413(.A1(KEYINPUT23), .A2(G107), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n311), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT24), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT24), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n610), .A2(new_n618), .A3(new_n615), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n434), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT25), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n273), .B2(G107), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n273), .A2(new_n621), .A3(G107), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n622), .A2(new_n624), .B1(new_n472), .B2(G107), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n605), .B1(new_n620), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n599), .A2(new_n601), .A3(new_n374), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n628), .B(KEYINPUT85), .C1(G200), .C2(new_n604), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n610), .A2(new_n618), .A3(new_n615), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n618), .B1(new_n610), .B2(new_n615), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n269), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT85), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n604), .A2(new_n633), .A3(new_n374), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n629), .A2(new_n632), .A3(new_n625), .A4(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n581), .B1(new_n586), .B2(G200), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n374), .B2(new_n586), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n589), .A2(new_n627), .A3(new_n635), .A4(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n460), .A2(new_n553), .A3(new_n638), .ZN(G372));
  INV_X1    g0439(.A(new_n455), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n433), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n430), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n400), .B1(new_n396), .B2(new_n390), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n372), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n306), .A2(new_n307), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n299), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n552), .A2(new_n491), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(KEYINPUT26), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n552), .A2(new_n491), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n541), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n649), .A2(new_n541), .A3(new_n535), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n604), .A2(new_n296), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(G169), .B2(new_n604), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n632), .B2(new_n625), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n635), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n491), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n460), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n648), .A2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n232), .A2(new_n666), .A3(new_n408), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G213), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT86), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n666), .B1(new_n232), .B2(new_n408), .ZN(new_n670));
  OR3_X1    g0470(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n668), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n581), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n589), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n637), .ZN(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n675), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n632), .B2(new_n625), .ZN(new_n683));
  INV_X1    g0483(.A(new_n635), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n627), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n659), .A2(new_n682), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n589), .A2(new_n675), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n686), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n689), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n210), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n462), .A2(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n229), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n696), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n663), .A2(new_n682), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT90), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT90), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(new_n706), .A3(new_n703), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n649), .A2(KEYINPUT91), .A3(KEYINPUT26), .A4(new_n650), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n708), .B(new_n491), .C1(new_n656), .C2(new_n661), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT91), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n651), .A2(new_n710), .A3(new_n654), .ZN(new_n711));
  OAI211_X1 g0511(.A(KEYINPUT29), .B(new_n682), .C1(new_n709), .C2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n705), .A2(new_n707), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n553), .A2(new_n638), .A3(new_n682), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n599), .A2(new_n601), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n549), .A2(new_n586), .A3(new_n296), .A4(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n509), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n564), .A2(new_n296), .A3(new_n570), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(new_n489), .A3(new_n533), .A4(new_n604), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT87), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT30), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n549), .A2(new_n715), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(KEYINPUT87), .A3(new_n533), .A4(new_n719), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n718), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n682), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n714), .B1(KEYINPUT31), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n675), .A2(KEYINPUT31), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n604), .A2(new_n501), .A3(new_n489), .A4(new_n506), .ZN(new_n732));
  INV_X1    g0532(.A(new_n564), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(G179), .A3(new_n584), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n721), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n724), .A3(new_n726), .ZN(new_n736));
  INV_X1    g0536(.A(new_n718), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n727), .B1(new_n738), .B2(KEYINPUT88), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT88), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n725), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n731), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(G330), .B1(new_n730), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT89), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(KEYINPUT89), .B(G330), .C1(new_n730), .C2(new_n742), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n713), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n701), .B1(new_n750), .B2(G1), .ZN(G364));
  NOR2_X1   g0551(.A1(new_n311), .A2(new_n407), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G45), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G1), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n695), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT92), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n233), .B1(G20), .B2(new_n342), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n311), .A2(new_n296), .A3(new_n374), .A4(new_n300), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT94), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(KEYINPUT94), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT95), .B(KEYINPUT32), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n765), .A2(G159), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n232), .A2(new_n296), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G190), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n374), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n220), .A2(new_n770), .B1(new_n772), .B2(new_n260), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n300), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n311), .A2(new_n374), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n222), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n774), .A2(G20), .A3(G190), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n374), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n232), .A2(new_n778), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n287), .B1(new_n216), .B2(new_n777), .C1(new_n779), .C2(new_n418), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n773), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n766), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n764), .B2(new_n324), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n768), .A2(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n374), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(G190), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G50), .A2(new_n785), .B1(new_n786), .B2(G68), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n767), .A2(new_n781), .A3(new_n783), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n765), .A2(G329), .ZN(new_n789));
  INV_X1    g0589(.A(G303), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n315), .B1(new_n777), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G294), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n779), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n770), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n791), .B(new_n793), .C1(new_n794), .C2(G311), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G326), .A2(new_n785), .B1(new_n786), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n772), .ZN(new_n798));
  INV_X1    g0598(.A(new_n775), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n798), .A2(G322), .B1(G283), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n789), .A2(new_n795), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n759), .B1(new_n788), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n758), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n694), .A2(new_n315), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(G355), .B1(new_n572), .B2(new_n694), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n210), .A2(new_n315), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT93), .Z(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(G45), .B2(new_n699), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n250), .A2(new_n475), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n808), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n757), .B(new_n802), .C1(new_n806), .C2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT96), .Z(new_n815));
  INV_X1    g0615(.A(new_n678), .ZN(new_n816));
  INV_X1    g0616(.A(new_n805), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n755), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n678), .A2(new_n679), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n681), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  NAND2_X1  g0623(.A1(new_n675), .A2(new_n456), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n455), .A2(new_n458), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n455), .B2(new_n824), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n702), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n682), .B(new_n826), .C1(new_n655), .C2(new_n662), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n819), .B1(new_n831), .B2(new_n747), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n747), .B2(new_n831), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n827), .A2(new_n803), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n758), .A2(new_n803), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n756), .B1(G77), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n785), .A2(G303), .B1(new_n794), .B2(G116), .ZN(new_n838));
  INV_X1    g0638(.A(G283), .ZN(new_n839));
  INV_X1    g0639(.A(new_n786), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT97), .Z(new_n842));
  INV_X1    g0642(.A(new_n777), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n287), .B1(new_n843), .B2(G107), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n844), .B1(new_n418), .B2(new_n779), .C1(new_n772), .C2(new_n792), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n775), .A2(new_n216), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n765), .B2(G311), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT98), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G159), .A2(new_n794), .B1(new_n798), .B2(G143), .ZN(new_n850));
  INV_X1    g0650(.A(G150), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n840), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G137), .B2(new_n785), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT34), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n775), .A2(new_n214), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G50), .B2(new_n843), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT99), .Z(new_n857));
  INV_X1    g0657(.A(new_n779), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n315), .B1(new_n858), .B2(new_n365), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n857), .B(new_n859), .C1(new_n860), .C2(new_n764), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n846), .A2(new_n849), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n837), .B1(new_n862), .B2(new_n758), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n833), .B1(new_n834), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  OAI211_X1 g0665(.A(new_n229), .B(G77), .C1(new_n214), .C2(new_n260), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n202), .A2(G68), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n206), .B(G13), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n526), .A2(KEYINPUT35), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n526), .A2(KEYINPUT35), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n869), .A2(G116), .A3(new_n234), .A4(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(KEYINPUT100), .B(KEYINPUT36), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n356), .A2(new_n673), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT16), .B1(new_n327), .B2(new_n334), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n360), .B1(new_n336), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n878), .B2(new_n396), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(new_n673), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n370), .B1(new_n358), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n389), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n877), .A2(new_n881), .ZN(new_n885));
  OAI211_X1 g0685(.A(KEYINPUT38), .B(new_n884), .C1(new_n401), .C2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT101), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n396), .A2(new_n390), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n398), .B(new_n370), .C1(new_n395), .C2(new_n387), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n645), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n885), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(KEYINPUT101), .A3(KEYINPUT38), .A4(new_n884), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n884), .B1(new_n401), .B2(new_n885), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n888), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT39), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n370), .A2(new_n881), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n643), .B2(new_n645), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n341), .B1(new_n356), .B2(new_n673), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n902), .B2(new_n396), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n903), .A2(new_n883), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n896), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(new_n886), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n899), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n428), .A2(new_n429), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n415), .A3(new_n682), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n640), .A2(new_n682), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n829), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n415), .A2(new_n675), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n433), .A2(new_n430), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n415), .A3(new_n675), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n920), .A2(new_n898), .B1(new_n372), .B2(new_n673), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n912), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n705), .A2(new_n460), .A3(new_n707), .A4(new_n712), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n648), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n922), .B(new_n924), .Z(new_n925));
  NAND2_X1  g0725(.A1(new_n905), .A2(new_n886), .ZN(new_n926));
  OR2_X1    g0726(.A1(KEYINPUT102), .A2(KEYINPUT31), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n729), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n729), .A2(new_n927), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n714), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n827), .B1(new_n916), .B2(new_n917), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n926), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT40), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT40), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n898), .A2(new_n934), .A3(new_n930), .A4(new_n931), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n936), .A2(new_n460), .A3(new_n930), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n460), .B2(new_n930), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n937), .A2(new_n938), .A3(new_n679), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n925), .A2(new_n939), .B1(new_n206), .B2(new_n752), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n925), .A2(new_n939), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n874), .B1(new_n940), .B2(new_n941), .ZN(G367));
  NAND2_X1  g0742(.A1(new_n810), .A2(new_n245), .ZN(new_n943));
  INV_X1    g0743(.A(new_n806), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n694), .B2(new_n439), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n757), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n682), .A2(new_n548), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n649), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n491), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n765), .A2(G137), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n287), .B1(new_n777), .B2(new_n260), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n779), .A2(new_n214), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n951), .B(new_n952), .C1(new_n794), .C2(G50), .ZN(new_n953));
  AOI22_X1  g0753(.A1(G143), .A2(new_n785), .B1(new_n786), .B2(G159), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n775), .A2(new_n220), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n798), .B2(G150), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n950), .A2(new_n953), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n799), .A2(G97), .ZN(new_n958));
  INV_X1    g0758(.A(G317), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n315), .B(new_n958), .C1(new_n764), .C2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT104), .Z(new_n961));
  OAI22_X1  g0761(.A1(new_n839), .A2(new_n770), .B1(new_n772), .B2(new_n790), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n843), .A2(KEYINPUT46), .A3(G116), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT46), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n777), .B2(new_n572), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n963), .B(new_n965), .C1(new_n222), .C2(new_n779), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n962), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(G311), .ZN(new_n968));
  INV_X1    g0768(.A(new_n785), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n967), .B1(new_n792), .B2(new_n840), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n957), .B1(new_n961), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT47), .Z(new_n972));
  OAI221_X1 g0772(.A(new_n946), .B1(new_n817), .B2(new_n949), .C1(new_n972), .C2(new_n759), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n538), .A2(new_n675), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n535), .A2(new_n541), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n541), .B2(new_n682), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n691), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT42), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n541), .B1(new_n975), .B2(new_n627), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT103), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(KEYINPUT103), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n682), .A3(new_n982), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n979), .A2(new_n983), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n689), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n977), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n986), .B(new_n988), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n692), .A2(new_n977), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n692), .A2(new_n977), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n993), .A2(KEYINPUT45), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(KEYINPUT45), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n689), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n992), .B(new_n987), .C1(new_n994), .C2(new_n995), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n687), .B(new_n690), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(new_n680), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n750), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n750), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n695), .B(KEYINPUT41), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n754), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n973), .B1(new_n989), .B2(new_n1006), .ZN(G387));
  INV_X1    g0807(.A(new_n807), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n1008), .A2(new_n697), .B1(G107), .B2(new_n210), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n435), .A2(G50), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n697), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT106), .B1(new_n810), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n242), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1015), .B1(G45), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n810), .A2(KEYINPUT106), .A3(new_n1014), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1009), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n756), .B1(new_n1019), .B2(new_n944), .ZN(new_n1020));
  INV_X1    g0820(.A(G326), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n315), .B1(new_n572), .B2(new_n775), .C1(new_n764), .C2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G303), .A2(new_n794), .B1(new_n798), .B2(G317), .ZN(new_n1023));
  INV_X1    g0823(.A(G322), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1023), .B1(new_n969), .B2(new_n1024), .C1(new_n968), .C2(new_n840), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n858), .A2(G283), .B1(G294), .B2(new_n843), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT49), .Z(new_n1031));
  AOI21_X1  g0831(.A(new_n1022), .B1(new_n1031), .B2(KEYINPUT108), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(KEYINPUT108), .B2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n786), .A2(new_n264), .B1(new_n794), .B2(G68), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT107), .Z(new_n1035));
  NAND2_X1  g0835(.A1(new_n798), .A2(G50), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n858), .A2(new_n439), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n315), .B1(new_n843), .B2(G77), .ZN(new_n1038));
  AND4_X1   g0838(.A1(new_n958), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n851), .B2(new_n764), .C1(new_n324), .C2(new_n969), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1033), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1020), .B1(new_n1041), .B2(new_n758), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT109), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1042), .A2(KEYINPUT109), .B1(new_n688), .B2(new_n805), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1043), .A2(new_n1044), .B1(new_n754), .B2(new_n1001), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1002), .A2(KEYINPUT110), .A3(new_n695), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n750), .B2(new_n1001), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT110), .B1(new_n1002), .B2(new_n695), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(G393));
  NAND2_X1  g0849(.A1(new_n810), .A2(new_n253), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n806), .C1(new_n418), .C2(new_n210), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT111), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n757), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1052), .B2(new_n1051), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n315), .B(new_n847), .C1(G68), .C2(new_n843), .ZN(new_n1055));
  INV_X1    g0855(.A(G143), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n1056), .B2(new_n764), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT112), .Z(new_n1058));
  AOI22_X1  g0858(.A1(new_n785), .A2(G150), .B1(new_n798), .B2(G159), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT51), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n779), .A2(new_n220), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n794), .B2(new_n436), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n840), .B2(new_n202), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n1058), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1065), .A2(KEYINPUT113), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n287), .B1(new_n843), .B2(G283), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n222), .B2(new_n775), .C1(new_n764), .C2(new_n1024), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT114), .Z(new_n1069));
  AOI22_X1  g0869(.A1(new_n785), .A2(G317), .B1(new_n798), .B2(G311), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT52), .Z(new_n1071));
  NAND2_X1  g0871(.A1(new_n786), .A2(G303), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n794), .A2(G294), .B1(G116), .B2(new_n858), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1065), .A2(KEYINPUT113), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1066), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1054), .B1(new_n1076), .B2(new_n758), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n817), .B2(new_n976), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n754), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n999), .A2(new_n1002), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n695), .B1(new_n999), .B2(new_n1002), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1078), .B1(new_n1079), .B2(new_n999), .C1(new_n1080), .C2(new_n1081), .ZN(G390));
  NAND2_X1  g0882(.A1(new_n930), .A2(G330), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n918), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1083), .A2(new_n827), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n919), .A2(new_n910), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n899), .A2(new_n907), .A3(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n682), .B(new_n826), .C1(new_n709), .C2(new_n711), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n913), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n918), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n911), .B1(new_n905), .B2(new_n886), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1086), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n747), .A2(new_n931), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1088), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT115), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT115), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1088), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1094), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n754), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n264), .A2(new_n836), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n765), .A2(G294), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n315), .B1(new_n777), .B2(new_n216), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n855), .A2(new_n1061), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G107), .A2(new_n786), .B1(new_n785), .B2(G283), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G97), .A2(new_n794), .B1(new_n798), .B2(G116), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1103), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n765), .A2(G125), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n777), .A2(new_n851), .ZN(new_n1110));
  XOR2_X1   g0910(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1111));
  XNOR2_X1  g0911(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G159), .B2(new_n858), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT54), .B(G143), .Z(new_n1114));
  AOI22_X1  g0914(.A1(new_n794), .A2(new_n1114), .B1(new_n798), .B2(G132), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G128), .A2(new_n785), .B1(new_n786), .B2(G137), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1109), .A2(new_n1113), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n287), .B1(new_n775), .B2(new_n202), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1108), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n757), .B(new_n1102), .C1(new_n1120), .C2(new_n758), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n908), .B2(new_n804), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1085), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1088), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1098), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1124), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n747), .A2(new_n931), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1084), .B1(new_n1083), .B2(new_n827), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1128), .A2(new_n913), .A3(new_n1089), .A4(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n589), .A2(new_n627), .A3(new_n635), .A4(new_n637), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n656), .A2(new_n1131), .A3(new_n675), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n736), .A2(new_n728), .A3(new_n737), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT31), .B1(new_n1133), .B2(new_n675), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n728), .B1(new_n725), .B2(new_n740), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n738), .A2(KEYINPUT88), .ZN(new_n1137));
  OAI211_X1 g0937(.A(KEYINPUT31), .B(new_n675), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT89), .B1(new_n1139), .B2(G330), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n746), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n826), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1085), .B1(new_n1142), .B2(new_n1084), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n914), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1130), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n460), .A2(G330), .A3(new_n930), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n923), .A2(new_n648), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT116), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1127), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n918), .B1(new_n747), .B2(new_n826), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n914), .B1(new_n1152), .B2(new_n1085), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1147), .B1(new_n1153), .B2(new_n1130), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT116), .B1(new_n1100), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT117), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1100), .B2(new_n1154), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1127), .A2(KEYINPUT117), .A3(new_n1149), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n695), .A3(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1101), .B(new_n1122), .C1(new_n1156), .C2(new_n1160), .ZN(G378));
  OAI21_X1  g0961(.A(new_n1148), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n679), .B1(new_n933), .B2(new_n935), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n922), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n936), .A2(G330), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n912), .A3(new_n921), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n274), .A2(new_n881), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n308), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n308), .A2(new_n1167), .ZN(new_n1169));
  OR3_X1    g0969(.A1(new_n1168), .A2(new_n1169), .A3(KEYINPUT120), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1171));
  OAI21_X1  g0971(.A(KEYINPUT120), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1171), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1164), .A2(new_n1166), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1175), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n696), .B1(new_n1162), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1150), .B1(new_n1127), .B2(new_n1149), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1100), .A2(KEYINPUT116), .A3(new_n1154), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1147), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1175), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1176), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1179), .B1(new_n1184), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1181), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1186), .A2(new_n803), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n755), .B1(G50), .B2(new_n836), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n775), .A2(new_n260), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n315), .A2(new_n278), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1194), .B(new_n952), .C1(G77), .C2(new_n843), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n222), .B2(new_n772), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1193), .B(new_n1196), .C1(new_n439), .C2(new_n794), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G97), .A2(new_n786), .B1(new_n785), .B2(G116), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n839), .C2(new_n764), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT58), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G50), .B1(new_n277), .B2(new_n278), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1199), .A2(new_n1200), .B1(new_n1194), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n843), .A2(new_n1114), .ZN(new_n1203));
  INV_X1    g1003(.A(G128), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1203), .B1(new_n851), .B2(new_n779), .C1(new_n772), .C2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n785), .A2(G125), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n840), .B2(new_n860), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(G137), .C2(new_n794), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n765), .A2(G124), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n799), .C2(G159), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT59), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1211), .B(new_n1212), .C1(new_n1208), .C2(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1202), .B1(new_n1200), .B2(new_n1199), .C1(new_n1210), .C2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1192), .B1(new_n1215), .B2(new_n758), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1191), .A2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1188), .B2(new_n1079), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT121), .B1(new_n1190), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT121), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1221), .B(new_n1218), .C1(new_n1181), .C2(new_n1189), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1220), .A2(new_n1222), .ZN(G375));
  INV_X1    g1023(.A(new_n1145), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1147), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT122), .ZN(new_n1226));
  OR3_X1    g1026(.A1(new_n1145), .A2(new_n1148), .A3(KEYINPUT122), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n1005), .A3(new_n1149), .A4(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1084), .A2(new_n803), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n836), .A2(G68), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1037), .B1(new_n839), .B2(new_n772), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT123), .Z(new_n1232));
  AOI22_X1  g1032(.A1(G116), .A2(new_n786), .B1(new_n785), .B2(G294), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n315), .B1(new_n777), .B2(new_n418), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1234), .B(new_n955), .C1(new_n794), .C2(G107), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1233), .B(new_n1235), .C1(new_n790), .C2(new_n764), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n764), .A2(new_n1204), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G132), .A2(new_n785), .B1(new_n786), .B2(new_n1114), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n287), .B1(new_n777), .B2(new_n324), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1239), .B(new_n1193), .C1(G50), .C2(new_n858), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G150), .A2(new_n794), .B1(new_n798), .B2(G137), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1232), .A2(new_n1236), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n757), .B(new_n1230), .C1(new_n1243), .C2(new_n758), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1145), .A2(new_n754), .B1(new_n1229), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1228), .A2(new_n1245), .ZN(G381));
  INV_X1    g1046(.A(G375), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1101), .A2(new_n1122), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1158), .A2(new_n695), .A3(new_n1159), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT124), .Z(new_n1253));
  NOR3_X1   g1053(.A1(G387), .A2(G381), .A3(G390), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1247), .A2(new_n1251), .A3(new_n1253), .A4(new_n1254), .ZN(G407));
  OAI21_X1  g1055(.A(new_n1251), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G407), .B(G213), .C1(G343), .C2(new_n1256), .ZN(G409));
  NAND2_X1  g1057(.A1(new_n1149), .A2(KEYINPUT60), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1226), .A2(new_n1258), .A3(new_n1227), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1225), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n696), .B1(new_n1260), .B2(KEYINPUT60), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1245), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n864), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(G384), .A3(new_n1245), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n674), .A2(G213), .A3(G2897), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1266), .ZN(new_n1268));
  AOI21_X1  g1068(.A(G384), .B1(new_n1262), .B2(new_n1245), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1245), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n864), .B(new_n1270), .C1(new_n1259), .C2(new_n1261), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1268), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1188), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT57), .B1(new_n1162), .B2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1187), .A2(KEYINPUT57), .A3(new_n1176), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n695), .B1(new_n1184), .B2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G378), .B(new_n1219), .C1(new_n1276), .C2(new_n1278), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1184), .A2(new_n1188), .A3(new_n1004), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1251), .B1(new_n1280), .B2(new_n1218), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n674), .A2(G213), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT61), .B1(new_n1274), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT63), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1286), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n989), .A2(new_n1006), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n973), .A3(G390), .ZN(new_n1291));
  INV_X1    g1091(.A(G390), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(G387), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(G393), .B(new_n822), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1294), .A2(KEYINPUT125), .A3(new_n1295), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT126), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1291), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1295), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1290), .A2(KEYINPUT126), .A3(new_n973), .A4(G390), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .A4(new_n1293), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1298), .A2(new_n1299), .A3(new_n1304), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n1279), .A2(new_n1281), .B1(G213), .B2(new_n674), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1285), .A2(new_n1289), .A3(new_n1305), .A4(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1306), .A2(new_n1309), .A3(new_n1287), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT61), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1306), .B2(new_n1273), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1309), .B1(new_n1306), .B2(new_n1287), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1310), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1308), .B1(new_n1314), .B2(new_n1305), .ZN(G405));
  INV_X1    g1115(.A(KEYINPUT127), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1219), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1221), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1190), .A2(KEYINPUT121), .A3(new_n1219), .ZN(new_n1319));
  AOI21_X1  g1119(.A(G378), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1317), .A2(G378), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1320), .A2(new_n1287), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1288), .B1(new_n1256), .B2(new_n1321), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1316), .B(new_n1305), .C1(new_n1323), .C2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1305), .A2(new_n1316), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1287), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1256), .A2(new_n1288), .A3(new_n1321), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1298), .A2(KEYINPUT127), .A3(new_n1304), .A4(new_n1299), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1326), .A2(new_n1327), .A3(new_n1328), .A4(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1325), .A2(new_n1330), .ZN(G402));
endmodule


