//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT64), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT65), .B(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT67), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n218), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT68), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND4_X1  g0051(.A1(KEYINPUT70), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n252), .A2(new_n215), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT70), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n254), .B1(new_n208), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G13), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n258), .A2(new_n216), .A3(G1), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(G50), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n259), .ZN(new_n264));
  INV_X1    g0064(.A(new_n257), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT8), .B(G58), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n216), .A2(G33), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n266), .A2(new_n267), .B1(new_n216), .B2(new_n201), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n216), .A2(new_n255), .A3(KEYINPUT71), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT71), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G20), .B2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n268), .B1(G150), .B2(new_n272), .ZN(new_n273));
  OAI221_X1 g0073(.A(new_n263), .B1(G50), .B2(new_n264), .C1(new_n265), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT9), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT69), .B(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(G222), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(G223), .A3(G1698), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n278), .B(new_n279), .C1(new_n222), .C2(new_n276), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n215), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n284), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n285), .B1(G226), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n282), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n274), .A2(new_n275), .B1(G200), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n293), .B1(new_n275), .B2(new_n274), .C1(new_n294), .C2(new_n292), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(new_n292), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n274), .B1(new_n297), .B2(G169), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n292), .A2(G179), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n269), .A2(new_n271), .ZN(new_n303));
  INV_X1    g0103(.A(G50), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n267), .A2(new_n202), .B1(new_n216), .B2(G68), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n257), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT11), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n259), .A2(new_n220), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT12), .ZN(new_n311));
  OAI211_X1 g0111(.A(KEYINPUT11), .B(new_n257), .C1(new_n305), .C2(new_n306), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n260), .A2(G68), .A3(new_n262), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n309), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT75), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT14), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n277), .A2(G226), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G232), .A2(G1698), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G97), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT74), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT74), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(G33), .A3(G97), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n281), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n285), .B1(G238), .B2(new_n290), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n329), .B2(new_n331), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n316), .B(G169), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT69), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT69), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G1698), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G226), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n322), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n328), .B1(new_n341), .B2(new_n276), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n331), .B1(new_n342), .B2(new_n288), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT13), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(G179), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n334), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n345), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n316), .B1(new_n348), .B2(G169), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n315), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n332), .A2(new_n333), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n314), .B1(new_n352), .B2(G190), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(G200), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n276), .B1(new_n221), .B2(new_n335), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n339), .A2(new_n235), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n281), .B1(G107), .B2(new_n276), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n285), .B1(G244), .B2(new_n290), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n294), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(G200), .B2(new_n360), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n260), .A2(G77), .A3(new_n262), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n222), .A2(new_n259), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT72), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n216), .A2(new_n222), .B1(new_n366), .B2(new_n267), .ZN(new_n367));
  INV_X1    g0167(.A(new_n266), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n367), .B1(new_n272), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n363), .B(new_n365), .C1(new_n265), .C2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT73), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n371), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n362), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G169), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n360), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n376), .B(new_n370), .C1(G179), .C2(new_n360), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NOR4_X1   g0178(.A1(new_n302), .A2(new_n351), .A3(new_n355), .A4(new_n378), .ZN(new_n379));
  XNOR2_X1  g0179(.A(G58), .B(G68), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n272), .A2(G159), .B1(new_n380), .B2(G20), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n276), .B2(G20), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT78), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n320), .A2(new_n216), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT78), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n386), .A3(new_n382), .ZN(new_n387));
  OR3_X1    g0187(.A1(new_n255), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n319), .A2(KEYINPUT79), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n388), .B(new_n389), .C1(new_n390), .C2(G33), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n382), .A2(G20), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n384), .A2(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n381), .B1(new_n393), .B2(new_n220), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n318), .A2(KEYINPUT76), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT76), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT3), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n399), .A3(G33), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n317), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(new_n382), .A3(new_n216), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G68), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n382), .B1(new_n401), .B2(new_n216), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT16), .B(new_n381), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT77), .ZN(new_n406));
  INV_X1    g0206(.A(new_n317), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n390), .B2(G33), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT7), .B1(new_n408), .B2(G20), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(G68), .A3(new_n402), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT77), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT16), .A4(new_n381), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n396), .A2(new_n406), .A3(new_n257), .A4(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n266), .B1(new_n261), .B2(G20), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n260), .A2(new_n414), .B1(new_n259), .B2(new_n266), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n288), .A2(G274), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n235), .A2(new_n289), .B1(new_n417), .B2(new_n284), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n277), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n419));
  INV_X1    g0219(.A(G87), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n419), .A2(new_n401), .B1(new_n255), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n418), .B1(new_n421), .B2(new_n281), .ZN(new_n422));
  INV_X1    g0222(.A(G179), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT80), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n422), .A2(G169), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT80), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n422), .A2(new_n427), .A3(new_n423), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n416), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT18), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n416), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n422), .A2(G190), .ZN(new_n436));
  INV_X1    g0236(.A(G200), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n437), .B2(new_n422), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n413), .A2(new_n415), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n413), .A2(new_n439), .A3(KEYINPUT17), .A4(new_n415), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n435), .A2(KEYINPUT81), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n432), .A2(new_n434), .A3(new_n442), .A4(new_n443), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n379), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n420), .A2(KEYINPUT22), .A3(G20), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n276), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT87), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT87), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n276), .A2(new_n454), .A3(new_n451), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n408), .A2(new_n216), .A3(G87), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(KEYINPUT22), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G116), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G20), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT23), .B1(new_n205), .B2(G20), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT24), .B1(new_n458), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n457), .A2(KEYINPUT22), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(new_n464), .C1(new_n468), .C2(new_n456), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n265), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n281), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G264), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(new_n472), .A3(new_n473), .ZN(new_n477));
  INV_X1    g0277(.A(G250), .ZN(new_n478));
  INV_X1    g0278(.A(G257), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n339), .A2(new_n478), .B1(new_n479), .B2(new_n335), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n480), .A2(new_n408), .B1(G33), .B2(G294), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n475), .B(new_n477), .C1(new_n481), .C2(new_n288), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G200), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n294), .B2(new_n482), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n259), .A2(new_n205), .ZN(new_n485));
  XOR2_X1   g0285(.A(new_n485), .B(KEYINPUT25), .Z(new_n486));
  NAND2_X1  g0286(.A1(new_n261), .A2(G33), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n260), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(new_n205), .ZN(new_n489));
  OR3_X1    g0289(.A1(new_n470), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT88), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n277), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n492));
  INV_X1    g0292(.A(G294), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n492), .A2(new_n401), .B1(new_n255), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(new_n281), .B1(G264), .B2(new_n474), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n375), .B1(new_n495), .B2(new_n477), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n482), .A2(new_n423), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n491), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n482), .A2(G169), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n499), .B(KEYINPUT88), .C1(new_n423), .C2(new_n482), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n498), .B(new_n500), .C1(new_n470), .C2(new_n489), .ZN(new_n501));
  AND2_X1   g0301(.A1(KEYINPUT5), .A2(G41), .ZN(new_n502));
  NOR2_X1   g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n472), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(G257), .A3(new_n288), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n477), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT83), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT83), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n477), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(KEYINPUT4), .A2(G244), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n276), .A2(new_n277), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G283), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  XOR2_X1   g0315(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n516));
  NAND2_X1  g0316(.A1(new_n277), .A2(G244), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n401), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n288), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n375), .B1(new_n510), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n509), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n508), .B1(new_n477), .B2(new_n505), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n516), .ZN(new_n524));
  INV_X1    g0324(.A(new_n517), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(new_n408), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n281), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n523), .A2(new_n423), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n520), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n264), .A2(G97), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n488), .B2(new_n204), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT6), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n534), .A2(new_n204), .A3(G107), .ZN(new_n535));
  XNOR2_X1  g0335(.A(G97), .B(G107), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n537), .A2(new_n216), .B1(new_n202), .B2(new_n303), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n393), .B2(new_n205), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n533), .B1(new_n540), .B2(new_n257), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n530), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n510), .A2(new_n519), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G190), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(new_n541), .C1(new_n437), .C2(new_n544), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n490), .A2(new_n501), .A3(new_n543), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n476), .A2(new_n472), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT84), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n261), .A3(G45), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT84), .B1(new_n471), .B2(G1), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n288), .A2(G250), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n336), .A2(new_n338), .A3(G238), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G244), .A2(G1698), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n408), .A2(new_n556), .B1(G33), .B2(G116), .ZN(new_n557));
  OAI211_X1 g0357(.A(G179), .B(new_n553), .C1(new_n557), .C2(new_n288), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT85), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n548), .A2(new_n552), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n277), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n459), .B1(new_n561), .B2(new_n401), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n560), .B1(new_n562), .B2(new_n281), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n558), .B(new_n559), .C1(new_n563), .C2(new_n375), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n553), .B1(new_n557), .B2(new_n288), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G169), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n559), .B1(new_n567), .B2(new_n558), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n400), .A2(new_n216), .A3(G68), .A4(new_n317), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n267), .B2(new_n204), .ZN(new_n572));
  AOI21_X1  g0372(.A(G20), .B1(new_n328), .B2(KEYINPUT19), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n206), .A2(G87), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n570), .B(new_n572), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n257), .ZN(new_n576));
  INV_X1    g0376(.A(new_n366), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n264), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT86), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT86), .ZN(new_n581));
  AOI211_X1 g0381(.A(new_n581), .B(new_n578), .C1(new_n575), .C2(new_n257), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n580), .A2(new_n582), .B1(new_n488), .B2(new_n366), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n570), .A2(new_n572), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n571), .B1(new_n325), .B2(new_n327), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n585), .A2(G20), .B1(G87), .B2(new_n206), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n265), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n581), .B1(new_n587), .B2(new_n578), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n576), .A2(KEYINPUT86), .A3(new_n579), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n265), .A2(new_n264), .A3(new_n487), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n588), .A2(new_n589), .B1(G87), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n563), .A2(G190), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n408), .A2(new_n556), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n288), .B1(new_n593), .B2(new_n459), .ZN(new_n594));
  OAI21_X1  g0394(.A(G200), .B1(new_n594), .B2(new_n560), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n569), .A2(new_n583), .B1(new_n591), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT21), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n265), .A2(G116), .A3(new_n264), .A4(new_n487), .ZN(new_n600));
  INV_X1    g0400(.A(G116), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n259), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(G20), .B1(G33), .B2(G283), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n255), .A2(G97), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n603), .A2(new_n604), .B1(G20), .B2(new_n601), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n257), .A2(KEYINPUT20), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT20), .B1(new_n257), .B2(new_n605), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n600), .B(new_n602), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n504), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n474), .A2(G270), .B1(new_n610), .B2(new_n476), .ZN(new_n611));
  NAND2_X1  g0411(.A1(G264), .A2(G1698), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n339), .B2(new_n479), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n613), .A2(new_n408), .B1(G303), .B2(new_n320), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n611), .B1(new_n614), .B2(new_n288), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G169), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n599), .B1(new_n609), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(G200), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n611), .B(G190), .C1(new_n614), .C2(new_n288), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n609), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n615), .A2(new_n423), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n608), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n608), .A2(new_n615), .A3(KEYINPUT21), .A4(G169), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n617), .A2(new_n620), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n598), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n450), .A2(new_n547), .A3(new_n625), .ZN(G372));
  OAI21_X1  g0426(.A(new_n350), .B1(new_n355), .B2(new_n377), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n444), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n435), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n300), .B1(new_n629), .B2(new_n296), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n617), .A2(new_n622), .A3(new_n623), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n470), .A2(new_n489), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n499), .B1(new_n423), .B2(new_n482), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n490), .A2(new_n543), .A3(new_n546), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT89), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n595), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n566), .A2(KEYINPUT89), .A3(G200), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n638), .A2(new_n592), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n567), .A2(new_n558), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n640), .A2(new_n591), .B1(new_n583), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n635), .A2(new_n636), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT91), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n583), .A2(new_n641), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT90), .B1(new_n530), .B2(new_n541), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n588), .A2(new_n589), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n590), .A2(G87), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n595), .A2(new_n637), .B1(G190), .B2(new_n563), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .A4(new_n639), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n531), .B1(new_n590), .B2(G97), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n391), .A2(new_n392), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n386), .B1(new_n385), .B2(new_n382), .ZN(new_n654));
  AOI211_X1 g0454(.A(KEYINPUT78), .B(KEYINPUT7), .C1(new_n320), .C2(new_n216), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n538), .B1(new_n656), .B2(G107), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n652), .B1(new_n657), .B2(new_n265), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT90), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(new_n529), .A4(new_n520), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n647), .A2(new_n651), .A3(new_n646), .A4(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n646), .B1(new_n661), .B2(KEYINPUT26), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n598), .B2(new_n542), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n645), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n569), .A2(new_n583), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n591), .A2(new_n597), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n542), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT26), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n642), .A2(new_n663), .A3(new_n647), .A4(new_n660), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(KEYINPUT91), .A4(new_n646), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n644), .B1(new_n665), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n630), .B1(new_n450), .B2(new_n672), .ZN(G369));
  AND2_X1   g0473(.A1(new_n490), .A2(new_n501), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n261), .A2(new_n216), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n632), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT92), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n682), .A2(KEYINPUT92), .ZN(new_n685));
  OAI22_X1  g0485(.A1(new_n684), .A2(new_n685), .B1(new_n501), .B2(new_n681), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n608), .A2(new_n680), .ZN(new_n687));
  MUX2_X1   g0487(.A(new_n631), .B(new_n624), .S(new_n687), .Z(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n684), .A2(new_n685), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n631), .A2(new_n681), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n680), .B(KEYINPUT93), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n633), .A2(new_n634), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT94), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT94), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n695), .A2(new_n700), .A3(new_n697), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n692), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT95), .ZN(G399));
  INV_X1    g0503(.A(new_n210), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n574), .A2(new_n601), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n213), .B2(new_n706), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT96), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n523), .A2(new_n495), .A3(new_n528), .A4(new_n563), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n615), .A2(new_n423), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n495), .A2(new_n563), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n544), .A3(KEYINPUT30), .A4(new_n621), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n482), .B1(new_n510), .B2(new_n519), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n615), .A2(new_n566), .A3(new_n423), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT97), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT97), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n615), .A2(new_n566), .A3(new_n724), .A4(new_n423), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n721), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n713), .B1(new_n727), .B2(new_n681), .ZN(new_n728));
  INV_X1    g0528(.A(new_n696), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT31), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n728), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n547), .A2(new_n625), .A3(new_n729), .ZN(new_n732));
  OAI21_X1  g0532(.A(G330), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT98), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT98), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n735), .B(G330), .C1(new_n731), .C2(new_n732), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n672), .A2(new_n729), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT29), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n661), .A2(KEYINPUT26), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n598), .A2(new_n663), .A3(new_n542), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(new_n646), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(KEYINPUT99), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n636), .A2(new_n643), .ZN(new_n744));
  INV_X1    g0544(.A(new_n501), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n745), .B2(new_n631), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n742), .A2(KEYINPUT99), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n680), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT29), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n737), .B1(new_n739), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n712), .B1(new_n751), .B2(G1), .ZN(G364));
  NOR2_X1   g0552(.A1(new_n258), .A2(G20), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G45), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(G1), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n705), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n690), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G330), .B2(new_n688), .ZN(new_n760));
  OAI21_X1  g0560(.A(G20), .B1(KEYINPUT103), .B2(G169), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(KEYINPUT103), .A2(G169), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n215), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n294), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n216), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n204), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n216), .A2(G179), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(new_n294), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G107), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n216), .A2(new_n423), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n437), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n772), .B1(new_n776), .B2(new_n304), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n774), .A2(G200), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n768), .B(new_n777), .C1(G58), .C2(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT104), .B(KEYINPUT32), .Z(new_n780));
  NOR2_X1   g0580(.A1(G190), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n769), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n769), .A2(G190), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n785), .B1(G87), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n773), .A2(new_n294), .A3(G200), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n276), .B1(new_n789), .B2(new_n220), .ZN(new_n790));
  INV_X1    g0590(.A(new_n222), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n773), .A2(new_n781), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n790), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n779), .A2(new_n784), .A3(new_n788), .A4(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n793), .A2(G311), .ZN(new_n796));
  INV_X1    g0596(.A(new_n789), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n276), .B(new_n796), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  INV_X1    g0600(.A(G329), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n770), .A2(new_n800), .B1(new_n782), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT105), .Z(new_n803));
  AOI22_X1  g0603(.A1(G322), .A2(new_n778), .B1(new_n775), .B2(G326), .ZN(new_n804));
  INV_X1    g0604(.A(new_n767), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n805), .A2(G294), .B1(new_n787), .B2(G303), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n799), .A2(new_n803), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n765), .B1(new_n795), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT102), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n764), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n210), .A2(new_n401), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT101), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n250), .A2(G45), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(G45), .C2(new_n213), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n704), .A2(new_n320), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n818), .A2(G355), .B1(new_n601), .B2(new_n704), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n813), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n758), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n808), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n811), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n688), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n760), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  NAND2_X1  g0626(.A1(new_n370), .A2(new_n680), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n374), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n377), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n377), .A2(new_n680), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n696), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n738), .A2(new_n832), .B1(new_n672), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n737), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n758), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  INV_X1    g0637(.A(new_n809), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n765), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G294), .A2(new_n778), .B1(new_n775), .B2(G303), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n205), .B2(new_n786), .ZN(new_n841));
  INV_X1    g0641(.A(new_n782), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G116), .A2(new_n793), .B1(new_n842), .B2(G311), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(new_n320), .C1(new_n800), .C2(new_n789), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n770), .A2(new_n420), .ZN(new_n845));
  NOR4_X1   g0645(.A1(new_n841), .A2(new_n844), .A3(new_n768), .A4(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n797), .A2(G150), .B1(new_n793), .B2(G159), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  INV_X1    g0648(.A(G143), .ZN(new_n849));
  INV_X1    g0649(.A(new_n778), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n847), .B1(new_n776), .B2(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n408), .B1(new_n854), .B2(new_n782), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n770), .A2(new_n220), .ZN(new_n856));
  INV_X1    g0656(.A(G58), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n767), .A2(new_n857), .B1(new_n786), .B2(new_n304), .ZN(new_n858));
  NOR4_X1   g0658(.A1(new_n853), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n851), .A2(new_n852), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n846), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n758), .B1(G77), .B2(new_n839), .C1(new_n861), .C2(new_n765), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT106), .Z(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n810), .B2(new_n832), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n837), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(G384));
  NOR2_X1   g0666(.A1(new_n753), .A2(new_n261), .ZN(new_n867));
  INV_X1    g0667(.A(new_n678), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n435), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n406), .A2(new_n257), .A3(new_n412), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT16), .B1(new_n410), .B2(new_n381), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n415), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n446), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n429), .A2(new_n678), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n440), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT37), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(KEYINPUT109), .B(KEYINPUT37), .Z(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n416), .A2(new_n874), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n440), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n877), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n873), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT39), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n446), .A2(new_n416), .A3(new_n868), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT110), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n881), .A2(new_n891), .A3(new_n879), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n880), .B(new_n440), .C1(new_n890), .C2(new_n878), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(KEYINPUT111), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT111), .B1(new_n892), .B2(new_n893), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n884), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(KEYINPUT112), .B(KEYINPUT39), .Z(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(new_n886), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT108), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n350), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n315), .B(KEYINPUT108), .C1(new_n347), .C2(new_n349), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(new_n680), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n869), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n315), .A2(new_n680), .B1(new_n353), .B2(new_n354), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n902), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n347), .A2(new_n349), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n315), .B(new_n680), .C1(new_n909), .C2(new_n355), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n830), .B1(new_n672), .B2(new_n833), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT107), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT107), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n915), .B(new_n830), .C1(new_n672), .C2(new_n833), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n912), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n887), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n906), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n739), .A2(new_n750), .A3(new_n449), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n630), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(KEYINPUT31), .B(new_n680), .C1(new_n720), .C2(new_n726), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n728), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n732), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n911), .A2(new_n832), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT113), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n624), .A2(new_n666), .A3(new_n667), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n543), .A2(new_n546), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n928), .A2(new_n674), .A3(new_n929), .A4(new_n696), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(new_n728), .A3(new_n923), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT113), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n831), .B1(new_n908), .B2(new_n910), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n873), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n873), .B2(new_n882), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n927), .B(new_n934), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n897), .A2(new_n886), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n931), .A2(KEYINPUT40), .A3(new_n933), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n937), .A2(new_n938), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n450), .B2(new_n925), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n449), .A3(new_n931), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n944), .A2(G330), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n867), .B1(new_n922), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n922), .B2(new_n946), .ZN(new_n948));
  INV_X1    g0748(.A(new_n537), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n949), .A2(KEYINPUT35), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(KEYINPUT35), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n950), .A2(G116), .A3(new_n217), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT36), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n214), .B1(new_n857), .B2(new_n220), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n954), .A2(new_n222), .B1(G50), .B2(new_n220), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(G1), .A3(new_n258), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n948), .A2(new_n953), .A3(new_n956), .ZN(G367));
  OAI21_X1  g0757(.A(new_n929), .B1(new_n541), .B2(new_n696), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n530), .A2(new_n541), .A3(new_n696), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT114), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n960), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n543), .B1(new_n964), .B2(new_n501), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n729), .B1(new_n965), .B2(KEYINPUT115), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(KEYINPUT115), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n695), .A2(new_n964), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT42), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n591), .A2(new_n681), .ZN(new_n970));
  MUX2_X1   g0770(.A(new_n643), .B(new_n646), .S(new_n970), .Z(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n967), .A2(new_n969), .B1(KEYINPUT43), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(KEYINPUT43), .B2(new_n972), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT43), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n967), .A2(new_n969), .A3(new_n975), .A4(new_n971), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n691), .A2(new_n964), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n705), .B(KEYINPUT41), .Z(new_n980));
  AOI21_X1  g0780(.A(new_n964), .B1(new_n699), .B2(new_n701), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT45), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n699), .A2(new_n701), .A3(new_n964), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT44), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n692), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n695), .B1(new_n686), .B2(new_n694), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(new_n689), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n982), .A2(new_n985), .A3(new_n691), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n987), .A2(new_n751), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n980), .B1(new_n992), .B2(new_n751), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n979), .B1(new_n993), .B2(new_n757), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n815), .A2(new_n241), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n813), .B1(new_n704), .B2(new_n577), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n821), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n776), .A2(new_n849), .B1(new_n786), .B2(new_n857), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G150), .B2(new_n778), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n792), .A2(new_n304), .B1(new_n782), .B2(new_n848), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n320), .B(new_n1000), .C1(G159), .C2(new_n797), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n805), .A2(G68), .B1(new_n771), .B2(new_n791), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G107), .A2(new_n805), .B1(new_n775), .B2(G311), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n204), .B2(new_n770), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n789), .A2(new_n493), .B1(new_n792), .B2(new_n800), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G317), .B2(new_n842), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n408), .B1(new_n778), .B2(G303), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT46), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n786), .B2(new_n601), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n787), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1003), .B1(new_n1005), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT47), .Z(new_n1014));
  OAI221_X1 g0814(.A(new_n997), .B1(new_n765), .B2(new_n1014), .C1(new_n972), .C2(new_n823), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n994), .A2(new_n1015), .ZN(G387));
  NAND2_X1  g0816(.A1(new_n751), .A2(new_n990), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n705), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n751), .A2(new_n990), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n686), .A2(new_n823), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n815), .B1(new_n238), .B2(new_n471), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n818), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1022), .B1(new_n708), .B2(new_n1023), .ZN(new_n1024));
  OR3_X1    g0824(.A1(new_n266), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1025));
  OAI21_X1  g0825(.A(KEYINPUT50), .B1(new_n266), .B2(G50), .ZN(new_n1026));
  AOI21_X1  g0826(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1025), .A2(new_n708), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1024), .A2(new_n1028), .B1(new_n205), .B2(new_n704), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n758), .B1(new_n1029), .B2(new_n813), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n776), .A2(new_n783), .B1(new_n222), .B2(new_n786), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n797), .A2(new_n368), .B1(new_n842), .B2(G150), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n220), .B2(new_n792), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n850), .A2(new_n304), .B1(new_n366), .B2(new_n767), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n408), .B1(new_n204), .B2(new_n770), .ZN(new_n1035));
  OR4_X1    g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n797), .A2(G311), .B1(new_n793), .B2(G303), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n778), .A2(G317), .ZN(new_n1038));
  INV_X1    g0838(.A(G322), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1037), .B(new_n1038), .C1(new_n1039), .C2(new_n776), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n800), .B2(new_n767), .C1(new_n493), .C2(new_n786), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(KEYINPUT49), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n770), .A2(new_n601), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n408), .B(new_n1047), .C1(G326), .C2(new_n842), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1045), .A2(KEYINPUT49), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1036), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1030), .B1(new_n1051), .B2(new_n764), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n990), .A2(new_n757), .B1(new_n1021), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1020), .A2(new_n1053), .ZN(G393));
  INV_X1    g0854(.A(new_n991), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n691), .B1(new_n982), .B2(new_n985), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1017), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(new_n992), .A3(new_n705), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n815), .A2(new_n247), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n812), .B1(new_n204), .B2(new_n210), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G311), .A2(new_n778), .B1(new_n775), .B2(G317), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT52), .Z(new_n1062));
  OAI221_X1 g0862(.A(new_n772), .B1(new_n800), .B2(new_n786), .C1(new_n601), .C2(new_n767), .ZN(new_n1063));
  INV_X1    g0863(.A(G303), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n320), .B1(new_n789), .B2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n792), .A2(new_n493), .B1(new_n782), .B2(new_n1039), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G150), .A2(new_n775), .B1(new_n778), .B2(G159), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT51), .Z(new_n1069));
  AOI22_X1  g0869(.A1(new_n797), .A2(G50), .B1(new_n842), .B2(G143), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n266), .B2(new_n792), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n767), .A2(new_n202), .B1(new_n786), .B2(new_n220), .ZN(new_n1072));
  NOR4_X1   g0872(.A1(new_n1071), .A2(new_n401), .A3(new_n845), .A4(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1062), .A2(new_n1067), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n758), .B1(new_n1059), .B2(new_n1060), .C1(new_n1074), .C2(new_n765), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n964), .B2(new_n811), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1076), .B1(new_n1077), .B2(new_n757), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1058), .A2(new_n1078), .ZN(G390));
  INV_X1    g0879(.A(new_n896), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1080), .A2(new_n889), .A3(new_n894), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n935), .B1(new_n1081), .B2(new_n884), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1082), .A2(new_n898), .B1(KEYINPUT39), .B2(new_n887), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n917), .B2(new_n905), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n905), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n830), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n749), .B2(new_n829), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n911), .B(KEYINPUT116), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1085), .B(new_n939), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n831), .B1(new_n734), .B2(new_n736), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n911), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1084), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n931), .A2(G330), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n933), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n449), .A2(new_n1094), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n920), .A2(new_n630), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1094), .A2(new_n832), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1090), .A2(new_n911), .B1(new_n1101), .B2(new_n1088), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n1087), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1095), .B1(new_n1090), .B2(new_n911), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n914), .A2(new_n916), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT117), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1097), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1108), .B(new_n1109), .C1(new_n1092), .C2(new_n1096), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n705), .A3(new_n1112), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n900), .A2(new_n810), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n758), .B1(new_n368), .B2(new_n839), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n601), .A2(new_n850), .B1(new_n776), .B2(new_n800), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n856), .B(new_n1116), .C1(G77), .C2(new_n805), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n320), .B1(new_n782), .B2(new_n493), .C1(new_n420), .C2(new_n786), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n789), .A2(new_n205), .B1(new_n792), .B2(new_n204), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(KEYINPUT119), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1117), .B(new_n1120), .C1(KEYINPUT119), .C2(new_n1119), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n789), .A2(new_n848), .B1(new_n792), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G159), .B2(new_n805), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT118), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n787), .A2(G150), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n320), .B1(new_n842), .B2(G125), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n850), .B2(new_n854), .ZN(new_n1129));
  INV_X1    g0929(.A(G128), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n776), .A2(new_n1130), .B1(new_n770), .B2(new_n304), .ZN(new_n1131));
  OR3_X1    g0931(.A1(new_n1127), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1121), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1115), .B1(new_n1133), .B2(new_n764), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1097), .A2(new_n757), .B1(new_n1114), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1113), .A2(new_n1135), .ZN(G378));
  NAND2_X1  g0936(.A1(new_n937), .A2(new_n938), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n939), .A2(new_n941), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n274), .A2(new_n868), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n296), .A2(new_n301), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1139), .B1(new_n296), .B2(new_n301), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OR3_X1    g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AND4_X1   g0947(.A1(G330), .A2(new_n1137), .A3(new_n1138), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(new_n942), .B2(G330), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n919), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1137), .A2(G330), .A3(new_n1138), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1147), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n942), .A2(G330), .A3(new_n1147), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1153), .A2(new_n1154), .A3(new_n918), .A4(new_n906), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1147), .A2(new_n810), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n758), .B1(G50), .B2(new_n839), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n771), .A2(G58), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n776), .B2(new_n601), .C1(new_n205), .C2(new_n850), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n408), .A2(G41), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n797), .A2(G97), .B1(new_n842), .B2(G283), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n366), .B2(new_n792), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n767), .A2(new_n220), .B1(new_n786), .B2(new_n222), .ZN(new_n1164));
  OR4_X1    g0964(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT58), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1161), .B(new_n304), .C1(G33), .C2(G41), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G150), .A2(new_n805), .B1(new_n775), .B2(G125), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1130), .B2(new_n850), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n786), .A2(new_n1122), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n789), .A2(new_n854), .B1(new_n792), .B2(new_n848), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n771), .A2(G159), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G33), .B(G41), .C1(new_n842), .C2(G124), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1169), .B1(new_n1166), .B2(new_n1165), .C1(new_n1176), .C2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1158), .B1(new_n1181), .B2(new_n764), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1156), .A2(new_n757), .B1(new_n1157), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1102), .A2(new_n1087), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1092), .A2(new_n1096), .A3(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1187), .B2(new_n1099), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n705), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1084), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n939), .A2(new_n1085), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n748), .A2(new_n743), .A3(new_n746), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n681), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n829), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n830), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1088), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1191), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1105), .A2(new_n911), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1085), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1197), .B1(new_n1199), .B2(new_n1083), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1190), .B(new_n1107), .C1(new_n1200), .C2(new_n1095), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1100), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1156), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1183), .B1(new_n1189), .B2(new_n1203), .ZN(G375));
  NAND2_X1  g1004(.A1(new_n1186), .A2(new_n1099), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n980), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1108), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1088), .A2(new_n809), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n758), .B1(G68), .B2(new_n839), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n202), .A2(new_n770), .B1(new_n786), .B2(new_n204), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n577), .A2(new_n805), .B1(new_n775), .B2(G294), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n276), .B1(new_n793), .B2(G107), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n797), .A2(G116), .B1(new_n842), .B2(G303), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1210), .B(new_n1214), .C1(G283), .C2(new_n778), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1216), .A2(KEYINPUT121), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n767), .A2(new_n304), .B1(new_n786), .B2(new_n783), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n793), .A2(G150), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n1130), .B2(new_n782), .C1(new_n789), .C2(new_n1122), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n854), .A2(new_n776), .B1(new_n850), .B2(new_n848), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1159), .A2(new_n408), .ZN(new_n1222));
  OR4_X1    g1022(.A1(new_n1218), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1216), .A2(KEYINPUT121), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1217), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1209), .B1(new_n1225), .B2(new_n764), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1107), .A2(new_n757), .B1(new_n1208), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1207), .A2(new_n1227), .ZN(G381));
  NAND3_X1  g1028(.A1(new_n1020), .A2(new_n825), .A3(new_n1053), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1058), .A2(new_n1078), .A3(new_n865), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(G387), .A2(G381), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(G378), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1201), .A2(new_n1100), .B1(new_n1155), .B2(new_n1150), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1188), .B(new_n705), .C1(new_n1233), .C2(KEYINPUT57), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1231), .A2(new_n1232), .A3(new_n1234), .A4(new_n1183), .ZN(G407));
  NAND2_X1  g1035(.A1(new_n679), .A2(G213), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT122), .ZN(new_n1237));
  OR3_X1    g1037(.A1(G375), .A2(G378), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G407), .A2(G213), .A3(new_n1238), .ZN(G409));
  NAND3_X1  g1039(.A1(new_n1234), .A2(G378), .A3(new_n1183), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1233), .A2(new_n1206), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1241), .A2(new_n1183), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(G378), .B2(new_n1242), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1243), .A2(new_n1237), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT123), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT60), .B1(new_n1205), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT60), .ZN(new_n1247));
  AOI211_X1 g1047(.A(KEYINPUT123), .B(new_n1247), .C1(new_n1186), .C2(new_n1099), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n705), .B(new_n1108), .C1(new_n1246), .C2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(G384), .A3(new_n1227), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G384), .B1(new_n1249), .B2(new_n1227), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1244), .A2(KEYINPUT63), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(G2897), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1236), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1253), .A2(KEYINPUT124), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT124), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1249), .A2(new_n1227), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n865), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1250), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1259), .B1(new_n1262), .B2(new_n1256), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1258), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1243), .A2(new_n1236), .ZN(new_n1265));
  OR3_X1    g1065(.A1(new_n1253), .A2(new_n1255), .A3(new_n1237), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1243), .A2(new_n1236), .A3(new_n1253), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT63), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G387), .A2(KEYINPUT125), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT125), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n994), .A2(new_n1272), .A3(new_n1015), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G390), .A2(new_n1229), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1229), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1058), .A3(new_n1078), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1271), .A2(new_n1273), .A3(new_n1275), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n994), .A2(new_n1272), .A3(new_n1015), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1272), .B1(new_n994), .B2(new_n1015), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1254), .A2(new_n1267), .A3(new_n1270), .A4(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1285), .B1(new_n1286), .B2(new_n1244), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1262), .A2(new_n1288), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1244), .A2(new_n1289), .B1(new_n1268), .B2(new_n1288), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1284), .B1(new_n1291), .B2(new_n1292), .ZN(G405));
  AND3_X1   g1093(.A1(new_n1234), .A2(G378), .A3(new_n1183), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G378), .B1(new_n1234), .B2(new_n1183), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1253), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G375), .A2(new_n1232), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(new_n1262), .A3(new_n1240), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1296), .A2(new_n1297), .A3(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1300), .A2(new_n1292), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1294), .A2(new_n1295), .A3(new_n1253), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1262), .B1(new_n1298), .B2(new_n1240), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT126), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT127), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT127), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(KEYINPUT126), .A3(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1301), .A2(new_n1305), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1300), .A2(new_n1292), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1307), .B1(new_n1306), .B2(KEYINPUT126), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n1297), .B(KEYINPUT127), .C1(new_n1296), .C2(new_n1299), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1310), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1309), .A2(new_n1313), .ZN(G402));
endmodule


