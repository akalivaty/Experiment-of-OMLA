//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(G13), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n204), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G87), .A2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n220));
  AND4_X1   g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT64), .B(G238), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G68), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n205), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n210), .B(new_n215), .C1(new_n216), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n216), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n225), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G87), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(G97), .B(G107), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(new_n213), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT72), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT68), .ZN(new_n247));
  NOR3_X1   g0047(.A1(new_n247), .A2(G20), .A3(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  AOI21_X1  g0049(.A(KEYINPUT68), .B1(new_n204), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G50), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n246), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n204), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G68), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n255), .A2(G77), .B1(G20), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n251), .A2(new_n246), .A3(new_n252), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n245), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT73), .B(KEYINPUT11), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n261), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n245), .B(new_n263), .C1(new_n258), .C2(new_n259), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n244), .A2(new_n213), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n203), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G68), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(KEYINPUT12), .A3(new_n256), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT12), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(new_n268), .B2(G68), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n267), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n262), .A2(new_n264), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(G226), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G97), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G232), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n277), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  OAI211_X1 g0082(.A(G1), .B(G13), .C1(new_n249), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT66), .B(G41), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n203), .B(G274), .C1(new_n286), .C2(G45), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT67), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n290), .B(new_n203), .C1(G41), .C2(G45), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n283), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G238), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n285), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT13), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT13), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n285), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(G179), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n297), .B2(new_n299), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT14), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n299), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n298), .B1(new_n285), .B2(new_n295), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n307), .A2(KEYINPUT14), .A3(new_n301), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n274), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(G190), .ZN(new_n310));
  INV_X1    g0110(.A(new_n274), .ZN(new_n311));
  INV_X1    g0111(.A(G200), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n310), .B(new_n311), .C1(new_n312), .C2(new_n307), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n275), .A2(G222), .A3(new_n276), .ZN(new_n315));
  INV_X1    g0115(.A(G77), .ZN(new_n316));
  INV_X1    g0116(.A(G223), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n315), .B1(new_n316), .B2(new_n275), .C1(new_n279), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n284), .ZN(new_n319));
  INV_X1    g0119(.A(new_n287), .ZN(new_n320));
  INV_X1    g0120(.A(new_n292), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(G226), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OR3_X1    g0126(.A1(new_n269), .A2(new_n245), .A3(KEYINPUT70), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT70), .B1(new_n269), .B2(new_n245), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(new_n266), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(new_n252), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n269), .A2(new_n252), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G58), .A2(G68), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n204), .B1(new_n332), .B2(new_n252), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT69), .ZN(new_n334));
  INV_X1    g0134(.A(G150), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT8), .B(G58), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n251), .A2(new_n335), .B1(new_n336), .B2(new_n254), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n245), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n330), .A2(new_n331), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n323), .A2(new_n301), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n326), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT9), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n324), .A2(G190), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n330), .A2(KEYINPUT9), .A3(new_n331), .A4(new_n338), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n323), .A2(G200), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n343), .A2(new_n344), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n347), .A2(KEYINPUT10), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(KEYINPUT10), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n341), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT3), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G33), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n351), .A2(new_n353), .A3(G232), .A4(new_n276), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT71), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n275), .A2(KEYINPUT71), .A3(G232), .A4(new_n276), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n222), .A2(new_n275), .A3(G1698), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n351), .A2(new_n353), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G107), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n356), .A2(new_n357), .A3(new_n358), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n284), .ZN(new_n362));
  INV_X1    g0162(.A(G244), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n287), .B1(new_n292), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n301), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n362), .A2(new_n325), .A3(new_n365), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n251), .A2(new_n336), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT15), .B(G87), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n370), .A2(new_n254), .B1(new_n204), .B2(new_n316), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n245), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n265), .A2(G77), .A3(new_n266), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n269), .A2(new_n316), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n367), .A2(new_n368), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n362), .A2(G190), .A3(new_n365), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n373), .A2(new_n374), .ZN(new_n378));
  XOR2_X1   g0178(.A(KEYINPUT15), .B(G87), .Z(new_n379));
  AOI22_X1  g0179(.A1(new_n379), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n251), .B2(new_n336), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n378), .B1(new_n381), .B2(new_n245), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n364), .B1(new_n284), .B2(new_n361), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n377), .B(new_n382), .C1(new_n312), .C2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n314), .A2(new_n350), .A3(new_n376), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n275), .B2(G20), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n359), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n256), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(G58), .A2(G68), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n390), .B2(new_n332), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT74), .ZN(new_n392));
  OAI21_X1  g0192(.A(G159), .B1(new_n248), .B2(new_n250), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT74), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(G20), .C1(new_n390), .C2(new_n332), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT75), .B1(new_n389), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT16), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT75), .B(new_n399), .C1(new_n389), .C2(new_n396), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n400), .A3(new_n245), .ZN(new_n401));
  INV_X1    g0201(.A(new_n336), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n268), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n329), .B2(new_n336), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n287), .B1(new_n292), .B2(new_n280), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n351), .A2(new_n353), .A3(G226), .A4(G1698), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n351), .A2(new_n353), .A3(G223), .A4(new_n276), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G87), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT76), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n283), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT76), .A4(new_n410), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n407), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G190), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(new_n412), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n414), .A3(new_n284), .ZN(new_n418));
  INV_X1    g0218(.A(new_n407), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G200), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n401), .A2(new_n406), .A3(new_n416), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT17), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n265), .B1(new_n397), .B2(KEYINPUT16), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n405), .B1(new_n424), .B2(new_n400), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(new_n416), .A4(new_n421), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n401), .A2(new_n406), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n418), .A2(new_n325), .A3(new_n419), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(G169), .B2(new_n415), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT18), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT77), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(new_n432), .A3(KEYINPUT18), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n429), .A2(new_n432), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT18), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n428), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n385), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G116), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n269), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n203), .A2(G33), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n265), .A2(new_n268), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n447), .B2(new_n444), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n244), .A2(new_n213), .B1(G20), .B2(new_n444), .ZN(new_n449));
  AOI21_X1  g0249(.A(G20), .B1(G33), .B2(G283), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n249), .A2(G97), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT87), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n452), .B1(new_n450), .B2(new_n451), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n449), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT20), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(KEYINPUT20), .B(new_n449), .C1(new_n453), .C2(new_n454), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n448), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT21), .ZN(new_n461));
  INV_X1    g0261(.A(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G1), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n282), .A2(KEYINPUT66), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT66), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G41), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT5), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n463), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(G270), .A3(new_n283), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT85), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n468), .B1(new_n286), .B2(KEYINPUT5), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n284), .B1(new_n474), .B2(new_n463), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(KEYINPUT85), .A3(G270), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT80), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n474), .A2(new_n478), .A3(G274), .A4(new_n463), .ZN(new_n479));
  OAI211_X1 g0279(.A(G274), .B(new_n463), .C1(new_n467), .C2(new_n469), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT80), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n351), .A2(new_n353), .A3(G264), .A4(G1698), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT86), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT86), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n275), .A2(new_n484), .A3(G264), .A4(G1698), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n359), .A2(G303), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n275), .A2(G257), .A3(new_n276), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n479), .A2(new_n481), .B1(new_n488), .B2(new_n284), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n461), .B(new_n301), .C1(new_n477), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n477), .A2(new_n489), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n325), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n460), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n460), .B1(new_n491), .B2(G200), .ZN(new_n494));
  INV_X1    g0294(.A(G190), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(new_n491), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT88), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n301), .B1(new_n477), .B2(new_n489), .ZN(new_n498));
  AOI211_X1 g0298(.A(new_n497), .B(KEYINPUT21), .C1(new_n498), .C2(new_n460), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT85), .B1(new_n475), .B2(G270), .ZN(new_n500));
  AND4_X1   g0300(.A1(KEYINPUT85), .A2(new_n470), .A3(G270), .A4(new_n283), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n481), .A2(new_n479), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n488), .A2(new_n284), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G169), .B(new_n460), .C1(new_n502), .C2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT88), .B1(new_n506), .B2(new_n461), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n493), .B(new_n496), .C1(new_n499), .C2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n351), .A2(new_n353), .A3(new_n204), .A4(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT22), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n275), .A2(new_n511), .A3(new_n204), .A4(G87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G20), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT89), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT23), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G107), .ZN(new_n519));
  NAND2_X1  g0319(.A1(KEYINPUT89), .A2(KEYINPUT23), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n518), .A2(G20), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n516), .B(new_n517), .C1(new_n204), .C2(G107), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n513), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT24), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n513), .A2(KEYINPUT24), .A3(new_n523), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n245), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n447), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT25), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n268), .B2(G107), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n269), .A2(KEYINPUT25), .A3(new_n519), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n529), .A2(G107), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n470), .A2(G264), .A3(new_n283), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT90), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT90), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n475), .A2(new_n537), .A3(G264), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n275), .A2(G250), .A3(new_n276), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n275), .A2(G257), .A3(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G294), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n284), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n536), .A2(new_n503), .A3(new_n538), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n312), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n481), .A2(new_n479), .B1(new_n284), .B2(new_n542), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(new_n495), .A3(new_n535), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n534), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n503), .A2(new_n535), .A3(new_n543), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G169), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n546), .A2(G179), .A3(new_n536), .A4(new_n538), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n550), .A2(new_n551), .B1(new_n528), .B2(new_n533), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT6), .ZN(new_n554));
  INV_X1    g0354(.A(G97), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n554), .A2(new_n555), .A3(G107), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n554), .B2(new_n238), .ZN(new_n557));
  OAI22_X1  g0357(.A1(new_n557), .A2(new_n204), .B1(new_n316), .B2(new_n251), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n519), .B1(new_n387), .B2(new_n388), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n245), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n268), .A2(G97), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n529), .B2(G97), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT81), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n481), .A2(new_n479), .B1(new_n475), .B2(G257), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n351), .A2(new_n353), .A3(G244), .A4(new_n276), .ZN(new_n566));
  XNOR2_X1  g0366(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g0368(.A1(KEYINPUT78), .A2(KEYINPUT4), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n275), .A2(G244), .A3(new_n276), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G283), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n275), .A2(G250), .A3(G1698), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n568), .A2(new_n570), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT79), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n573), .A2(new_n574), .A3(new_n284), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n573), .B2(new_n284), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n325), .B(new_n565), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n573), .A2(new_n284), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n475), .A2(G257), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n503), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n301), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT81), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n560), .A2(new_n582), .A3(new_n562), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n564), .A2(new_n577), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n580), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n563), .B1(new_n585), .B2(G190), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n565), .B1(new_n575), .B2(new_n576), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G200), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n275), .A2(G244), .A3(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n351), .A2(new_n353), .A3(G238), .A4(new_n276), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n514), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n284), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n203), .A2(G45), .ZN(new_n594));
  INV_X1    g0394(.A(G274), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT82), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT82), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n463), .A2(new_n597), .A3(G274), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n283), .A2(G250), .A3(new_n594), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G200), .ZN(new_n604));
  INV_X1    g0404(.A(G87), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n447), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n606), .B(KEYINPUT84), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT19), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n254), .B2(new_n555), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT83), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n275), .A2(new_n204), .A3(G68), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n204), .B1(new_n278), .B2(new_n608), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n605), .A2(new_n555), .A3(new_n519), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT83), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(new_n608), .C1(new_n254), .C2(new_n555), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n610), .A2(new_n611), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n617), .A2(new_n245), .B1(new_n269), .B2(new_n370), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n593), .A2(new_n602), .A3(G190), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n604), .A2(new_n607), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n529), .A2(new_n379), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n603), .A2(new_n301), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n601), .B1(new_n284), .B2(new_n592), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n325), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n553), .A2(new_n584), .A3(new_n589), .A4(new_n627), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n443), .A2(new_n508), .A3(new_n628), .ZN(G372));
  NAND2_X1  g0429(.A1(new_n348), .A2(new_n349), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n428), .A2(new_n313), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT92), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n382), .B1(new_n366), .B2(new_n301), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n632), .B1(new_n633), .B2(new_n368), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n375), .B1(new_n383), .B2(G169), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n362), .A2(new_n325), .A3(new_n365), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n635), .A2(new_n636), .A3(KEYINPUT92), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n309), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n631), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n438), .B1(new_n425), .B2(new_n431), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n435), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n630), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n341), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n623), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT91), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n647), .A2(new_n648), .B1(new_n618), .B2(new_n621), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n623), .A2(KEYINPUT91), .B1(new_n325), .B2(new_n624), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n528), .A2(new_n533), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n537), .B1(new_n475), .B2(G264), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n537), .A2(new_n470), .A3(G264), .A4(new_n283), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(G200), .B1(new_n655), .B2(new_n546), .ZN(new_n656));
  INV_X1    g0456(.A(new_n547), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AND4_X1   g0458(.A1(new_n584), .A2(new_n589), .A3(new_n658), .A4(new_n620), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n550), .A2(new_n551), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n534), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n493), .B(new_n661), .C1(new_n499), .C2(new_n507), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n651), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n620), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n649), .B2(new_n650), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n577), .A2(new_n581), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n665), .A2(new_n666), .A3(new_n668), .A4(new_n563), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n620), .A2(new_n626), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT26), .B1(new_n584), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n663), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n646), .B1(new_n442), .B2(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT93), .Z(G369));
  INV_X1    g0475(.A(G330), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n677));
  OAI21_X1  g0477(.A(G213), .B1(new_n677), .B2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT94), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT94), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n459), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n508), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n493), .B1(new_n499), .B2(new_n507), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n687), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n676), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n534), .A2(new_n685), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n553), .A2(new_n692), .B1(new_n552), .B2(new_n685), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n661), .A2(new_n685), .ZN(new_n696));
  AOI211_X1 g0496(.A(new_n301), .B(new_n459), .C1(new_n477), .C2(new_n489), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n497), .B1(new_n697), .B2(KEYINPUT21), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n506), .A2(KEYINPUT88), .A3(new_n461), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n685), .B1(new_n700), .B2(new_n493), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n696), .B1(new_n701), .B2(new_n553), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n695), .A2(new_n702), .ZN(G399));
  NOR2_X1   g0503(.A1(new_n207), .A2(new_n286), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n613), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n211), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n673), .A2(new_n710), .A3(new_n686), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n584), .A2(new_n670), .A3(KEYINPUT26), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n665), .A2(new_n668), .A3(new_n563), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(KEYINPUT26), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n685), .B1(new_n663), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n711), .B1(new_n710), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n536), .A2(new_n624), .A3(new_n538), .A4(new_n543), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT95), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n543), .A2(new_n593), .A3(new_n602), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n655), .A2(KEYINPUT95), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n585), .A2(G179), .A3(new_n477), .A4(new_n489), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n717), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n491), .A2(new_n325), .A3(new_n580), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(KEYINPUT30), .A3(new_n720), .A4(new_n722), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n624), .A2(G179), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n587), .A2(new_n491), .A3(new_n544), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT96), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n725), .A2(new_n727), .A3(KEYINPUT96), .A4(new_n729), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(new_n685), .A3(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n628), .A2(new_n508), .A3(new_n685), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n676), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n716), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n709), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n206), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n203), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n704), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n691), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n688), .A2(new_n676), .A3(new_n690), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT97), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n688), .A2(new_n690), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n208), .A2(new_n275), .ZN(new_n752));
  INV_X1    g0552(.A(G355), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n752), .A2(new_n753), .B1(G116), .B2(new_n208), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n242), .A2(new_n462), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n208), .A2(new_n359), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n462), .B2(new_n212), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n754), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n213), .B1(G20), .B2(new_n301), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n749), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n745), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n204), .A2(new_n495), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n312), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G87), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n325), .A2(new_n312), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n204), .A2(G190), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n767), .B1(new_n256), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n763), .A2(new_n768), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n359), .B(new_n772), .C1(G50), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  OAI21_X1  g0577(.A(KEYINPUT32), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n776), .A2(KEYINPUT32), .A3(new_n777), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n204), .B1(new_n775), .B2(G190), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n555), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n325), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n763), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G58), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n769), .A2(new_n764), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n784), .A2(new_n785), .B1(new_n786), .B2(new_n519), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n769), .A2(new_n783), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(G77), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n774), .A2(new_n778), .A3(new_n782), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n359), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT33), .B(G317), .Z(new_n794));
  NOR2_X1   g0594(.A1(new_n771), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n776), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n793), .B(new_n795), .C1(G329), .C2(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n766), .A2(G303), .B1(new_n773), .B2(G326), .ZN(new_n798));
  INV_X1    g0598(.A(new_n784), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G322), .A2(new_n799), .B1(new_n789), .B2(G311), .ZN(new_n800));
  INV_X1    g0600(.A(new_n780), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G294), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n797), .A2(new_n798), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n791), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n762), .B1(new_n804), .B2(new_n759), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n751), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n748), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n759), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT98), .Z(new_n811));
  INV_X1    g0611(.A(new_n786), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G87), .A2(new_n812), .B1(new_n796), .B2(G311), .ZN(new_n813));
  INV_X1    g0613(.A(G303), .ZN(new_n814));
  INV_X1    g0614(.A(new_n773), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n813), .B1(new_n519), .B2(new_n765), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n359), .B1(new_n784), .B2(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n771), .A2(new_n792), .B1(new_n788), .B2(new_n444), .ZN(new_n819));
  NOR4_X1   g0619(.A1(new_n816), .A2(new_n781), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G143), .A2(new_n799), .B1(new_n770), .B2(G150), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n822), .B2(new_n815), .C1(new_n777), .C2(new_n788), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT34), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n275), .B1(new_n776), .B2(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n765), .A2(new_n252), .B1(new_n786), .B2(new_n256), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(G58), .C2(new_n801), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n820), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n759), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n745), .B1(G77), .B2(new_n811), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n685), .A2(new_n375), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n634), .B2(new_n637), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT99), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n376), .A2(new_n384), .A3(new_n832), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT92), .B1(new_n635), .B2(new_n636), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n367), .A2(new_n632), .A3(new_n368), .A4(new_n375), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n832), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n376), .A2(new_n384), .A3(new_n832), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT99), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n831), .B1(new_n843), .B2(new_n809), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT100), .Z(new_n845));
  AOI21_X1  g0645(.A(new_n685), .B1(new_n663), .B2(new_n672), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(new_n843), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n847), .A2(new_n739), .B1(new_n704), .B2(new_n744), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n847), .A2(new_n739), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(G384));
  INV_X1    g0650(.A(new_n557), .ZN(new_n851));
  OAI211_X1 g0651(.A(G116), .B(new_n214), .C1(new_n851), .C2(KEYINPUT35), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(KEYINPUT35), .B2(new_n851), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT36), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n211), .A2(new_n390), .A3(new_n316), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n856), .A2(KEYINPUT101), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n856), .A2(KEYINPUT101), .B1(new_n252), .B2(G68), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n203), .B(G13), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT40), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n422), .B1(new_n425), .B2(new_n431), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n425), .A2(new_n683), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT37), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n429), .A2(new_n682), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n437), .A2(new_n865), .A3(new_n866), .A4(new_n422), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n425), .A2(new_n438), .A3(new_n431), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n641), .B1(new_n869), .B2(KEYINPUT77), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n870), .A2(new_n439), .B1(new_n423), .B2(new_n427), .ZN(new_n871));
  OAI211_X1 g0671(.A(KEYINPUT38), .B(new_n868), .C1(new_n871), .C2(new_n865), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n428), .A2(new_n642), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n863), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n868), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT103), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT103), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n878), .B(KEYINPUT38), .C1(new_n874), .C2(new_n868), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n872), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT102), .B1(new_n311), .B2(new_n686), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT102), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n274), .A2(new_n882), .A3(new_n685), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n309), .A2(new_n313), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n274), .B(new_n685), .C1(new_n304), .C2(new_n308), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n843), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n686), .B1(new_n730), .B2(new_n731), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(KEYINPUT31), .A3(new_n733), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n888), .B1(new_n737), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n861), .B1(new_n880), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n870), .A2(new_n439), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n865), .B1(new_n893), .B2(new_n428), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n864), .A2(new_n867), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n876), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT40), .B1(new_n896), .B2(new_n872), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(new_n891), .ZN(new_n898));
  OAI21_X1  g0698(.A(G330), .B1(new_n892), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n737), .A2(new_n890), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(G330), .A3(new_n442), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n863), .A2(new_n873), .B1(new_n864), .B2(new_n867), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n878), .B1(new_n903), .B2(KEYINPUT38), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n865), .B1(new_n428), .B2(new_n642), .ZN(new_n905));
  OAI211_X1 g0705(.A(KEYINPUT103), .B(new_n876), .C1(new_n895), .C2(new_n905), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n441), .A2(new_n863), .B1(new_n864), .B2(new_n867), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n904), .A2(new_n906), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n843), .B1(new_n884), .B2(new_n885), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n658), .A2(new_n661), .A3(new_n627), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n589), .A2(new_n584), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n491), .A2(G169), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n913), .A2(new_n461), .B1(new_n325), .B2(new_n491), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n698), .A2(new_n699), .B1(new_n914), .B2(new_n460), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n912), .A2(new_n915), .A3(new_n496), .A4(new_n686), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n916), .A2(KEYINPUT31), .B1(new_n889), .B2(new_n733), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n889), .A2(KEYINPUT31), .A3(new_n733), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n909), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT40), .B1(new_n908), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n897), .A2(new_n891), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n442), .A3(new_n900), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n902), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n646), .B1(new_n716), .B2(new_n442), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n924), .B(new_n925), .Z(new_n926));
  OR2_X1    g0726(.A1(new_n309), .A2(new_n685), .ZN(new_n927));
  XOR2_X1   g0727(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n928));
  OAI211_X1 g0728(.A(new_n872), .B(new_n928), .C1(new_n877), .C2(new_n879), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n441), .A2(new_n863), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n930), .B2(new_n868), .ZN(new_n931));
  INV_X1    g0731(.A(new_n872), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT39), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n927), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n673), .A2(new_n686), .A3(new_n887), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n376), .A2(new_n685), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n896), .A2(new_n872), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(new_n886), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n642), .A2(new_n682), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n934), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT105), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n926), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n203), .B2(new_n742), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n926), .A2(new_n945), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n860), .B1(new_n947), .B2(new_n948), .ZN(G367));
  XNOR2_X1  g0749(.A(new_n704), .B(KEYINPUT41), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n693), .B1(new_n915), .B2(new_n685), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n689), .A2(new_n553), .A3(new_n686), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n695), .B1(new_n691), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n740), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT108), .ZN(new_n957));
  INV_X1    g0757(.A(new_n696), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n563), .A2(new_n685), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n589), .A2(new_n584), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n667), .B2(new_n960), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n957), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  AOI211_X1 g0764(.A(KEYINPUT108), .B(new_n962), .C1(new_n952), .C2(new_n958), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n702), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n967), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n959), .B2(new_n963), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n966), .A2(KEYINPUT44), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n964), .B2(new_n965), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n971), .A2(KEYINPUT110), .A3(new_n695), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT108), .B1(new_n702), .B2(new_n962), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n959), .A2(new_n957), .A3(new_n963), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(KEYINPUT44), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n968), .A2(new_n970), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n973), .A2(new_n977), .A3(new_n695), .A4(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT110), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n956), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n740), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n950), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n743), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n584), .B1(new_n963), .B2(new_n661), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n686), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT42), .B1(new_n952), .B2(new_n911), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n952), .A2(KEYINPUT42), .A3(new_n911), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT106), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n686), .B1(new_n607), .B2(new_n618), .ZN(new_n992));
  MUX2_X1   g0792(.A(new_n665), .B(new_n651), .S(new_n992), .Z(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT106), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n987), .A2(new_n995), .A3(new_n989), .A4(new_n988), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n991), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n991), .A2(new_n996), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n993), .B(KEYINPUT43), .Z(new_n999));
  OAI221_X1 g0799(.A(new_n997), .B1(new_n695), .B2(new_n963), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n695), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n997), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n999), .B1(new_n991), .B2(new_n996), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1001), .B(new_n962), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n985), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n750), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n993), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n235), .A2(new_n756), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n760), .B1(new_n208), .B2(new_n370), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n745), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n765), .A2(new_n785), .B1(new_n788), .B2(new_n252), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n359), .B(new_n1013), .C1(G159), .C2(new_n770), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n786), .A2(new_n316), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n784), .A2(new_n335), .B1(new_n776), .B2(new_n822), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(G143), .C2(new_n773), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1014), .B(new_n1017), .C1(new_n256), .C2(new_n780), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n555), .A2(new_n786), .B1(new_n788), .B2(new_n792), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n275), .B(new_n1019), .C1(G303), .C2(new_n799), .ZN(new_n1020));
  INV_X1    g0820(.A(G311), .ZN(new_n1021));
  INV_X1    g0821(.A(G317), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n815), .A2(new_n1021), .B1(new_n776), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G294), .B2(new_n770), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n766), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT46), .B1(new_n766), .B2(G116), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G107), .B2(new_n801), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1020), .A2(new_n1024), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(KEYINPUT47), .B1(new_n1018), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1029), .A2(new_n830), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1018), .A2(new_n1028), .A3(KEYINPUT47), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1012), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1009), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1007), .A2(new_n1033), .ZN(G387));
  INV_X1    g0834(.A(KEYINPUT114), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n740), .B2(new_n955), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n954), .B(KEYINPUT114), .C1(new_n716), .C2(new_n739), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1036), .A2(new_n704), .A3(new_n956), .A4(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(KEYINPUT113), .B(G322), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n773), .A2(new_n1039), .B1(new_n770), .B2(G311), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n814), .B2(new_n788), .C1(new_n1022), .C2(new_n784), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT48), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n792), .B2(new_n780), .C1(new_n817), .C2(new_n765), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT49), .Z(new_n1044));
  AOI21_X1  g0844(.A(new_n275), .B1(new_n796), .B2(G326), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n444), .B2(new_n786), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n773), .A2(G159), .B1(new_n796), .B2(G150), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n275), .C1(new_n555), .C2(new_n786), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n771), .A2(new_n336), .B1(new_n252), .B2(new_n784), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n765), .A2(new_n316), .B1(new_n788), .B2(new_n256), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n780), .A2(new_n370), .ZN(new_n1052));
  NOR4_X1   g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n759), .B1(new_n1047), .B2(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n752), .A2(new_n706), .B1(G107), .B2(new_n208), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n232), .A2(G45), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n706), .B(new_n462), .C1(new_n256), .C2(new_n316), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n336), .A2(G50), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n756), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1055), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n745), .B1(new_n1063), .B2(new_n761), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT112), .Z(new_n1065));
  NAND2_X1  g0865(.A1(new_n1054), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n693), .B2(new_n750), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n744), .B2(new_n955), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1038), .A2(new_n1068), .ZN(G393));
  NAND2_X1  g0869(.A1(new_n971), .A2(new_n973), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n974), .A2(new_n981), .B1(new_n1070), .B2(new_n1001), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n963), .A2(new_n749), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n239), .A2(new_n756), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n760), .B1(new_n208), .B2(new_n555), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n745), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n815), .A2(new_n1022), .B1(new_n784), .B2(new_n1021), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT116), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1077), .B(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G303), .A2(new_n770), .B1(new_n796), .B2(new_n1039), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n792), .B2(new_n765), .C1(new_n817), .C2(new_n788), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n359), .B1(new_n780), .B2(new_n444), .C1(new_n519), .C2(new_n786), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n799), .A2(G159), .B1(new_n773), .B2(G150), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT51), .ZN(new_n1085));
  INV_X1    g0885(.A(G143), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n788), .A2(new_n336), .B1(new_n776), .B2(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n771), .A2(new_n252), .B1(new_n256), .B2(new_n765), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n275), .B1(new_n780), .B2(new_n316), .C1(new_n605), .C2(new_n786), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1083), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1075), .B1(new_n1091), .B2(new_n759), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1071), .A2(new_n744), .B1(new_n1072), .B2(new_n1092), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n982), .A2(new_n705), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n956), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1071), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1093), .B1(new_n1094), .B2(new_n1096), .ZN(G390));
  OAI211_X1 g0897(.A(G330), .B(new_n887), .C1(new_n917), .C2(new_n918), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n739), .B(new_n909), .C1(new_n1098), .C2(KEYINPUT117), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n685), .B(new_n843), .C1(new_n663), .C2(new_n714), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n886), .B1(new_n1100), .B2(new_n936), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n880), .A3(new_n927), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n929), .A2(new_n933), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n927), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n938), .B2(new_n886), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1099), .B(new_n1102), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n908), .A2(new_n928), .B1(KEYINPUT39), .B2(new_n939), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n936), .B1(new_n846), .B2(new_n887), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n886), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n927), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n904), .A2(new_n906), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1104), .B1(new_n1111), .B2(new_n872), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1107), .A2(new_n1110), .B1(new_n1101), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n676), .B1(new_n737), .B2(new_n890), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(KEYINPUT117), .A3(new_n909), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1106), .B(new_n744), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n745), .B1(new_n811), .B2(new_n402), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n815), .A2(new_n1118), .B1(new_n786), .B2(new_n252), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n359), .B(new_n1119), .C1(G125), .C2(new_n796), .ZN(new_n1120));
  OAI21_X1  g0920(.A(KEYINPUT53), .B1(new_n765), .B2(new_n335), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n765), .A2(KEYINPUT53), .A3(new_n335), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G159), .B2(new_n801), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n784), .A2(new_n825), .B1(new_n788), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G137), .B2(new_n770), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .A4(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n784), .A2(new_n444), .B1(new_n780), .B2(new_n316), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT120), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n815), .A2(new_n792), .B1(new_n771), .B2(new_n519), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G97), .B2(new_n789), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n786), .A2(new_n256), .B1(new_n776), .B2(new_n817), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT119), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1131), .A2(new_n359), .A3(new_n767), .A4(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1127), .B1(new_n1129), .B2(new_n1134), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1135), .A2(KEYINPUT121), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n830), .B1(new_n1135), .B2(KEYINPUT121), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1117), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n809), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1138), .B1(new_n1103), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1116), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1106), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT118), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n901), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1114), .A2(KEYINPUT118), .A3(new_n442), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1144), .A2(new_n925), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n738), .ZN(new_n1147));
  OAI211_X1 g0947(.A(G330), .B(new_n887), .C1(new_n917), .C2(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1109), .A2(new_n1148), .B1(new_n1114), .B2(new_n909), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1100), .A2(new_n936), .ZN(new_n1150));
  OAI21_X1  g0950(.A(G330), .B1(new_n917), .B2(new_n1147), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n888), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n886), .B1(new_n1114), .B2(new_n887), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1149), .A2(new_n1108), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1146), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n705), .B1(new_n1142), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1102), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1115), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1159), .A2(new_n1106), .A3(new_n1154), .A4(new_n1146), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1141), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(G378));
  XNOR2_X1  g0962(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n339), .A2(new_n682), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n350), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n350), .A2(new_n1165), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1164), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1168), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n1166), .A3(new_n1163), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n809), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n810), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n745), .B1(G50), .B2(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n773), .A2(G116), .B1(new_n801), .B2(G68), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT122), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G77), .A2(new_n766), .B1(new_n796), .B2(G283), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n555), .B2(new_n771), .C1(new_n370), .C2(new_n788), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n275), .A2(new_n286), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n785), .B2(new_n786), .C1(new_n519), .C2(new_n784), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1177), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1180), .ZN(new_n1183));
  AOI21_X1  g0983(.A(G50), .B1(new_n249), .B2(new_n282), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1182), .A2(KEYINPUT58), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n1118), .A2(new_n784), .B1(new_n765), .B2(new_n1124), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT123), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n780), .A2(new_n335), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n773), .A2(G125), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n771), .A2(new_n825), .B1(new_n788), .B2(new_n822), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n812), .A2(G159), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n796), .C2(G124), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1185), .B1(KEYINPUT58), .B2(new_n1182), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1175), .B1(new_n1198), .B2(new_n759), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1173), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n944), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1172), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n922), .B2(G330), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n676), .B(new_n1172), .C1(new_n920), .C2(new_n921), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1202), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n899), .A2(new_n1172), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n922), .A2(G330), .A3(new_n1203), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n944), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1201), .B1(new_n1210), .B2(new_n744), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1146), .B1(new_n1142), .B2(new_n1155), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(KEYINPUT57), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n704), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1209), .A2(new_n1206), .B1(new_n1160), .B2(new_n1146), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT57), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1211), .B1(new_n1214), .B2(new_n1216), .ZN(G375));
  NAND2_X1  g1017(.A1(new_n1109), .A2(new_n809), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n745), .B1(new_n811), .B2(G68), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n555), .A2(new_n765), .B1(new_n784), .B2(new_n792), .ZN(new_n1220));
  OR4_X1    g1020(.A1(new_n275), .A2(new_n1220), .A3(new_n1015), .A4(new_n1052), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G116), .A2(new_n770), .B1(new_n796), .B2(G303), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n519), .B2(new_n788), .C1(new_n817), .C2(new_n815), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G150), .A2(new_n789), .B1(new_n796), .B2(G128), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n777), .B2(new_n765), .C1(new_n771), .C2(new_n1124), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n799), .A2(G137), .B1(new_n773), .B2(G132), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n359), .B1(new_n812), .B2(G58), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n252), .C2(new_n780), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1221), .A2(new_n1223), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1219), .B1(new_n1229), .B2(new_n759), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1154), .A2(new_n744), .B1(new_n1218), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1155), .A2(new_n950), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1146), .A2(new_n1154), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1231), .B1(new_n1232), .B2(new_n1233), .ZN(G381));
  NAND2_X1  g1034(.A1(new_n1210), .A2(new_n744), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1200), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n705), .B1(new_n1215), .B2(KEYINPUT57), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT57), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1236), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1033), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n985), .B2(new_n1006), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1038), .A2(new_n1068), .A3(new_n807), .ZN(new_n1244));
  NOR4_X1   g1044(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1244), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1241), .A2(new_n1243), .A3(new_n1161), .A4(new_n1245), .ZN(G407));
  NAND2_X1  g1046(.A1(new_n1241), .A2(new_n1161), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G407), .B(G213), .C1(G343), .C2(new_n1247), .ZN(G409));
  NAND2_X1  g1048(.A1(new_n684), .A2(G213), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1210), .A2(new_n950), .A3(new_n1212), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1211), .A2(new_n1161), .A3(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1249), .B(new_n1251), .C1(new_n1241), .C2(new_n1161), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n684), .A2(G213), .A3(G2897), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT60), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1146), .B2(new_n1154), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1149), .A2(new_n1108), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1144), .A2(new_n925), .A3(new_n1145), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(KEYINPUT60), .A4(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1256), .A2(new_n1260), .A3(new_n704), .A4(new_n1155), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(G384), .A3(new_n1231), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G384), .B1(new_n1261), .B2(new_n1231), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1254), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1264), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(new_n1262), .A3(new_n1253), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT61), .B1(new_n1252), .B2(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1251), .A2(new_n1249), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1270), .B(new_n1271), .C1(new_n1161), .C2(new_n1241), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT62), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1251), .A2(new_n1249), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(G378), .B2(G375), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1271), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1269), .A2(new_n1273), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1243), .B2(G390), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G393), .A2(G396), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1244), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT125), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1281), .A2(new_n1284), .A3(new_n1244), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n974), .A2(new_n981), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1070), .A2(new_n1001), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n744), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1092), .A2(new_n1072), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1071), .A2(new_n1095), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n982), .A2(new_n705), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1005), .B1(new_n984), .B2(new_n743), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1294), .A2(new_n1295), .A3(new_n1242), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G390), .B1(new_n1007), .B2(new_n1033), .ZN(new_n1297));
  OAI22_X1  g1097(.A1(new_n1280), .A2(new_n1286), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G387), .A2(new_n1294), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1281), .A2(new_n1284), .A3(new_n1244), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1284), .B1(new_n1281), .B2(new_n1244), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1243), .A2(G390), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1299), .A2(new_n1279), .A3(new_n1302), .A4(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1278), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT124), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1307), .B1(new_n1275), .B2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1252), .A2(KEYINPUT124), .A3(new_n1268), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1275), .A2(KEYINPUT63), .A3(new_n1271), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT61), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1298), .A2(new_n1304), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1315), .B2(new_n1272), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1311), .A2(new_n1312), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1306), .A2(new_n1317), .ZN(G405));
  NAND2_X1  g1118(.A1(G375), .A2(G378), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1247), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1271), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1247), .A2(new_n1319), .A3(new_n1271), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT127), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1325), .A3(new_n1305), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1305), .A2(new_n1325), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1298), .A2(new_n1304), .A3(KEYINPUT127), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1322), .A2(new_n1327), .A3(new_n1328), .A4(new_n1323), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1326), .A2(new_n1329), .ZN(G402));
endmodule


