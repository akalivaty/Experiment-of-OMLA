//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT65), .B(G77), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n214), .A2(G244), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(G58), .A2(G68), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n225), .A2(G50), .A3(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n212), .B1(KEYINPUT1), .B2(new_n221), .C1(new_n223), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G50), .B(G68), .Z(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G1), .A2(G13), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(KEYINPUT68), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G50), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n207), .B1(new_n224), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n256), .A2(new_n259), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n253), .B1(new_n255), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n248), .B(new_n250), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n267), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n206), .A2(G20), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G50), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n264), .B1(G50), .B2(new_n267), .C1(new_n269), .C2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT9), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n278), .A3(G274), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n278), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n276), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n280), .B1(G226), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n289), .A2(G223), .B1(new_n214), .B2(new_n287), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT3), .B(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G222), .A3(new_n288), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n283), .B1(new_n293), .B2(new_n278), .ZN(new_n294));
  XOR2_X1   g0094(.A(new_n294), .B(KEYINPUT67), .Z(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n273), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n294), .B(KEYINPUT67), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT10), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n298), .A2(KEYINPUT70), .A3(new_n299), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT70), .B1(new_n298), .B2(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT69), .B(KEYINPUT10), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n273), .B(new_n305), .C1(new_n296), .C2(new_n295), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n301), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n298), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n272), .C1(G169), .C2(new_n298), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n284), .A2(new_n286), .A3(G232), .A4(G1698), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n284), .A2(new_n286), .A3(G226), .A4(new_n288), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n281), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT13), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n278), .A2(G238), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n279), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n317), .B1(new_n316), .B2(new_n321), .ZN(new_n323));
  OAI21_X1  g0123(.A(G200), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n258), .A2(G77), .ZN(new_n325));
  INV_X1    g0125(.A(G68), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n251), .A2(new_n252), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT73), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n249), .A2(new_n267), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n270), .A2(G68), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n265), .A2(new_n207), .A3(G1), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n248), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n335), .A2(KEYINPUT73), .A3(G68), .A4(new_n270), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n334), .A2(KEYINPUT12), .A3(new_n326), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT12), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n267), .B2(G68), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n339), .B(new_n341), .C1(new_n328), .C2(KEYINPUT11), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n324), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n316), .A2(new_n321), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT71), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n320), .B1(new_n281), .B2(new_n315), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n317), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n317), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT72), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n322), .A2(KEYINPUT72), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n350), .A2(G190), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n344), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT74), .B1(new_n338), .B2(new_n342), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n341), .A2(new_n339), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n327), .A2(new_n325), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n253), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT11), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT74), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(new_n329), .A4(new_n337), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  AND4_X1   g0165(.A1(G179), .A2(new_n350), .A3(new_n353), .A4(new_n354), .ZN(new_n366));
  OAI21_X1  g0166(.A(G169), .B1(new_n322), .B2(new_n323), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT14), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT14), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(G169), .C1(new_n322), .C2(new_n323), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n365), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n311), .A2(new_n356), .A3(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(G58), .A2(G68), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n374), .B2(new_n224), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n261), .A2(G159), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n375), .A2(KEYINPUT76), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT76), .B1(new_n375), .B2(new_n376), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n291), .B2(G20), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n287), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n326), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(KEYINPUT75), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT75), .ZN(new_n385));
  AOI211_X1 g0185(.A(new_n385), .B(new_n326), .C1(new_n381), .C2(new_n382), .ZN(new_n386));
  OAI211_X1 g0186(.A(KEYINPUT16), .B(new_n379), .C1(new_n384), .C2(new_n386), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n291), .A2(new_n380), .A3(G20), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT7), .B1(new_n287), .B2(new_n207), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n379), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n249), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n291), .A2(G226), .A3(G1698), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n291), .A2(G223), .A3(new_n288), .ZN(new_n396));
  INV_X1    g0196(.A(G87), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n395), .B(new_n396), .C1(new_n257), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n281), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n280), .B1(G232), .B2(new_n282), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n399), .A2(G190), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n299), .B1(new_n399), .B2(new_n400), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n256), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n270), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n269), .A2(new_n405), .B1(new_n267), .B2(new_n404), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n394), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n394), .A2(new_n407), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  INV_X1    g0212(.A(G169), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n399), .B2(new_n400), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n399), .A2(new_n400), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n308), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n411), .A2(new_n412), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n406), .B1(new_n387), .B2(new_n393), .ZN(new_n419));
  INV_X1    g0219(.A(new_n416), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n414), .B1(new_n420), .B2(G179), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT18), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(KEYINPUT17), .A3(new_n403), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n410), .A2(new_n418), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n289), .A2(G238), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n291), .A2(G232), .A3(new_n288), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n426), .B(new_n427), .C1(new_n203), .C2(new_n291), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n281), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n280), .B1(G244), .B2(new_n282), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G200), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT15), .B(G87), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n214), .A2(G20), .B1(new_n434), .B2(new_n258), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n404), .A2(new_n261), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n249), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n335), .A2(G77), .A3(new_n270), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n214), .B2(new_n267), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n432), .B(new_n440), .C1(new_n296), .C2(new_n431), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n440), .B1(new_n431), .B2(new_n413), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n429), .A2(new_n308), .A3(new_n430), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n425), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n373), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n284), .A2(new_n286), .A3(G264), .A4(G1698), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT85), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT85), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n291), .A2(new_n450), .A3(G264), .A4(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n287), .A2(G303), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n291), .A2(G257), .A3(new_n288), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n449), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n281), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(new_n274), .A3(KEYINPUT5), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(KEYINPUT79), .B2(G41), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n275), .A2(G1), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G270), .A3(new_n278), .ZN(new_n462));
  INV_X1    g0262(.A(G274), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n222), .B2(new_n277), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(new_n457), .A3(new_n459), .A4(new_n460), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n455), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT86), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n454), .B2(new_n281), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT86), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(G200), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT82), .ZN(new_n474));
  INV_X1    g0274(.A(G116), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(KEYINPUT82), .A2(G116), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(G20), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n479), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n248), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT20), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n266), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n475), .B1(new_n206), .B2(G33), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n485), .B1(new_n335), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n470), .B(KEYINPUT86), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n473), .B(new_n489), .C1(new_n490), .C2(new_n296), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n284), .A2(new_n286), .A3(new_n207), .A4(G87), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT22), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT22), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n291), .A2(new_n494), .A3(new_n207), .A4(G87), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n257), .B1(new_n476), .B2(new_n477), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n207), .A2(G107), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT23), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT23), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n207), .B2(G107), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n497), .A2(new_n207), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT24), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n496), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n249), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n266), .A2(new_n498), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(KEYINPUT87), .A3(KEYINPUT25), .ZN(new_n510));
  OR2_X1    g0310(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n511));
  NAND2_X1  g0311(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n266), .A2(new_n498), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n268), .B(new_n267), .C1(G1), .C2(new_n257), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n510), .B(new_n513), .C1(new_n514), .C2(new_n203), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n284), .A2(new_n286), .A3(G257), .A4(G1698), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n284), .A2(new_n286), .A3(G250), .A4(new_n288), .ZN(new_n518));
  XOR2_X1   g0318(.A(KEYINPUT88), .B(G294), .Z(new_n519));
  OAI211_X1 g0319(.A(new_n517), .B(new_n518), .C1(new_n519), .C2(new_n257), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n281), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n461), .A2(new_n278), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G264), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n521), .A2(new_n523), .A3(new_n465), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G190), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n281), .A2(new_n520), .B1(new_n522), .B2(G264), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n465), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G200), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n508), .A2(new_n516), .A3(new_n525), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n491), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n413), .B1(new_n483), .B2(new_n487), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n469), .A2(new_n472), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT21), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI211_X1 g0334(.A(new_n308), .B(new_n466), .C1(new_n281), .C2(new_n454), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n488), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n469), .A2(KEYINPUT21), .A3(new_n472), .A4(new_n531), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n527), .A2(new_n413), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n524), .A2(new_n308), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n538), .B(new_n539), .C1(new_n507), .C2(new_n515), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n534), .A2(new_n536), .A3(new_n537), .A4(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n530), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT84), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT83), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT81), .ZN(new_n545));
  AND2_X1   g0345(.A1(G244), .A2(G1698), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n291), .B2(new_n546), .ZN(new_n547));
  AND4_X1   g0347(.A1(new_n545), .A2(new_n284), .A3(new_n286), .A4(new_n546), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n284), .A2(new_n286), .A3(G238), .A4(new_n288), .ZN(new_n550));
  INV_X1    g0350(.A(new_n477), .ZN(new_n551));
  NOR2_X1   g0351(.A1(KEYINPUT82), .A2(G116), .ZN(new_n552));
  OAI21_X1  g0352(.A(G33), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n278), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n464), .A2(new_n460), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n206), .A2(G45), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n278), .A2(G250), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n544), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n284), .A2(new_n286), .A3(new_n546), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT81), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n291), .A2(new_n545), .A3(new_n546), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(new_n553), .A4(new_n550), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n559), .B1(new_n564), .B2(new_n281), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT83), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n299), .B1(new_n560), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n259), .B2(new_n202), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n291), .A2(new_n207), .A3(G68), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n207), .B1(new_n314), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G87), .B2(new_n204), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n248), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n433), .A2(new_n334), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n574), .B(new_n575), .C1(new_n514), .C2(new_n397), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n543), .B1(new_n567), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n576), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n565), .A2(KEYINPUT83), .ZN(new_n579));
  AOI211_X1 g0379(.A(new_n544), .B(new_n559), .C1(new_n564), .C2(new_n281), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(KEYINPUT84), .B(new_n578), .C1(new_n581), .C2(new_n299), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n560), .A2(G190), .A3(new_n566), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n577), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n560), .A2(new_n308), .A3(new_n566), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n574), .B(new_n575), .C1(new_n514), .C2(new_n433), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n585), .B(new_n586), .C1(new_n581), .C2(G169), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n284), .A2(new_n286), .A3(G250), .A4(G1698), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n284), .A2(new_n286), .A3(G244), .A4(new_n288), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n479), .B(new_n589), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT78), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n589), .A2(new_n479), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT78), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n590), .A2(new_n591), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n291), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n595), .A2(new_n596), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n278), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT80), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n461), .A2(new_n278), .ZN(new_n602));
  INV_X1    g0402(.A(G257), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n461), .A2(KEYINPUT80), .A3(G257), .A4(new_n278), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n465), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(G169), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n267), .A2(G97), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n514), .B2(new_n202), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT6), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n614), .A2(new_n202), .A3(G107), .ZN(new_n615));
  XNOR2_X1  g0415(.A(G97), .B(G107), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(G77), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n617), .A2(new_n207), .B1(new_n618), .B2(new_n262), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n203), .B1(new_n381), .B2(new_n382), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n248), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT77), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT77), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n623), .B(new_n248), .C1(new_n619), .C2(new_n620), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n613), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n600), .A2(new_n607), .A3(G179), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n594), .A2(new_n599), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n281), .ZN(new_n629));
  INV_X1    g0429(.A(new_n465), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n604), .B2(new_n605), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n296), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(G200), .B2(new_n608), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n610), .A2(new_n627), .B1(new_n633), .B2(new_n625), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n447), .A2(new_n542), .A3(new_n588), .A4(new_n634), .ZN(G372));
  NOR3_X1   g0435(.A1(new_n609), .A2(new_n625), .A3(new_n626), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n584), .A2(KEYINPUT26), .A3(new_n636), .A4(new_n587), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n627), .A2(new_n610), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n583), .B(new_n578), .C1(new_n299), .C2(new_n565), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n413), .B1(new_n555), .B2(new_n559), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n585), .A2(new_n586), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n638), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n541), .A2(KEYINPUT89), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n537), .A2(new_n536), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT89), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n647), .A2(new_n648), .A3(new_n534), .A4(new_n540), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n640), .A2(new_n642), .A3(new_n529), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n646), .A2(new_n649), .A3(new_n634), .A4(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n645), .A2(new_n651), .A3(new_n642), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n447), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n350), .A2(G179), .A3(new_n353), .A4(new_n354), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(new_n368), .A3(new_n370), .ZN(new_n655));
  INV_X1    g0455(.A(new_n444), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n365), .A2(new_n655), .B1(new_n656), .B2(new_n356), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n410), .A2(new_n423), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n418), .A2(new_n422), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n307), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n653), .A2(new_n310), .A3(new_n661), .ZN(G369));
  NAND2_X1  g0462(.A1(new_n647), .A2(new_n534), .ZN(new_n663));
  OR3_X1    g0463(.A1(new_n484), .A2(KEYINPUT27), .A3(G20), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT27), .B1(new_n484), .B2(G20), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n489), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n663), .B(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(new_n491), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  INV_X1    g0473(.A(new_n540), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n668), .B1(new_n507), .B2(new_n515), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n674), .B1(new_n529), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n540), .A2(new_n668), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n668), .B1(new_n647), .B2(new_n534), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n677), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n210), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G1), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n227), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n588), .A2(new_n638), .A3(new_n636), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n634), .A2(new_n650), .A3(new_n541), .ZN(new_n694));
  INV_X1    g0494(.A(new_n642), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n636), .A2(new_n642), .A3(new_n640), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(KEYINPUT26), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .A3(new_n669), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(KEYINPUT91), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n699), .A2(KEYINPUT91), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n652), .A2(new_n669), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n700), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n588), .A2(new_n542), .A3(new_n634), .A4(new_n669), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n669), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n565), .A2(G179), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n469), .A2(new_n472), .A3(new_n709), .A4(new_n527), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n535), .A2(new_n560), .A3(new_n526), .A4(new_n566), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n629), .A2(KEYINPUT30), .A3(new_n631), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n710), .A2(new_n608), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g0513(.A(KEYINPUT90), .B(KEYINPUT30), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n470), .A2(G179), .A3(new_n526), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n716), .A2(new_n579), .A3(new_n580), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n715), .B1(new_n717), .B2(new_n608), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n708), .B1(new_n713), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n608), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n629), .A2(new_n631), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n714), .B1(new_n711), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n490), .A2(new_n527), .A3(new_n721), .A4(new_n709), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT31), .B1(new_n724), .B2(new_n668), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n706), .A2(new_n719), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n705), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n692), .B1(new_n730), .B2(G1), .ZN(G364));
  NOR2_X1   g0531(.A1(new_n265), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n206), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n687), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n672), .B2(G330), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G330), .B2(new_n672), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT92), .Z(new_n738));
  INV_X1    g0538(.A(new_n735), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n210), .A2(G355), .A3(new_n291), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n686), .A2(new_n291), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G45), .B2(new_n227), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n241), .A2(new_n275), .ZN(new_n743));
  OAI221_X1 g0543(.A(new_n740), .B1(G116), .B2(new_n210), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n247), .B1(G20), .B2(new_n413), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n739), .B1(new_n744), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n748), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n207), .A2(G190), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(new_n308), .A3(new_n299), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT94), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT94), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G329), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT95), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n308), .B2(G200), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n299), .A2(KEYINPUT95), .A3(G179), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n207), .A2(new_n296), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G303), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n756), .A2(new_n757), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n752), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n761), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n308), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n763), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n291), .B1(new_n774), .B2(G322), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n752), .A2(new_n772), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G190), .ZN(new_n780));
  INV_X1    g0580(.A(G317), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n781), .A2(KEYINPUT33), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(KEYINPUT33), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n779), .A2(new_n296), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT96), .B(G326), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n296), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n207), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n784), .B1(new_n786), .B2(new_n787), .C1(new_n519), .C2(new_n789), .ZN(new_n790));
  NOR4_X1   g0590(.A1(new_n766), .A2(new_n771), .A3(new_n778), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n764), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n792), .A2(G87), .B1(G107), .B2(new_n768), .ZN(new_n793));
  INV_X1    g0593(.A(new_n789), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G97), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n287), .B1(new_n780), .B2(G68), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT32), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n756), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n756), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n801), .A2(KEYINPUT32), .A3(G159), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n797), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n777), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n774), .A2(G58), .B1(new_n804), .B2(new_n214), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n254), .B2(new_n786), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT93), .Z(new_n807));
  AOI21_X1  g0607(.A(new_n791), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n747), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n750), .B1(new_n751), .B2(new_n808), .C1(new_n672), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n738), .A2(new_n810), .ZN(G396));
  NOR2_X1   g0611(.A1(new_n748), .A2(new_n745), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n739), .B1(new_n618), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n780), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n795), .B1(new_n814), .B2(new_n770), .C1(new_n765), .C2(new_n786), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n756), .A2(new_n776), .B1(new_n764), .B2(new_n203), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n769), .A2(new_n397), .ZN(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n476), .A2(new_n477), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n287), .B1(new_n773), .B2(new_n818), .C1(new_n820), .C2(new_n777), .ZN(new_n821));
  NOR4_X1   g0621(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G137), .A2(new_n785), .B1(new_n780), .B2(G150), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT97), .ZN(new_n824));
  INV_X1    g0624(.A(G143), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n825), .B2(new_n773), .C1(new_n799), .C2(new_n777), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT34), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n768), .A2(G68), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n254), .B2(new_n764), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n830), .A2(KEYINPUT98), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(KEYINPUT98), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n287), .B1(new_n794), .B2(G58), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n756), .B2(new_n834), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n822), .B1(new_n827), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n444), .A2(new_n668), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n441), .B1(new_n440), .B2(new_n669), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n839), .B2(new_n444), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n813), .B1(new_n837), .B2(new_n751), .C1(new_n840), .C2(new_n746), .ZN(new_n841));
  INV_X1    g0641(.A(new_n840), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n702), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n445), .A2(new_n669), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n652), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n735), .B1(new_n846), .B2(new_n728), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n846), .A2(new_n728), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n841), .B1(new_n848), .B2(new_n849), .ZN(G384));
  INV_X1    g0650(.A(KEYINPUT103), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n387), .A2(new_n253), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n390), .A2(new_n385), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n383), .A2(KEYINPUT75), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT16), .B1(new_n855), .B2(new_n379), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n407), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n666), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n424), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n857), .A2(new_n858), .B1(new_n419), .B2(new_n403), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n857), .A2(new_n417), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n408), .B1(new_n419), .B2(new_n421), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n419), .A2(new_n666), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n865), .A2(KEYINPUT37), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n860), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n860), .B(KEYINPUT38), .C1(new_n864), .C2(new_n867), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n357), .A2(new_n364), .A3(new_n668), .ZN(new_n873));
  AOI221_X4 g0673(.A(new_n873), .B1(new_n355), .B2(new_n344), .C1(new_n655), .C2(new_n365), .ZN(new_n874));
  INV_X1    g0674(.A(new_n873), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n372), .B2(new_n356), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n840), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT102), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n719), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n724), .A2(KEYINPUT102), .A3(new_n708), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n725), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n877), .B1(new_n881), .B2(new_n706), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n872), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n851), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI211_X1 g0685(.A(KEYINPUT103), .B(KEYINPUT40), .C1(new_n872), .C2(new_n882), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n865), .B2(new_n866), .ZN(new_n888));
  INV_X1    g0688(.A(new_n866), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n411), .A2(new_n417), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n889), .A2(new_n861), .A3(new_n890), .A4(new_n408), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n424), .A2(new_n866), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n869), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n884), .B1(new_n895), .B2(new_n871), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n887), .B1(new_n882), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n881), .A2(new_n706), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n373), .A2(new_n446), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(G330), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n897), .A2(new_n899), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n874), .A2(new_n876), .ZN(new_n905));
  INV_X1    g0705(.A(new_n838), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n845), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT101), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n845), .A2(KEYINPUT101), .A3(new_n906), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n872), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n660), .A2(new_n666), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT39), .B1(new_n895), .B2(new_n871), .ZN(new_n914));
  INV_X1    g0714(.A(new_n872), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(KEYINPUT39), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n372), .A2(new_n668), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(new_n913), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n661), .A2(new_n310), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n701), .A2(new_n704), .ZN(new_n921));
  INV_X1    g0721(.A(new_n700), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n920), .B1(new_n923), .B2(new_n447), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n919), .B(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n904), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n904), .A2(new_n925), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(new_n206), .C2(new_n732), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n616), .A2(new_n614), .ZN(new_n929));
  INV_X1    g0729(.A(new_n615), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n931), .A2(KEYINPUT35), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n932), .A2(new_n475), .A3(new_n223), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(KEYINPUT35), .B2(new_n931), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT99), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n936), .A2(KEYINPUT36), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(KEYINPUT36), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n213), .A2(new_n374), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n939), .A2(new_n227), .B1(G50), .B2(new_n326), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(G1), .A3(new_n265), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT100), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n928), .A2(new_n937), .A3(new_n938), .A4(new_n942), .ZN(G367));
  OAI21_X1  g0743(.A(new_n634), .B1(new_n625), .B2(new_n669), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(new_n540), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n668), .B1(new_n945), .B2(new_n639), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n944), .B1(new_n639), .B2(new_n669), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n683), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n948), .B2(KEYINPUT42), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n578), .A2(new_n669), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n643), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n695), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n949), .A2(new_n950), .B1(KEYINPUT43), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n955), .B(new_n956), .Z(new_n957));
  NAND2_X1  g0757(.A1(new_n680), .A2(new_n947), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n687), .B(KEYINPUT41), .Z(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n678), .B(new_n682), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n673), .B(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n684), .A2(new_n947), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n684), .A2(new_n947), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT45), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT104), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n680), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n970), .A3(new_n681), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n963), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n961), .B1(new_n974), .B2(new_n729), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n959), .B1(new_n975), .B2(new_n733), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n741), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n749), .B1(new_n210), .B2(new_n433), .C1(new_n978), .C2(new_n237), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n735), .ZN(new_n980));
  INV_X1    g0780(.A(G137), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n756), .A2(new_n981), .B1(new_n769), .B2(new_n213), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G58), .B2(new_n792), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n287), .B1(new_n774), .B2(G150), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n794), .A2(G68), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n984), .B(new_n985), .C1(new_n786), .C2(new_n825), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT107), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n804), .A2(G50), .B1(G159), .B2(new_n780), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n983), .B(new_n989), .C1(new_n987), .C2(new_n988), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n764), .A2(new_n820), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(KEYINPUT46), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n792), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n992), .B1(KEYINPUT106), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(KEYINPUT106), .B2(new_n993), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n769), .A2(new_n202), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G317), .B2(new_n801), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n789), .A2(new_n203), .B1(new_n770), .B2(new_n777), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT105), .Z(new_n999));
  OAI221_X1 g0799(.A(new_n287), .B1(new_n773), .B2(new_n765), .C1(new_n776), .C2(new_n786), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n519), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n780), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n997), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n990), .B1(new_n995), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n980), .B1(new_n1005), .B2(new_n748), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n952), .A2(new_n747), .A3(new_n953), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n977), .A2(new_n1008), .ZN(G387));
  INV_X1    g0809(.A(new_n963), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n730), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n729), .A2(new_n963), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1011), .A2(new_n687), .A3(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n678), .A2(new_n809), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n749), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n689), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1016), .A2(new_n210), .A3(new_n291), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(G107), .B2(new_n210), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n234), .A2(new_n275), .ZN(new_n1019));
  AOI211_X1 g0819(.A(G45), .B(new_n1016), .C1(G68), .C2(G77), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n256), .A2(G50), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n978), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1018), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n789), .A2(new_n433), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n404), .B2(new_n780), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n799), .B2(new_n786), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n756), .A2(new_n260), .B1(new_n764), .B2(new_n213), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n291), .B1(new_n777), .B2(new_n326), .C1(new_n254), .C2(new_n773), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n996), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G317), .A2(new_n774), .B1(new_n804), .B2(G303), .ZN(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT108), .B(G322), .Z(new_n1032));
  OAI221_X1 g0832(.A(new_n1031), .B1(new_n814), .B2(new_n776), .C1(new_n786), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT48), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n792), .A2(new_n1001), .B1(G283), .B2(new_n794), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n287), .B1(new_n769), .B2(new_n820), .C1(new_n787), .C2(new_n756), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1030), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n735), .B1(new_n1015), .B2(new_n1024), .C1(new_n1044), .C2(new_n751), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1013), .B1(new_n733), .B2(new_n963), .C1(new_n1014), .C2(new_n1045), .ZN(G393));
  OAI221_X1 g0846(.A(new_n749), .B1(new_n202), .B2(new_n210), .C1(new_n978), .C2(new_n244), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n735), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1032), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n801), .A2(new_n1049), .B1(G107), .B2(new_n768), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n786), .A2(new_n781), .B1(new_n773), .B2(new_n776), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT52), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n287), .B1(new_n777), .B2(new_n818), .C1(new_n814), .C2(new_n765), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n819), .B2(new_n794), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n792), .A2(G283), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1050), .A2(new_n1052), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n756), .A2(new_n825), .B1(new_n764), .B2(new_n326), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT109), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n291), .B1(new_n397), .B2(new_n769), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT110), .Z(new_n1061));
  AOI22_X1  g0861(.A1(new_n774), .A2(G159), .B1(G150), .B2(new_n785), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT51), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n794), .A2(G77), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n256), .B2(new_n777), .C1(new_n814), .C2(new_n254), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1056), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1048), .B1(new_n1067), .B2(new_n748), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n947), .B2(new_n809), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n972), .A2(new_n687), .A3(new_n973), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n1011), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n969), .B(new_n680), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1011), .A2(new_n687), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1072), .B1(new_n733), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(G390));
  OAI21_X1  g0876(.A(new_n1064), .B1(new_n786), .B2(new_n770), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n287), .B1(new_n777), .B2(new_n202), .C1(new_n475), .C2(new_n773), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n792), .B2(G87), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1079), .B(new_n828), .C1(new_n818), .C2(new_n756), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1077), .B(new_n1080), .C1(G107), .C2(new_n780), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT114), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(KEYINPUT54), .B(G143), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n789), .A2(new_n799), .B1(new_n1083), .B2(new_n777), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G137), .B2(new_n780), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT112), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT53), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n792), .B2(G150), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n774), .A2(G132), .B1(G128), .B2(new_n785), .ZN(new_n1089));
  INV_X1    g0889(.A(G125), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1089), .B1(new_n756), .B2(new_n1090), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n764), .A2(KEYINPUT53), .A3(new_n260), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n287), .B1(new_n768), .B2(G50), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT113), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1086), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n748), .B1(new_n1082), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n812), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n735), .C1(new_n404), .C2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n916), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n745), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n911), .B2(new_n917), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n905), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n727), .A2(G330), .A3(new_n840), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n895), .A2(new_n871), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n917), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n839), .A2(new_n444), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n698), .A2(new_n669), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n906), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n1110), .B2(new_n1103), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1102), .A2(new_n1104), .A3(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n898), .A2(new_n902), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n840), .A3(new_n1103), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT101), .B1(new_n845), .B2(new_n906), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n908), .B(new_n838), .C1(new_n652), .C2(new_n844), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1103), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n916), .B1(new_n1119), .B2(new_n1106), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1116), .B1(new_n1120), .B2(new_n1111), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1113), .A2(new_n1121), .A3(KEYINPUT111), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT111), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1123), .B(new_n1116), .C1(new_n1120), .C2(new_n1111), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1101), .B1(new_n1125), .B2(new_n734), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1126), .A2(KEYINPUT115), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(KEYINPUT115), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n447), .A2(new_n1114), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1114), .A2(new_n840), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n905), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1110), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1131), .A2(new_n1104), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n905), .B1(new_n728), .B2(new_n842), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1115), .A2(new_n1134), .B1(new_n909), .B2(new_n910), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n924), .B(new_n1129), .C1(new_n1133), .C2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1122), .A2(new_n1136), .A3(new_n1124), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n687), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1127), .A2(new_n1128), .B1(new_n1137), .B2(new_n1139), .ZN(G378));
  NAND2_X1  g0940(.A1(new_n924), .A2(new_n1129), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1124), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1102), .A2(new_n1112), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1123), .B1(new_n1144), .B2(new_n1116), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n1145), .B2(new_n1113), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1142), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT57), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n902), .B1(new_n896), .B2(new_n882), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n885), .B2(new_n886), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT118), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(KEYINPUT118), .B(new_n1150), .C1(new_n885), .C2(new_n886), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n272), .A2(new_n858), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n311), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n307), .A2(new_n310), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n272), .A3(new_n858), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1159), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1153), .A2(new_n1154), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n887), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1165), .A2(KEYINPUT118), .A3(new_n1162), .A4(new_n1150), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n919), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(new_n1166), .A3(new_n919), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1149), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n688), .B1(new_n1148), .B2(new_n1171), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1164), .A2(new_n1166), .A3(new_n919), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n919), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT119), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1136), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1141), .B1(new_n1125), .B2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1167), .A2(KEYINPUT119), .A3(new_n1168), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1172), .B1(new_n1180), .B2(KEYINPUT57), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1162), .A2(new_n745), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n735), .B1(G50), .B2(new_n1098), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n985), .B1(new_n814), .B2(new_n202), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n287), .A2(new_n274), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n773), .A2(new_n203), .B1(new_n777), .B2(new_n433), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n792), .C2(new_n214), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n768), .A2(G58), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n770), .C2(new_n756), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1185), .B(new_n1190), .C1(G116), .C2(new_n785), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT58), .Z(new_n1192));
  AOI22_X1  g0992(.A1(new_n804), .A2(G137), .B1(G125), .B2(new_n785), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n794), .A2(G150), .B1(G132), .B2(new_n780), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1083), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n792), .A2(new_n1195), .B1(G128), .B2(new_n774), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT116), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1193), .B(new_n1194), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n257), .B(new_n274), .C1(new_n769), .C2(new_n799), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G124), .B2(new_n801), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1186), .B(new_n254), .C1(G33), .C2(G41), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1192), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT117), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n751), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1184), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1182), .A2(new_n734), .B1(new_n1183), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1181), .A2(new_n1212), .ZN(G375));
  INV_X1    g1013(.A(new_n1147), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n905), .A2(new_n745), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n735), .B1(G68), .B2(new_n1098), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n801), .A2(G303), .B1(G77), .B2(new_n768), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n202), .B2(new_n764), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n291), .B(new_n1025), .C1(G283), .C2(new_n774), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n804), .A2(G107), .B1(new_n819), .B2(new_n780), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1220), .A2(KEYINPUT120), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(KEYINPUT120), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n785), .A2(G294), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1219), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n801), .A2(G128), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n291), .B1(new_n773), .B2(new_n981), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G150), .B2(new_n804), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n792), .A2(G159), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1225), .A2(new_n1189), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1195), .A2(new_n780), .B1(G132), .B2(new_n785), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n254), .B2(new_n789), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1218), .A2(new_n1224), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1216), .B1(new_n1232), .B2(new_n748), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT121), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1214), .A2(new_n734), .B1(new_n1215), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1136), .A2(new_n961), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(G381));
  NOR2_X1   g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1075), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(G387), .A2(new_n1240), .A3(G384), .A4(G381), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1126), .B1(new_n1139), .B2(new_n1137), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1241), .A2(new_n1181), .A3(new_n1212), .A4(new_n1243), .ZN(G407));
  NAND2_X1  g1044(.A1(new_n667), .A2(G213), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G407), .B(G213), .C1(G375), .C2(new_n1247), .ZN(G409));
  NAND3_X1  g1048(.A1(new_n977), .A2(G390), .A3(new_n1008), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1008), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1075), .B1(new_n976), .B2(new_n1250), .ZN(new_n1251));
  AND2_X1   g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1252), .A2(new_n1239), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1249), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1253), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT126), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1169), .A2(KEYINPUT119), .A3(new_n1170), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1148), .A2(new_n961), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1262), .A2(new_n734), .B1(new_n1183), .B2(new_n1211), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1243), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT122), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1181), .A2(G378), .A3(new_n1212), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1264), .A2(KEYINPUT122), .A3(new_n1243), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1245), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1246), .A2(G2897), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(KEYINPUT123), .B(new_n1136), .C1(new_n1237), .C2(KEYINPUT60), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT123), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT60), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(new_n1177), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n688), .B1(new_n1237), .B2(KEYINPUT60), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1274), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1279), .A2(G384), .A3(new_n1235), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G384), .B1(new_n1279), .B2(new_n1235), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1273), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(new_n1235), .ZN(new_n1283));
  INV_X1    g1083(.A(G384), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1279), .A2(G384), .A3(new_n1235), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n1286), .A3(new_n1272), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1282), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1271), .B2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1270), .A2(new_n1245), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT62), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1292), .A2(KEYINPUT62), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1258), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1280), .A2(new_n1281), .A3(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1270), .A2(new_n1245), .A3(new_n1298), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1255), .A2(new_n1256), .A3(KEYINPUT61), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT122), .B1(new_n1264), .B2(new_n1243), .ZN(new_n1302));
  AOI211_X1 g1102(.A(new_n1266), .B(new_n1242), .C1(new_n1261), .C2(new_n1263), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1246), .B1(new_n1304), .B2(new_n1268), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT124), .B1(new_n1305), .B2(new_n1288), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1292), .A2(new_n1297), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT124), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1271), .A2(new_n1308), .A3(new_n1289), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1301), .A2(new_n1306), .A3(new_n1307), .A4(new_n1309), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1310), .A2(KEYINPUT125), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT125), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1308), .B1(new_n1271), .B2(new_n1289), .ZN(new_n1313));
  AOI211_X1 g1113(.A(KEYINPUT124), .B(new_n1288), .C1(new_n1270), .C2(new_n1245), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT63), .B1(new_n1305), .B2(new_n1291), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1312), .B1(new_n1315), .B2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1296), .B1(new_n1311), .B2(new_n1319), .ZN(G405));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1243), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1268), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1291), .A2(KEYINPUT127), .ZN(new_n1323));
  XOR2_X1   g1123(.A(new_n1322), .B(new_n1323), .Z(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(new_n1258), .ZN(G402));
endmodule


