

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U558 ( .A1(n709), .A2(n538), .ZN(n537) );
  NOR2_X1 U559 ( .A1(G651), .A2(n584), .ZN(n814) );
  AND2_X1 U560 ( .A1(n548), .A2(n547), .ZN(n546) );
  NAND2_X1 U561 ( .A1(n546), .A2(n543), .ZN(n786) );
  NAND2_X1 U562 ( .A1(n545), .A2(n544), .ZN(n543) );
  BUF_X1 U563 ( .A(n640), .Z(n587) );
  XOR2_X1 U564 ( .A(KEYINPUT17), .B(n563), .Z(n903) );
  AND2_X1 U565 ( .A1(n1019), .A2(G1348), .ZN(n648) );
  INV_X1 U566 ( .A(n707), .ZN(n535) );
  NAND2_X1 U567 ( .A1(n707), .A2(KEYINPUT32), .ZN(n538) );
  OR2_X1 U568 ( .A1(n700), .A2(n538), .ZN(n536) );
  AND2_X1 U569 ( .A1(n553), .A2(n643), .ZN(n552) );
  INV_X1 U570 ( .A(KEYINPUT66), .ZN(n579) );
  OR2_X1 U571 ( .A1(n585), .A2(n584), .ZN(n580) );
  INV_X1 U572 ( .A(KEYINPUT28), .ZN(n678) );
  NAND2_X1 U573 ( .A1(n555), .A2(n524), .ZN(n554) );
  NAND2_X1 U574 ( .A1(n525), .A2(n523), .ZN(n555) );
  XNOR2_X1 U575 ( .A(KEYINPUT100), .B(KEYINPUT31), .ZN(n695) );
  AND2_X1 U576 ( .A1(n536), .A2(n534), .ZN(n533) );
  NAND2_X1 U577 ( .A1(n535), .A2(n708), .ZN(n534) );
  AND2_X1 U578 ( .A1(n700), .A2(n708), .ZN(n532) );
  AND2_X1 U579 ( .A1(n557), .A2(n733), .ZN(n718) );
  XNOR2_X1 U580 ( .A(n645), .B(n644), .ZN(n1019) );
  XNOR2_X1 U581 ( .A(n551), .B(KEYINPUT15), .ZN(n645) );
  NAND2_X1 U582 ( .A1(n552), .A2(n639), .ZN(n551) );
  AND2_X1 U583 ( .A1(n785), .A2(n529), .ZN(n547) );
  INV_X1 U584 ( .A(KEYINPUT106), .ZN(n544) );
  INV_X1 U585 ( .A(G543), .ZN(n556) );
  NOR2_X1 U586 ( .A1(n571), .A2(n570), .ZN(G160) );
  OR2_X1 U587 ( .A1(n668), .A2(n701), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n556), .B(KEYINPUT0), .ZN(n584) );
  AND2_X1 U589 ( .A1(n676), .A2(n561), .ZN(n524) );
  NOR2_X1 U590 ( .A1(n664), .A2(n663), .ZN(n525) );
  AND2_X1 U591 ( .A1(G92), .A2(n818), .ZN(n526) );
  OR2_X1 U592 ( .A1(KEYINPUT33), .A2(n727), .ZN(n527) );
  AND2_X1 U593 ( .A1(n537), .A2(n533), .ZN(n528) );
  XNOR2_X2 U594 ( .A(n567), .B(KEYINPUT65), .ZN(n743) );
  OR2_X1 U595 ( .A1(n771), .A2(KEYINPUT106), .ZN(n529) );
  NAND2_X1 U596 ( .A1(n701), .A2(G8), .ZN(n733) );
  AND2_X1 U597 ( .A1(G8), .A2(n711), .ZN(n530) );
  NAND2_X1 U598 ( .A1(n528), .A2(n531), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n709), .A2(n532), .ZN(n531) );
  NAND2_X1 U600 ( .A1(n542), .A2(n539), .ZN(n712) );
  NAND2_X1 U601 ( .A1(n541), .A2(n540), .ZN(n539) );
  NOR2_X1 U602 ( .A1(n710), .A2(n530), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n709), .B(KEYINPUT102), .ZN(n541) );
  INV_X1 U604 ( .A(n550), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n548) );
  AND2_X1 U606 ( .A1(n771), .A2(KEYINPUT106), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n736), .A2(n735), .ZN(n550) );
  NOR2_X1 U608 ( .A1(n642), .A2(n526), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n680), .A2(n554), .ZN(n682) );
  XNOR2_X1 U610 ( .A(n558), .B(KEYINPUT105), .ZN(n557) );
  NOR2_X1 U611 ( .A1(n719), .A2(n714), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n903), .A2(G138), .ZN(n559) );
  XOR2_X1 U613 ( .A(KEYINPUT64), .B(G2104), .Z(n560) );
  OR2_X1 U614 ( .A1(n1019), .A2(n675), .ZN(n561) );
  OR2_X1 U615 ( .A1(n733), .A2(n732), .ZN(n562) );
  XNOR2_X1 U616 ( .A(n669), .B(KEYINPUT27), .ZN(n672) );
  NOR2_X1 U617 ( .A1(n672), .A2(n671), .ZN(n677) );
  XNOR2_X1 U618 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U619 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U620 ( .A1(G1966), .A2(n733), .ZN(n710) );
  INV_X1 U621 ( .A(KEYINPUT32), .ZN(n708) );
  INV_X1 U622 ( .A(n1009), .ZN(n723) );
  NOR2_X1 U623 ( .A1(n724), .A2(n723), .ZN(n725) );
  AND2_X1 U624 ( .A1(n726), .A2(n725), .ZN(n727) );
  AND2_X1 U625 ( .A1(n999), .A2(n562), .ZN(n734) );
  NAND2_X1 U626 ( .A1(n819), .A2(G68), .ZN(n653) );
  NAND2_X1 U627 ( .A1(G160), .A2(G40), .ZN(n738) );
  INV_X1 U628 ( .A(KEYINPUT13), .ZN(n655) );
  XNOR2_X1 U629 ( .A(n656), .B(n655), .ZN(n659) );
  NOR2_X1 U630 ( .A1(n659), .A2(n658), .ZN(n661) );
  NOR2_X1 U631 ( .A1(G2105), .A2(G2104), .ZN(n563) );
  NAND2_X1 U632 ( .A1(n903), .A2(G137), .ZN(n566) );
  NOR2_X1 U633 ( .A1(G2105), .A2(n560), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G101), .A2(n574), .ZN(n564) );
  XOR2_X1 U635 ( .A(KEYINPUT23), .B(n564), .Z(n565) );
  NAND2_X1 U636 ( .A1(n566), .A2(n565), .ZN(n571) );
  AND2_X1 U637 ( .A1(G2105), .A2(G2104), .ZN(n899) );
  NAND2_X1 U638 ( .A1(G113), .A2(n899), .ZN(n569) );
  NAND2_X1 U639 ( .A1(n560), .A2(G2105), .ZN(n567) );
  NAND2_X1 U640 ( .A1(G125), .A2(n743), .ZN(n568) );
  NAND2_X1 U641 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U642 ( .A1(G126), .A2(n743), .ZN(n572) );
  XNOR2_X1 U643 ( .A(n572), .B(KEYINPUT90), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n559), .A2(n573), .ZN(n578) );
  NAND2_X1 U645 ( .A1(G114), .A2(n899), .ZN(n576) );
  BUF_X1 U646 ( .A(n574), .Z(n904) );
  NAND2_X1 U647 ( .A1(G102), .A2(n904), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X2 U649 ( .A1(n578), .A2(n577), .ZN(G164) );
  NOR2_X1 U650 ( .A1(G543), .A2(G651), .ZN(n818) );
  NAND2_X1 U651 ( .A1(G91), .A2(n818), .ZN(n582) );
  INV_X1 U652 ( .A(G651), .ZN(n585) );
  XNOR2_X2 U653 ( .A(n580), .B(n579), .ZN(n819) );
  NAND2_X1 U654 ( .A1(G78), .A2(n819), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U656 ( .A(KEYINPUT67), .B(n583), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G53), .A2(n814), .ZN(n589) );
  NOR2_X1 U658 ( .A1(G543), .A2(n585), .ZN(n586) );
  XOR2_X1 U659 ( .A(KEYINPUT1), .B(n586), .Z(n640) );
  NAND2_X1 U660 ( .A1(G65), .A2(n587), .ZN(n588) );
  AND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(G299) );
  NAND2_X1 U663 ( .A1(G52), .A2(n814), .ZN(n593) );
  NAND2_X1 U664 ( .A1(G64), .A2(n587), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n598) );
  NAND2_X1 U666 ( .A1(G90), .A2(n818), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G77), .A2(n819), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U669 ( .A(KEYINPUT9), .B(n596), .Z(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(G171) );
  INV_X1 U671 ( .A(KEYINPUT75), .ZN(n611) );
  NAND2_X1 U672 ( .A1(G51), .A2(n814), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G63), .A2(n587), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U675 ( .A(KEYINPUT6), .B(n601), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G76), .A2(n819), .ZN(n602) );
  XNOR2_X1 U677 ( .A(KEYINPUT74), .B(n602), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n818), .A2(G89), .ZN(n603) );
  XNOR2_X1 U679 ( .A(KEYINPUT4), .B(n603), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U681 ( .A(n606), .B(KEYINPUT5), .Z(n607) );
  NOR2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U683 ( .A(KEYINPUT7), .B(n609), .Z(n610) );
  XNOR2_X1 U684 ( .A(n611), .B(n610), .ZN(G168) );
  XOR2_X1 U685 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U686 ( .A1(G75), .A2(n819), .ZN(n614) );
  NAND2_X1 U687 ( .A1(G88), .A2(n818), .ZN(n612) );
  XOR2_X1 U688 ( .A(KEYINPUT83), .B(n612), .Z(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U690 ( .A1(G50), .A2(n814), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G62), .A2(n587), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U693 ( .A1(n618), .A2(n617), .ZN(G166) );
  INV_X1 U694 ( .A(G166), .ZN(G303) );
  NAND2_X1 U695 ( .A1(G86), .A2(n818), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G48), .A2(n814), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n819), .A2(G73), .ZN(n621) );
  XOR2_X1 U699 ( .A(KEYINPUT2), .B(n621), .Z(n622) );
  NOR2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n587), .A2(G61), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(G305) );
  NAND2_X1 U703 ( .A1(G87), .A2(n584), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n626), .B(KEYINPUT82), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G49), .A2(n814), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U708 ( .A1(n587), .A2(n629), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(G288) );
  AND2_X1 U710 ( .A1(G72), .A2(n819), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G85), .A2(n818), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G47), .A2(n814), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n587), .A2(G60), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(G290) );
  NOR2_X2 U717 ( .A1(G164), .A2(G1384), .ZN(n737) );
  INV_X1 U718 ( .A(n738), .ZN(n638) );
  NAND2_X2 U719 ( .A1(n737), .A2(n638), .ZN(n701) );
  INV_X1 U720 ( .A(n733), .ZN(n722) );
  NAND2_X1 U721 ( .A1(G54), .A2(n814), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n819), .A2(G79), .ZN(n639) );
  NAND2_X1 U723 ( .A1(G66), .A2(n640), .ZN(n641) );
  XNOR2_X1 U724 ( .A(KEYINPUT71), .B(n641), .ZN(n642) );
  INV_X1 U725 ( .A(KEYINPUT72), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G1341), .A2(KEYINPUT98), .ZN(n646) );
  NAND2_X1 U727 ( .A1(KEYINPUT26), .A2(n646), .ZN(n647) );
  NOR2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n649) );
  INV_X2 U729 ( .A(n701), .ZN(n684) );
  NOR2_X1 U730 ( .A1(n649), .A2(n684), .ZN(n664) );
  NOR2_X1 U731 ( .A1(G1341), .A2(KEYINPUT98), .ZN(n651) );
  NOR2_X1 U732 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n650) );
  OR2_X1 U733 ( .A1(n651), .A2(n650), .ZN(n662) );
  NAND2_X1 U734 ( .A1(n818), .A2(G81), .ZN(n652) );
  XNOR2_X1 U735 ( .A(n652), .B(KEYINPUT12), .ZN(n654) );
  NAND2_X1 U736 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U737 ( .A1(G56), .A2(n587), .ZN(n657) );
  XOR2_X1 U738 ( .A(KEYINPUT14), .B(n657), .Z(n658) );
  NAND2_X1 U739 ( .A1(n814), .A2(G43), .ZN(n660) );
  NAND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(n1010) );
  OR2_X1 U741 ( .A1(n662), .A2(n1010), .ZN(n663) );
  AND2_X1 U742 ( .A1(G2067), .A2(n1019), .ZN(n667) );
  NAND2_X1 U743 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n665) );
  NAND2_X1 U744 ( .A1(KEYINPUT98), .A2(n665), .ZN(n666) );
  NOR2_X1 U745 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n684), .A2(G2072), .ZN(n669) );
  NAND2_X1 U747 ( .A1(G1956), .A2(n701), .ZN(n670) );
  XNOR2_X1 U748 ( .A(KEYINPUT97), .B(n670), .ZN(n671) );
  INV_X1 U749 ( .A(G299), .ZN(n1002) );
  NAND2_X1 U750 ( .A1(n677), .A2(n1002), .ZN(n676) );
  NAND2_X1 U751 ( .A1(G1348), .A2(n701), .ZN(n674) );
  NAND2_X1 U752 ( .A1(G2067), .A2(n684), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U754 ( .A1(n677), .A2(n1002), .ZN(n679) );
  XNOR2_X1 U755 ( .A(n679), .B(n678), .ZN(n680) );
  XOR2_X1 U756 ( .A(KEYINPUT29), .B(KEYINPUT99), .Z(n681) );
  XNOR2_X1 U757 ( .A(n682), .B(n681), .ZN(n688) );
  OR2_X1 U758 ( .A1(n684), .A2(G1961), .ZN(n686) );
  XNOR2_X1 U759 ( .A(G2078), .B(KEYINPUT96), .ZN(n683) );
  XNOR2_X1 U760 ( .A(n683), .B(KEYINPUT25), .ZN(n974) );
  NAND2_X1 U761 ( .A1(n684), .A2(n974), .ZN(n685) );
  NAND2_X1 U762 ( .A1(n686), .A2(n685), .ZN(n689) );
  AND2_X1 U763 ( .A1(G171), .A2(n689), .ZN(n687) );
  NOR2_X1 U764 ( .A1(n688), .A2(n687), .ZN(n698) );
  NOR2_X1 U765 ( .A1(G171), .A2(n689), .ZN(n694) );
  NOR2_X1 U766 ( .A1(G2084), .A2(n701), .ZN(n711) );
  NOR2_X1 U767 ( .A1(n710), .A2(n711), .ZN(n690) );
  NAND2_X1 U768 ( .A1(G8), .A2(n690), .ZN(n691) );
  XNOR2_X1 U769 ( .A(KEYINPUT30), .B(n691), .ZN(n692) );
  NOR2_X1 U770 ( .A1(G168), .A2(n692), .ZN(n693) );
  NOR2_X1 U771 ( .A1(n694), .A2(n693), .ZN(n696) );
  XNOR2_X1 U772 ( .A(n699), .B(KEYINPUT101), .ZN(n709) );
  AND2_X1 U773 ( .A1(G286), .A2(G8), .ZN(n700) );
  INV_X1 U774 ( .A(G8), .ZN(n706) );
  NOR2_X1 U775 ( .A1(G1971), .A2(n733), .ZN(n703) );
  NOR2_X1 U776 ( .A1(G2090), .A2(n701), .ZN(n702) );
  NOR2_X1 U777 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U778 ( .A1(G303), .A2(n704), .ZN(n705) );
  OR2_X1 U779 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U780 ( .A(n712), .B(KEYINPUT103), .ZN(n719) );
  NAND2_X1 U781 ( .A1(G166), .A2(G8), .ZN(n713) );
  NOR2_X1 U782 ( .A1(G2090), .A2(n713), .ZN(n714) );
  NOR2_X1 U783 ( .A1(G1981), .A2(G305), .ZN(n715) );
  XOR2_X1 U784 ( .A(n715), .B(KEYINPUT24), .Z(n716) );
  NOR2_X1 U785 ( .A1(n733), .A2(n716), .ZN(n717) );
  NOR2_X1 U786 ( .A1(n718), .A2(n717), .ZN(n736) );
  INV_X1 U787 ( .A(n719), .ZN(n721) );
  NOR2_X1 U788 ( .A1(G1976), .A2(G288), .ZN(n1005) );
  NOR2_X1 U789 ( .A1(G1971), .A2(G303), .ZN(n1007) );
  NOR2_X1 U790 ( .A1(n1005), .A2(n1007), .ZN(n720) );
  NAND2_X1 U791 ( .A1(n721), .A2(n720), .ZN(n726) );
  NAND2_X1 U792 ( .A1(n722), .A2(KEYINPUT104), .ZN(n724) );
  NAND2_X1 U793 ( .A1(G1976), .A2(G288), .ZN(n1009) );
  XOR2_X1 U794 ( .A(G1981), .B(G305), .Z(n999) );
  INV_X1 U795 ( .A(KEYINPUT104), .ZN(n728) );
  NAND2_X1 U796 ( .A1(n728), .A2(n1005), .ZN(n731) );
  NAND2_X1 U797 ( .A1(n1005), .A2(KEYINPUT33), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n729), .A2(KEYINPUT104), .ZN(n730) );
  NAND2_X1 U799 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U800 ( .A1(n527), .A2(n734), .ZN(n735) );
  NOR2_X1 U801 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U802 ( .A(n739), .B(KEYINPUT91), .Z(n784) );
  INV_X1 U803 ( .A(n784), .ZN(n769) );
  XNOR2_X1 U804 ( .A(KEYINPUT37), .B(G2067), .ZN(n781) );
  NAND2_X1 U805 ( .A1(G140), .A2(n903), .ZN(n741) );
  NAND2_X1 U806 ( .A1(G104), .A2(n904), .ZN(n740) );
  NAND2_X1 U807 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U808 ( .A(KEYINPUT34), .B(n742), .ZN(n748) );
  NAND2_X1 U809 ( .A1(G116), .A2(n899), .ZN(n745) );
  NAND2_X1 U810 ( .A1(G128), .A2(n743), .ZN(n744) );
  NAND2_X1 U811 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U812 ( .A(n746), .B(KEYINPUT35), .Z(n747) );
  NOR2_X1 U813 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U814 ( .A(KEYINPUT36), .B(n749), .Z(n750) );
  XOR2_X1 U815 ( .A(KEYINPUT92), .B(n750), .Z(n923) );
  OR2_X1 U816 ( .A1(n781), .A2(n923), .ZN(n949) );
  NOR2_X1 U817 ( .A1(n769), .A2(n949), .ZN(n777) );
  XNOR2_X1 U818 ( .A(G1986), .B(G290), .ZN(n1016) );
  XOR2_X1 U819 ( .A(KEYINPUT94), .B(G1991), .Z(n983) );
  NAND2_X1 U820 ( .A1(G107), .A2(n899), .ZN(n752) );
  NAND2_X1 U821 ( .A1(G119), .A2(n743), .ZN(n751) );
  NAND2_X1 U822 ( .A1(n752), .A2(n751), .ZN(n756) );
  NAND2_X1 U823 ( .A1(G131), .A2(n903), .ZN(n754) );
  NAND2_X1 U824 ( .A1(G95), .A2(n904), .ZN(n753) );
  NAND2_X1 U825 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U826 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U827 ( .A(KEYINPUT93), .B(n757), .Z(n914) );
  NOR2_X1 U828 ( .A1(n983), .A2(n914), .ZN(n758) );
  XNOR2_X1 U829 ( .A(n758), .B(KEYINPUT95), .ZN(n767) );
  NAND2_X1 U830 ( .A1(G117), .A2(n899), .ZN(n760) );
  NAND2_X1 U831 ( .A1(G141), .A2(n903), .ZN(n759) );
  NAND2_X1 U832 ( .A1(n760), .A2(n759), .ZN(n763) );
  NAND2_X1 U833 ( .A1(n904), .A2(G105), .ZN(n761) );
  XOR2_X1 U834 ( .A(KEYINPUT38), .B(n761), .Z(n762) );
  NOR2_X1 U835 ( .A1(n763), .A2(n762), .ZN(n765) );
  NAND2_X1 U836 ( .A1(n743), .A2(G129), .ZN(n764) );
  NAND2_X1 U837 ( .A1(n765), .A2(n764), .ZN(n913) );
  NAND2_X1 U838 ( .A1(G1996), .A2(n913), .ZN(n766) );
  NAND2_X1 U839 ( .A1(n767), .A2(n766), .ZN(n957) );
  NOR2_X1 U840 ( .A1(n1016), .A2(n957), .ZN(n768) );
  NOR2_X1 U841 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U842 ( .A1(n777), .A2(n770), .ZN(n771) );
  NOR2_X1 U843 ( .A1(G1996), .A2(n913), .ZN(n963) );
  NOR2_X1 U844 ( .A1(G1986), .A2(G290), .ZN(n773) );
  NAND2_X1 U845 ( .A1(n983), .A2(n914), .ZN(n772) );
  XNOR2_X1 U846 ( .A(KEYINPUT107), .B(n772), .ZN(n958) );
  NOR2_X1 U847 ( .A1(n773), .A2(n958), .ZN(n774) );
  NOR2_X1 U848 ( .A1(n957), .A2(n774), .ZN(n775) );
  NOR2_X1 U849 ( .A1(n963), .A2(n775), .ZN(n776) );
  XNOR2_X1 U850 ( .A(n776), .B(KEYINPUT39), .ZN(n779) );
  INV_X1 U851 ( .A(n777), .ZN(n778) );
  NAND2_X1 U852 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U853 ( .A(n780), .B(KEYINPUT108), .ZN(n782) );
  NAND2_X1 U854 ( .A1(n923), .A2(n781), .ZN(n950) );
  NAND2_X1 U855 ( .A1(n782), .A2(n950), .ZN(n783) );
  NAND2_X1 U856 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U857 ( .A(n786), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U858 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U859 ( .A(G57), .ZN(G237) );
  INV_X1 U860 ( .A(G132), .ZN(G219) );
  INV_X1 U861 ( .A(G82), .ZN(G220) );
  NAND2_X1 U862 ( .A1(G7), .A2(G661), .ZN(n787) );
  XOR2_X1 U863 ( .A(n787), .B(KEYINPUT10), .Z(n948) );
  NAND2_X1 U864 ( .A1(n948), .A2(G567), .ZN(n788) );
  XOR2_X1 U865 ( .A(KEYINPUT11), .B(n788), .Z(G234) );
  INV_X1 U866 ( .A(G860), .ZN(n797) );
  OR2_X1 U867 ( .A1(n1010), .A2(n797), .ZN(n789) );
  XNOR2_X1 U868 ( .A(KEYINPUT68), .B(n789), .ZN(G153) );
  XNOR2_X1 U869 ( .A(G171), .B(KEYINPUT69), .ZN(G301) );
  INV_X1 U870 ( .A(n1019), .ZN(n926) );
  NOR2_X1 U871 ( .A1(G868), .A2(n926), .ZN(n790) );
  XNOR2_X1 U872 ( .A(KEYINPUT73), .B(n790), .ZN(n793) );
  NAND2_X1 U873 ( .A1(G868), .A2(G301), .ZN(n791) );
  XNOR2_X1 U874 ( .A(KEYINPUT70), .B(n791), .ZN(n792) );
  NAND2_X1 U875 ( .A1(n793), .A2(n792), .ZN(G284) );
  XOR2_X1 U876 ( .A(KEYINPUT76), .B(G868), .Z(n794) );
  NOR2_X1 U877 ( .A1(G286), .A2(n794), .ZN(n796) );
  NOR2_X1 U878 ( .A1(G868), .A2(G299), .ZN(n795) );
  NOR2_X1 U879 ( .A1(n796), .A2(n795), .ZN(G297) );
  NAND2_X1 U880 ( .A1(n797), .A2(G559), .ZN(n798) );
  NAND2_X1 U881 ( .A1(n798), .A2(n926), .ZN(n799) );
  XNOR2_X1 U882 ( .A(n799), .B(KEYINPUT77), .ZN(n800) );
  XOR2_X1 U883 ( .A(KEYINPUT16), .B(n800), .Z(G148) );
  NOR2_X1 U884 ( .A1(G868), .A2(n1010), .ZN(n803) );
  NAND2_X1 U885 ( .A1(n926), .A2(G868), .ZN(n801) );
  NOR2_X1 U886 ( .A1(G559), .A2(n801), .ZN(n802) );
  NOR2_X1 U887 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U888 ( .A(KEYINPUT78), .B(n804), .ZN(G282) );
  NAND2_X1 U889 ( .A1(G111), .A2(n899), .ZN(n806) );
  NAND2_X1 U890 ( .A1(G135), .A2(n903), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n806), .A2(n805), .ZN(n811) );
  NAND2_X1 U892 ( .A1(G123), .A2(n743), .ZN(n807) );
  XNOR2_X1 U893 ( .A(n807), .B(KEYINPUT18), .ZN(n809) );
  NAND2_X1 U894 ( .A1(n904), .A2(G99), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U896 ( .A1(n811), .A2(n810), .ZN(n956) );
  XNOR2_X1 U897 ( .A(G2096), .B(n956), .ZN(n812) );
  INV_X1 U898 ( .A(G2100), .ZN(n874) );
  NAND2_X1 U899 ( .A1(n812), .A2(n874), .ZN(G156) );
  NAND2_X1 U900 ( .A1(n926), .A2(G559), .ZN(n813) );
  XOR2_X1 U901 ( .A(n1010), .B(n813), .Z(n856) );
  NAND2_X1 U902 ( .A1(G55), .A2(n814), .ZN(n816) );
  NAND2_X1 U903 ( .A1(G67), .A2(n587), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U905 ( .A(KEYINPUT80), .B(n817), .ZN(n823) );
  NAND2_X1 U906 ( .A1(G93), .A2(n818), .ZN(n821) );
  NAND2_X1 U907 ( .A1(G80), .A2(n819), .ZN(n820) );
  NAND2_X1 U908 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U909 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U910 ( .A(KEYINPUT81), .B(n824), .Z(n859) );
  XOR2_X1 U911 ( .A(G299), .B(n859), .Z(n830) );
  XNOR2_X1 U912 ( .A(KEYINPUT19), .B(G305), .ZN(n825) );
  XNOR2_X1 U913 ( .A(n825), .B(G288), .ZN(n826) );
  XNOR2_X1 U914 ( .A(KEYINPUT84), .B(n826), .ZN(n828) );
  XOR2_X1 U915 ( .A(G290), .B(G303), .Z(n827) );
  XNOR2_X1 U916 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U917 ( .A(n830), .B(n829), .ZN(n929) );
  XNOR2_X1 U918 ( .A(n856), .B(n929), .ZN(n831) );
  XNOR2_X1 U919 ( .A(n831), .B(KEYINPUT85), .ZN(n832) );
  NAND2_X1 U920 ( .A1(n832), .A2(G868), .ZN(n833) );
  XNOR2_X1 U921 ( .A(n833), .B(KEYINPUT86), .ZN(n835) );
  OR2_X1 U922 ( .A1(G868), .A2(n859), .ZN(n834) );
  NAND2_X1 U923 ( .A1(n835), .A2(n834), .ZN(G295) );
  NAND2_X1 U924 ( .A1(G2084), .A2(G2078), .ZN(n836) );
  XOR2_X1 U925 ( .A(KEYINPUT20), .B(n836), .Z(n837) );
  NAND2_X1 U926 ( .A1(G2090), .A2(n837), .ZN(n838) );
  XNOR2_X1 U927 ( .A(KEYINPUT21), .B(n838), .ZN(n839) );
  NAND2_X1 U928 ( .A1(n839), .A2(G2072), .ZN(n840) );
  XOR2_X1 U929 ( .A(KEYINPUT87), .B(n840), .Z(G158) );
  XNOR2_X1 U930 ( .A(KEYINPUT88), .B(G44), .ZN(n841) );
  XNOR2_X1 U931 ( .A(n841), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U932 ( .A1(G220), .A2(G219), .ZN(n842) );
  XOR2_X1 U933 ( .A(KEYINPUT22), .B(n842), .Z(n843) );
  NOR2_X1 U934 ( .A1(G218), .A2(n843), .ZN(n844) );
  NAND2_X1 U935 ( .A1(G96), .A2(n844), .ZN(n854) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n854), .ZN(n848) );
  NAND2_X1 U937 ( .A1(G120), .A2(G108), .ZN(n845) );
  NOR2_X1 U938 ( .A1(G237), .A2(n845), .ZN(n846) );
  NAND2_X1 U939 ( .A1(G69), .A2(n846), .ZN(n855) );
  NAND2_X1 U940 ( .A1(G567), .A2(n855), .ZN(n847) );
  NAND2_X1 U941 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U942 ( .A(KEYINPUT89), .B(n849), .Z(n860) );
  NAND2_X1 U943 ( .A1(G661), .A2(G483), .ZN(n850) );
  NOR2_X1 U944 ( .A1(n860), .A2(n850), .ZN(n853) );
  NAND2_X1 U945 ( .A1(n853), .A2(G36), .ZN(G176) );
  NAND2_X1 U946 ( .A1(G2106), .A2(n948), .ZN(G217) );
  AND2_X1 U947 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U948 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U949 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U950 ( .A1(n853), .A2(n852), .ZN(G188) );
  XNOR2_X1 U951 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U953 ( .A(G120), .ZN(G236) );
  INV_X1 U954 ( .A(G96), .ZN(G221) );
  NOR2_X1 U955 ( .A1(n855), .A2(n854), .ZN(G325) );
  INV_X1 U956 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U957 ( .A(KEYINPUT79), .B(n856), .ZN(n857) );
  NOR2_X1 U958 ( .A1(G860), .A2(n857), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(G145) );
  INV_X1 U960 ( .A(n860), .ZN(G319) );
  XNOR2_X1 U961 ( .A(G1996), .B(KEYINPUT41), .ZN(n870) );
  XOR2_X1 U962 ( .A(G1976), .B(G1956), .Z(n862) );
  XNOR2_X1 U963 ( .A(G1991), .B(G1961), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U965 ( .A(G1981), .B(G1971), .Z(n864) );
  XNOR2_X1 U966 ( .A(G1986), .B(G1966), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U968 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U969 ( .A(KEYINPUT112), .B(G2474), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U971 ( .A(n870), .B(n869), .ZN(G229) );
  XNOR2_X1 U972 ( .A(G2067), .B(G2072), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n871), .B(KEYINPUT42), .ZN(n882) );
  XOR2_X1 U974 ( .A(G2678), .B(KEYINPUT43), .Z(n873) );
  XNOR2_X1 U975 ( .A(KEYINPUT110), .B(G2096), .ZN(n872) );
  XNOR2_X1 U976 ( .A(n873), .B(n872), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n874), .B(G2078), .ZN(n876) );
  XNOR2_X1 U978 ( .A(G2090), .B(G2084), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U980 ( .A(n878), .B(n877), .Z(n880) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(KEYINPUT109), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n882), .B(n881), .ZN(G227) );
  NAND2_X1 U984 ( .A1(G112), .A2(n899), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G136), .A2(n903), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n890) );
  NAND2_X1 U987 ( .A1(G124), .A2(n743), .ZN(n885) );
  XOR2_X1 U988 ( .A(KEYINPUT113), .B(n885), .Z(n886) );
  XNOR2_X1 U989 ( .A(n886), .B(KEYINPUT44), .ZN(n888) );
  NAND2_X1 U990 ( .A1(G100), .A2(n904), .ZN(n887) );
  NAND2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n889) );
  NOR2_X1 U992 ( .A1(n890), .A2(n889), .ZN(G162) );
  NAND2_X1 U993 ( .A1(G115), .A2(n899), .ZN(n892) );
  NAND2_X1 U994 ( .A1(G127), .A2(n743), .ZN(n891) );
  NAND2_X1 U995 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U996 ( .A(n893), .B(KEYINPUT47), .ZN(n895) );
  NAND2_X1 U997 ( .A1(G139), .A2(n903), .ZN(n894) );
  NAND2_X1 U998 ( .A1(n895), .A2(n894), .ZN(n898) );
  NAND2_X1 U999 ( .A1(G103), .A2(n904), .ZN(n896) );
  XNOR2_X1 U1000 ( .A(KEYINPUT117), .B(n896), .ZN(n897) );
  NOR2_X1 U1001 ( .A1(n898), .A2(n897), .ZN(n951) );
  NAND2_X1 U1002 ( .A1(G118), .A2(n899), .ZN(n901) );
  NAND2_X1 U1003 ( .A1(G130), .A2(n743), .ZN(n900) );
  NAND2_X1 U1004 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1005 ( .A(KEYINPUT114), .B(n902), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(G142), .A2(n903), .ZN(n906) );
  NAND2_X1 U1007 ( .A1(G106), .A2(n904), .ZN(n905) );
  NAND2_X1 U1008 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(KEYINPUT45), .B(n907), .ZN(n908) );
  XNOR2_X1 U1010 ( .A(KEYINPUT115), .B(n908), .ZN(n909) );
  NOR2_X1 U1011 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n951), .B(n911), .ZN(n922) );
  XOR2_X1 U1013 ( .A(G162), .B(n956), .Z(n912) );
  XNOR2_X1 U1014 ( .A(n913), .B(n912), .ZN(n918) );
  XOR2_X1 U1015 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n916) );
  XNOR2_X1 U1016 ( .A(n914), .B(KEYINPUT48), .ZN(n915) );
  XNOR2_X1 U1017 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1018 ( .A(n918), .B(n917), .Z(n920) );
  XNOR2_X1 U1019 ( .A(G164), .B(G160), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(n922), .B(n921), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(n924), .B(n923), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(G37), .A2(n925), .ZN(G395) );
  XNOR2_X1 U1024 ( .A(n1010), .B(G286), .ZN(n928) );
  XOR2_X1 U1025 ( .A(G171), .B(n926), .Z(n927) );
  XNOR2_X1 U1026 ( .A(n928), .B(n927), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(n930), .B(n929), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(G37), .A2(n931), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(KEYINPUT118), .B(n932), .ZN(G397) );
  XOR2_X1 U1030 ( .A(G2451), .B(G2430), .Z(n934) );
  XNOR2_X1 U1031 ( .A(G2438), .B(G2443), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(n934), .B(n933), .ZN(n940) );
  XOR2_X1 U1033 ( .A(G2435), .B(G2454), .Z(n936) );
  INV_X1 U1034 ( .A(G1348), .ZN(n1020) );
  XOR2_X1 U1035 ( .A(n1020), .B(G1341), .Z(n935) );
  XNOR2_X1 U1036 ( .A(n936), .B(n935), .ZN(n938) );
  XOR2_X1 U1037 ( .A(G2446), .B(G2427), .Z(n937) );
  XNOR2_X1 U1038 ( .A(n938), .B(n937), .ZN(n939) );
  XOR2_X1 U1039 ( .A(n940), .B(n939), .Z(n941) );
  NAND2_X1 U1040 ( .A1(G14), .A2(n941), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(G319), .A2(n947), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(G229), .A2(G227), .ZN(n942) );
  XNOR2_X1 U1043 ( .A(KEYINPUT49), .B(n942), .ZN(n943) );
  NOR2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(G395), .A2(G397), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(G225) );
  INV_X1 U1047 ( .A(G225), .ZN(G308) );
  INV_X1 U1048 ( .A(G69), .ZN(G235) );
  INV_X1 U1049 ( .A(n947), .ZN(G401) );
  INV_X1 U1050 ( .A(n948), .ZN(G223) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n970) );
  XOR2_X1 U1052 ( .A(G2072), .B(n951), .Z(n953) );
  XOR2_X1 U1053 ( .A(G164), .B(G2078), .Z(n952) );
  NOR2_X1 U1054 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1055 ( .A(KEYINPUT50), .B(n954), .ZN(n968) );
  XOR2_X1 U1056 ( .A(G2084), .B(G160), .Z(n955) );
  NOR2_X1 U1057 ( .A1(n956), .A2(n955), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n966) );
  XOR2_X1 U1060 ( .A(G2090), .B(G162), .Z(n961) );
  XNOR2_X1 U1061 ( .A(KEYINPUT120), .B(n961), .ZN(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1063 ( .A(KEYINPUT51), .B(n964), .ZN(n965) );
  NOR2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(KEYINPUT52), .B(n971), .ZN(n972) );
  INV_X1 U1068 ( .A(KEYINPUT55), .ZN(n994) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n994), .ZN(n973) );
  NAND2_X1 U1070 ( .A1(n973), .A2(G29), .ZN(n1056) );
  XOR2_X1 U1071 ( .A(G29), .B(KEYINPUT124), .Z(n997) );
  XNOR2_X1 U1072 ( .A(n974), .B(G27), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G2067), .B(G26), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(G2072), .B(G33), .ZN(n975) );
  NOR2_X1 U1075 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1076 ( .A1(G28), .A2(n977), .ZN(n980) );
  XNOR2_X1 U1077 ( .A(KEYINPUT122), .B(G1996), .ZN(n978) );
  XNOR2_X1 U1078 ( .A(G32), .B(n978), .ZN(n979) );
  NOR2_X1 U1079 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1080 ( .A1(n982), .A2(n981), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(KEYINPUT121), .B(n983), .ZN(n984) );
  XNOR2_X1 U1082 ( .A(G25), .B(n984), .ZN(n985) );
  NOR2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1084 ( .A(n987), .B(KEYINPUT53), .ZN(n988) );
  XNOR2_X1 U1085 ( .A(n988), .B(KEYINPUT123), .ZN(n991) );
  XOR2_X1 U1086 ( .A(G2084), .B(G34), .Z(n989) );
  XNOR2_X1 U1087 ( .A(KEYINPUT54), .B(n989), .ZN(n990) );
  NAND2_X1 U1088 ( .A1(n991), .A2(n990), .ZN(n993) );
  XNOR2_X1 U1089 ( .A(G35), .B(G2090), .ZN(n992) );
  NOR2_X1 U1090 ( .A1(n993), .A2(n992), .ZN(n995) );
  XOR2_X1 U1091 ( .A(n995), .B(n994), .Z(n996) );
  NAND2_X1 U1092 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1093 ( .A1(G11), .A2(n998), .ZN(n1054) );
  INV_X1 U1094 ( .A(G16), .ZN(n1050) );
  XOR2_X1 U1095 ( .A(n1050), .B(KEYINPUT56), .Z(n1027) );
  XNOR2_X1 U1096 ( .A(G1966), .B(G168), .ZN(n1000) );
  NAND2_X1 U1097 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1098 ( .A(n1001), .B(KEYINPUT57), .ZN(n1025) );
  XOR2_X1 U1099 ( .A(G171), .B(G1961), .Z(n1004) );
  XOR2_X1 U1100 ( .A(n1002), .B(G1956), .Z(n1003) );
  NOR2_X1 U1101 ( .A1(n1004), .A2(n1003), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(KEYINPUT126), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1103 ( .A1(n1007), .A2(n1006), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(G1971), .A2(G303), .ZN(n1008) );
  NAND2_X1 U1105 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XNOR2_X1 U1106 ( .A(G1341), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1107 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1108 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1109 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1110 ( .A1(n1018), .A2(n1017), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(n1020), .B(n1019), .ZN(n1021) );
  XNOR2_X1 U1112 ( .A(KEYINPUT125), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1052) );
  XOR2_X1 U1116 ( .A(G1986), .B(G24), .Z(n1031) );
  XNOR2_X1 U1117 ( .A(G1971), .B(G22), .ZN(n1029) );
  XNOR2_X1 U1118 ( .A(G23), .B(G1976), .ZN(n1028) );
  NOR2_X1 U1119 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1033) );
  XNOR2_X1 U1121 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n1032) );
  XNOR2_X1 U1122 ( .A(n1033), .B(n1032), .ZN(n1037) );
  XNOR2_X1 U1123 ( .A(G1966), .B(G21), .ZN(n1035) );
  XNOR2_X1 U1124 ( .A(G1961), .B(G5), .ZN(n1034) );
  NOR2_X1 U1125 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1126 ( .A1(n1037), .A2(n1036), .ZN(n1047) );
  XNOR2_X1 U1127 ( .A(KEYINPUT59), .B(G4), .ZN(n1038) );
  XOR2_X1 U1128 ( .A(n1038), .B(G1348), .Z(n1040) );
  XNOR2_X1 U1129 ( .A(G20), .B(G1956), .ZN(n1039) );
  NOR2_X1 U1130 ( .A1(n1040), .A2(n1039), .ZN(n1044) );
  XNOR2_X1 U1131 ( .A(G1341), .B(G19), .ZN(n1042) );
  XNOR2_X1 U1132 ( .A(G1981), .B(G6), .ZN(n1041) );
  NOR2_X1 U1133 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NAND2_X1 U1134 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XNOR2_X1 U1135 ( .A(KEYINPUT60), .B(n1045), .ZN(n1046) );
  NOR2_X1 U1136 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  XNOR2_X1 U1137 ( .A(KEYINPUT61), .B(n1048), .ZN(n1049) );
  NAND2_X1 U1138 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  NAND2_X1 U1139 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
  NOR2_X1 U1140 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
  NAND2_X1 U1141 ( .A1(n1056), .A2(n1055), .ZN(n1057) );
  XNOR2_X1 U1142 ( .A(KEYINPUT62), .B(n1057), .ZN(G150) );
  INV_X1 U1143 ( .A(G150), .ZN(G311) );
endmodule

