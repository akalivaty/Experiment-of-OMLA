//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n550, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n458), .A2(G125), .ZN(new_n459));
  AND2_X1   g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(KEYINPUT66), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n463), .A2(G2105), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G112), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n464), .A2(new_n466), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT67), .Z(new_n479));
  AOI211_X1 g054(.A(new_n474), .B(new_n479), .C1(G136), .C2(new_n467), .ZN(G162));
  INV_X1    g055(.A(G126), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G114), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  OAI22_X1  g059(.A1(new_n476), .A2(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n458), .A2(new_n486), .A3(G138), .A4(new_n482), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n475), .A2(G138), .A3(new_n482), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n489), .A2(KEYINPUT68), .A3(KEYINPUT4), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n485), .B1(new_n492), .B2(new_n493), .ZN(G164));
  NOR2_X1   g069(.A1(KEYINPUT5), .A2(G543), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n498), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT69), .B(G651), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n500), .B2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(new_n498), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G88), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT69), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT69), .A2(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT6), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n503), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n502), .A2(new_n507), .A3(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  INV_X1    g092(.A(G51), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n514), .A2(KEYINPUT70), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(KEYINPUT70), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n506), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n498), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n521), .A2(new_n526), .ZN(G168));
  NAND2_X1  g102(.A1(new_n519), .A2(new_n520), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n528), .A2(G52), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n506), .A2(G90), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n505), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n500), .B1(new_n533), .B2(new_n534), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n529), .A2(new_n537), .ZN(G171));
  NAND2_X1  g113(.A1(new_n528), .A2(G43), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT72), .B(G81), .Z(new_n540));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n505), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n506), .A2(new_n540), .B1(new_n543), .B2(new_n500), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  XOR2_X1   g124(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n550));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G188));
  INV_X1    g128(.A(KEYINPUT6), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT69), .ZN(new_n555));
  INV_X1    g130(.A(G651), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n554), .B1(new_n557), .B2(new_n509), .ZN(new_n558));
  OAI211_X1 g133(.A(G91), .B(new_n498), .C1(new_n558), .C2(new_n503), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT75), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n512), .A2(new_n513), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n561), .A2(new_n562), .A3(G91), .A4(new_n498), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n505), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n560), .A2(new_n563), .B1(G651), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n514), .A2(G53), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  NOR3_X1   g145(.A1(new_n504), .A2(new_n570), .A3(new_n508), .ZN(new_n571));
  INV_X1    g146(.A(new_n568), .ZN(new_n572));
  NOR2_X1   g147(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n569), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n567), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G168), .ZN(G286));
  NAND2_X1  g153(.A1(new_n506), .A2(G87), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n514), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n498), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n514), .A2(G48), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n561), .A2(G86), .A3(new_n498), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n497), .ZN(new_n586));
  OAI21_X1  g161(.A(G61), .B1(new_n586), .B2(new_n495), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(KEYINPUT76), .B1(G73), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n496), .B2(new_n497), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n501), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n585), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n501), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT77), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(G85), .B2(new_n506), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n528), .A2(G47), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(new_n506), .A2(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n528), .A2(G54), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n498), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n556), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n609), .B2(G171), .ZN(G284));
  OAI21_X1  g186(.A(new_n610), .B1(new_n609), .B2(G171), .ZN(G321));
  NAND2_X1  g187(.A1(G299), .A2(new_n609), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n609), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n609), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(new_n608), .ZN(new_n616));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n620), .B(KEYINPUT78), .C1(G868), .C2(new_n546), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(KEYINPUT78), .B2(new_n620), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n458), .A2(new_n468), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n467), .A2(G135), .ZN(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n482), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n631), .C1(new_n632), .C2(new_n476), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n628), .A2(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT80), .Z(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n651), .A3(G14), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT81), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT17), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(KEYINPUT18), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT82), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n662), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n671), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n671), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G35), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G162), .B2(new_n689), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT29), .Z(new_n692));
  INV_X1    g267(.A(G2090), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(KEYINPUT90), .B1(G16), .B2(G21), .ZN(new_n695));
  NAND2_X1  g270(.A1(G168), .A2(G16), .ZN(new_n696));
  MUX2_X1   g271(.A(KEYINPUT90), .B(new_n695), .S(new_n696), .Z(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT91), .B(G1966), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(G164), .A2(G29), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G27), .B2(G29), .ZN(new_n701));
  INV_X1    g276(.A(G2078), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n697), .A2(new_n698), .ZN(new_n704));
  NOR4_X1   g279(.A1(new_n694), .A2(new_n699), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n701), .A2(new_n702), .ZN(new_n706));
  NOR2_X1   g281(.A1(G4), .A2(G16), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n616), .B2(G16), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1348), .ZN(new_n709));
  AOI211_X1 g284(.A(new_n706), .B(new_n709), .C1(new_n693), .C2(new_n692), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n689), .A2(G32), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n468), .A2(G105), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT89), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(KEYINPUT89), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT26), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n714), .A2(new_n715), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n477), .A2(G129), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n467), .A2(G141), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n712), .B1(new_n724), .B2(new_n689), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT27), .B(G1996), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n633), .A2(new_n689), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT92), .Z(new_n729));
  INV_X1    g304(.A(G34), .ZN(new_n730));
  AOI21_X1  g305(.A(G29), .B1(new_n730), .B2(KEYINPUT24), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(KEYINPUT24), .B2(new_n730), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n470), .B2(new_n689), .ZN(new_n733));
  INV_X1    g308(.A(G2084), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n727), .A2(new_n729), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n689), .A2(G26), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT28), .Z(new_n739));
  INV_X1    g314(.A(G104), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n740), .A2(new_n482), .A3(KEYINPUT87), .ZN(new_n741));
  AOI21_X1  g316(.A(KEYINPUT87), .B1(new_n740), .B2(new_n482), .ZN(new_n742));
  OAI221_X1 g317(.A(G2104), .B1(G116), .B2(new_n482), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n467), .A2(G140), .ZN(new_n744));
  INV_X1    g319(.A(G128), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n743), .B(new_n744), .C1(new_n745), .C2(new_n476), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n739), .B1(new_n746), .B2(G29), .ZN(new_n747));
  INV_X1    g322(.A(G2067), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT30), .B(G28), .ZN(new_n750));
  OR2_X1    g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  NAND2_X1  g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n750), .A2(new_n689), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n725), .B2(new_n726), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n737), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G16), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G5), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G171), .B2(new_n756), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n756), .A2(G20), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT94), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT93), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT23), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G299), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1956), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n689), .A2(G33), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n467), .A2(G139), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n458), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n770), .B(new_n771), .C1(new_n482), .C2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT88), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n768), .B1(new_n774), .B2(new_n689), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(G2072), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n756), .A2(G19), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n546), .B2(new_n756), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G1341), .Z(new_n779));
  NAND4_X1  g354(.A1(new_n761), .A2(new_n767), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n711), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G6), .A2(G16), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n594), .B2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  INV_X1    g360(.A(G1981), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n756), .A2(G23), .ZN(new_n788));
  INV_X1    g363(.A(G288), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n756), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT33), .B(G1976), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G22), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G166), .B2(G16), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT85), .B(G1971), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n787), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT86), .Z(new_n798));
  INV_X1    g373(.A(KEYINPUT34), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  MUX2_X1   g376(.A(G24), .B(G290), .S(G16), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1986), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n689), .A2(G25), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n467), .A2(G131), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT83), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n808));
  INV_X1    g383(.A(G107), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G2105), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n477), .B2(G119), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n804), .B1(new_n813), .B2(new_n689), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT35), .B(G1991), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT84), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n803), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n800), .A2(new_n801), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n801), .A2(new_n819), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n822), .A2(new_n823), .A3(new_n800), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n782), .B1(new_n821), .B2(new_n824), .ZN(G311));
  NOR2_X1   g400(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n823), .B1(new_n822), .B2(new_n800), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n781), .B1(new_n826), .B2(new_n827), .ZN(G150));
  NOR2_X1   g403(.A1(new_n608), .A2(new_n617), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n528), .A2(G55), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n506), .A2(G93), .ZN(new_n833));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  INV_X1    g409(.A(G67), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n505), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n500), .B1(new_n836), .B2(new_n837), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n546), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n545), .B1(new_n832), .B2(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n831), .B(new_n844), .Z(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n841), .A2(new_n847), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  XNOR2_X1  g427(.A(new_n470), .B(KEYINPUT97), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n633), .ZN(new_n854));
  XNOR2_X1  g429(.A(G162), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n485), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n486), .B1(new_n467), .B2(G138), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n487), .B1(new_n857), .B2(KEYINPUT68), .ZN(new_n858));
  INV_X1    g433(.A(G138), .ZN(new_n859));
  AOI211_X1 g434(.A(new_n859), .B(G2105), .C1(new_n464), .C2(new_n466), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n860), .A2(new_n491), .A3(new_n486), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n856), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n746), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n723), .ZN(new_n864));
  INV_X1    g439(.A(new_n774), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n773), .B2(new_n864), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n812), .B(new_n626), .ZN(new_n868));
  OR2_X1    g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(G2104), .C1(G118), .C2(new_n482), .ZN(new_n870));
  INV_X1    g445(.A(G130), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n476), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(G142), .B2(new_n467), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n868), .B(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n867), .A2(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT98), .B1(new_n867), .B2(new_n874), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n855), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n855), .B(KEYINPUT99), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(new_n877), .ZN(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n882), .B2(new_n875), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g460(.A(new_n844), .B(new_n619), .ZN(new_n886));
  INV_X1    g461(.A(G299), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n608), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT101), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n886), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n886), .A2(new_n888), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G288), .B(KEYINPUT102), .ZN(new_n899));
  XNOR2_X1  g474(.A(G290), .B(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n594), .B(G303), .Z(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(KEYINPUT103), .B2(KEYINPUT42), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n898), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n898), .B2(new_n904), .ZN(new_n906));
  OAI21_X1  g481(.A(G868), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(G868), .B2(new_n841), .ZN(G295));
  OAI21_X1  g483(.A(new_n907), .B1(G868), .B2(new_n841), .ZN(G331));
  XOR2_X1   g484(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n891), .A2(new_n894), .ZN(new_n912));
  XNOR2_X1  g487(.A(G171), .B(G168), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n913), .A2(new_n844), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n844), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(KEYINPUT105), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n914), .A2(new_n888), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n912), .A2(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n919), .B2(new_n902), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n912), .A2(new_n916), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n917), .A2(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n902), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n911), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n921), .A2(new_n902), .A3(new_n922), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  INV_X1    g503(.A(new_n890), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n917), .A2(new_n914), .B1(new_n892), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n918), .A2(new_n915), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n924), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND4_X1   g507(.A1(new_n911), .A2(new_n927), .A3(new_n928), .A4(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n910), .B1(new_n926), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n927), .A2(new_n932), .A3(new_n928), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n920), .A2(new_n925), .A3(new_n911), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(G397));
  OAI21_X1  g514(.A(new_n491), .B1(new_n860), .B2(new_n486), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n493), .A3(new_n487), .ZN(new_n941));
  AOI21_X1  g516(.A(G1384), .B1(new_n941), .B2(new_n856), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(KEYINPUT45), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n461), .A2(G40), .A3(new_n469), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(G290), .A2(new_n945), .A3(G1986), .ZN(new_n946));
  AND2_X1   g521(.A1(G290), .A2(G1986), .ZN(new_n947));
  INV_X1    g522(.A(new_n945), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT106), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n723), .B(G1996), .Z(new_n951));
  XNOR2_X1  g526(.A(new_n746), .B(new_n748), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT107), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n813), .A2(new_n816), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n813), .A2(new_n816), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n948), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n950), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n961));
  INV_X1    g536(.A(new_n944), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n862), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n964), .B2(KEYINPUT50), .ZN(new_n965));
  AOI211_X1 g540(.A(KEYINPUT50), .B(G1384), .C1(new_n941), .C2(new_n856), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(G1348), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n862), .A2(new_n944), .A3(new_n963), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n942), .A2(KEYINPUT115), .A3(new_n944), .ZN(new_n972));
  AOI21_X1  g547(.A(G2067), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n961), .B1(new_n968), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n969), .A2(new_n970), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT115), .B1(new_n942), .B2(new_n944), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n748), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1348), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n944), .B1(new_n942), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n980), .B2(new_n966), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(KEYINPUT116), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n974), .A2(new_n616), .A3(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT113), .B(KEYINPUT57), .Z(new_n984));
  NOR4_X1   g559(.A1(new_n504), .A2(new_n570), .A3(new_n508), .A4(new_n572), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n574), .B1(new_n514), .B2(G53), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT114), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n567), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n575), .A2(KEYINPUT114), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(G1956), .B1(new_n965), .B2(new_n967), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(G164), .B2(G1384), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n862), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT56), .B(G2072), .ZN(new_n998));
  AND4_X1   g573(.A1(new_n996), .A2(new_n944), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n993), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT117), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1002), .B(new_n993), .C1(new_n994), .C2(new_n999), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n983), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1956), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n980), .B2(new_n966), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n962), .B1(new_n942), .B2(KEYINPUT45), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(new_n996), .A3(new_n998), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n992), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1009), .A2(KEYINPUT61), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1001), .A2(new_n1011), .A3(new_n1003), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n968), .A2(new_n973), .A3(new_n961), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT116), .B1(new_n977), .B2(new_n981), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT60), .B(new_n608), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1000), .A2(new_n1009), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT61), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT58), .B(G1341), .Z(new_n1019));
  NAND3_X1  g594(.A1(new_n971), .A2(new_n972), .A3(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT118), .B(G1996), .Z(new_n1021));
  NAND3_X1  g596(.A1(new_n1007), .A2(new_n996), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT59), .B1(new_n1023), .B2(new_n546), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n1025));
  AOI211_X1 g600(.A(new_n1025), .B(new_n545), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1012), .A2(new_n1015), .A3(new_n1018), .A4(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT60), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT60), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n974), .A2(new_n1030), .A3(new_n982), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1029), .A2(new_n616), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1010), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1007), .A2(KEYINPUT53), .A3(new_n996), .A4(new_n702), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1035), .A2(KEYINPUT121), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n965), .A2(new_n967), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n996), .A2(new_n702), .A3(new_n944), .A4(new_n997), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1037), .A2(new_n759), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1035), .A2(KEYINPUT121), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1036), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT122), .B1(new_n1042), .B2(G171), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1035), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G171), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1042), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1034), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n980), .A2(G2084), .A3(new_n966), .ZN(new_n1049));
  INV_X1    g624(.A(new_n698), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n1007), .B2(new_n996), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n521), .B2(new_n526), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT119), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1052), .B(new_n1055), .C1(KEYINPUT120), .C2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1054), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1007), .A2(new_n996), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n698), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n965), .A2(new_n734), .A3(new_n967), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1058), .B1(new_n1063), .B2(new_n1054), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT51), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1057), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n759), .B1(new_n980), .B2(new_n966), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(G301), .A3(new_n1069), .A4(new_n1035), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT54), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(G171), .B2(new_n1042), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1059), .B1(new_n942), .B2(new_n944), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n789), .A2(G1976), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1073), .B1(new_n1076), .B2(KEYINPUT52), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n1078));
  AOI211_X1 g653(.A(KEYINPUT109), .B(new_n1078), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n588), .A2(new_n592), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n500), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1082), .A2(new_n786), .A3(new_n584), .A4(new_n583), .ZN(new_n1083));
  OAI21_X1  g658(.A(G1981), .B1(new_n585), .B2(new_n593), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT49), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT49), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT110), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1074), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1093), .A2(new_n1074), .A3(new_n1085), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT110), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1076), .ZN(new_n1096));
  INV_X1    g671(.A(G1976), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(G288), .B2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1090), .A2(new_n1095), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n980), .A2(G2090), .A3(new_n966), .ZN(new_n1100));
  AOI21_X1  g675(.A(G1971), .B1(new_n1007), .B2(new_n996), .ZN(new_n1101));
  OAI21_X1  g676(.A(G8), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(G303), .A2(G8), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT55), .ZN(new_n1104));
  OR3_X1    g679(.A1(new_n1103), .A2(KEYINPUT108), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT108), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1102), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1108), .B(G8), .C1(new_n1101), .C2(new_n1100), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1080), .A2(new_n1099), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1067), .A2(new_n1072), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1033), .A2(new_n1048), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1099), .A2(new_n1080), .A3(new_n1110), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT112), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1080), .A2(new_n1099), .A3(new_n1110), .A4(KEYINPUT112), .ZN(new_n1118));
  AND4_X1   g693(.A1(KEYINPUT63), .A2(new_n1111), .A3(G168), .A4(new_n1063), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1063), .A2(G168), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1112), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT111), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1089), .B1(new_n1088), .B2(new_n1074), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1094), .A2(KEYINPUT110), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1128), .A2(new_n1111), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1074), .ZN(new_n1131));
  NOR2_X1   g706(.A1(G288), .A2(G1976), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1131), .B1(new_n1133), .B2(new_n1083), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1124), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1132), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1083), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1074), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1099), .A2(new_n1080), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1139), .B(KEYINPUT111), .C1(new_n1140), .C2(new_n1111), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1120), .A2(new_n1123), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1114), .A2(KEYINPUT123), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1067), .A2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1057), .B(KEYINPUT62), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1112), .A2(new_n1045), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT124), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1145), .A2(new_n1150), .A3(new_n1147), .A4(new_n1146), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1143), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT123), .B1(new_n1114), .B2(new_n1142), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n960), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n954), .A2(new_n957), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n746), .A2(G2067), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n945), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n945), .A2(G1996), .ZN(new_n1159));
  NAND2_X1  g734(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n952), .A2(new_n724), .ZN(new_n1162));
  OAI221_X1 g737(.A(new_n1161), .B1(KEYINPUT125), .B2(KEYINPUT46), .C1(new_n945), .C2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT47), .Z(new_n1164));
  INV_X1    g739(.A(new_n959), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n946), .B(KEYINPUT48), .Z(new_n1166));
  AOI211_X1 g741(.A(new_n1158), .B(new_n1164), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1155), .A2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g743(.A(G319), .ZN(new_n1170));
  NOR2_X1   g744(.A1(G227), .A2(new_n1170), .ZN(new_n1171));
  XOR2_X1   g745(.A(new_n1171), .B(KEYINPUT126), .Z(new_n1172));
  NOR3_X1   g746(.A1(G229), .A2(G401), .A3(new_n1172), .ZN(new_n1173));
  OAI211_X1 g747(.A(new_n884), .B(new_n1173), .C1(new_n926), .C2(new_n933), .ZN(G225));
  INV_X1    g748(.A(G225), .ZN(G308));
endmodule


