//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT85), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G148gat), .ZN(new_n205));
  INV_X1    g004(.A(G148gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G141gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT79), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT2), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(G155gat), .B(G162gat), .Z(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n213), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT3), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n218));
  INV_X1    g017(.A(G127gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(G134gat), .ZN(new_n220));
  INV_X1    g019(.A(G134gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G127gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G120gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G113gat), .ZN(new_n225));
  INV_X1    g024(.A(G113gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G120gat), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT1), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n221), .A2(G127gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(G134gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT70), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n223), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT71), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n220), .A2(new_n222), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n234), .A2(new_n228), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT71), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n223), .A2(new_n236), .A3(new_n228), .A4(new_n231), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n214), .A2(new_n215), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n217), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT81), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n217), .A2(new_n244), .A3(new_n238), .A4(new_n241), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n233), .A2(new_n235), .A3(new_n237), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT82), .ZN(new_n248));
  INV_X1    g047(.A(new_n213), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n212), .B(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT82), .B1(new_n238), .B2(new_n216), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G225gat), .A2(G233gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n238), .A2(new_n216), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(KEYINPUT4), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n246), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT83), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n238), .A2(new_n216), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n261), .B1(new_n263), .B2(new_n257), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n251), .A2(new_n252), .B1(new_n216), .B2(new_n238), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n265), .A2(KEYINPUT83), .A3(new_n256), .ZN(new_n266));
  OAI211_X1 g065(.A(KEYINPUT5), .B(new_n260), .C1(new_n264), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT4), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n254), .B1(new_n238), .B2(new_n216), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT84), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT84), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n272), .A3(new_n269), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n257), .A2(KEYINPUT5), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n271), .A2(new_n246), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G1gat), .B(G29gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT0), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(G57gat), .ZN(new_n279));
  INV_X1    g078(.A(G85gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n203), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n281), .B1(new_n267), .B2(new_n275), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n267), .A2(new_n281), .A3(new_n275), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n284), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n291));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(G183gat), .A3(G190gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT24), .ZN(new_n296));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT23), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT25), .B1(new_n300), .B2(G169gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(KEYINPUT23), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n298), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n298), .B(KEYINPUT64), .ZN(new_n306));
  INV_X1    g105(.A(new_n304), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT65), .B(G169gat), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n306), .B(new_n307), .C1(new_n308), .C2(new_n300), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT26), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n302), .A3(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n315), .A2(new_n295), .ZN(new_n316));
  AND2_X1   g115(.A1(KEYINPUT66), .A2(KEYINPUT27), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT66), .A2(KEYINPUT27), .ZN(new_n318));
  OAI21_X1  g117(.A(G183gat), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT67), .ZN(new_n320));
  INV_X1    g119(.A(G183gat), .ZN(new_n321));
  AOI211_X1 g120(.A(KEYINPUT28), .B(G190gat), .C1(new_n321), .C2(KEYINPUT27), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n323), .B(G183gat), .C1(new_n317), .C2(new_n318), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n326));
  XOR2_X1   g125(.A(KEYINPUT27), .B(G183gat), .Z(new_n327));
  OAI21_X1  g126(.A(KEYINPUT28), .B1(new_n327), .B2(G190gat), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n326), .B1(new_n325), .B2(new_n328), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n316), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT69), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(KEYINPUT69), .B(new_n316), .C1(new_n329), .C2(new_n330), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n311), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n292), .B1(new_n335), .B2(KEYINPUT29), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT76), .ZN(new_n337));
  XNOR2_X1  g136(.A(G197gat), .B(G204gat), .ZN(new_n338));
  INV_X1    g137(.A(G211gat), .ZN(new_n339));
  INV_X1    g138(.A(G218gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n338), .B1(KEYINPUT22), .B2(new_n341), .ZN(new_n342));
  XOR2_X1   g141(.A(G211gat), .B(G218gat), .Z(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n328), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT68), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n311), .B1(new_n349), .B2(new_n316), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n350), .A2(new_n292), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n352), .B(new_n292), .C1(new_n335), .C2(KEYINPUT29), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n337), .A2(new_n345), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n292), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n311), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT69), .B1(new_n349), .B2(new_n316), .ZN(new_n358));
  INV_X1    g157(.A(new_n334), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI221_X1 g159(.A(new_n344), .B1(new_n350), .B2(new_n356), .C1(new_n360), .C2(new_n292), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363));
  INV_X1    g162(.A(G64gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n365), .B(G92gat), .Z(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT78), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n369));
  AOI211_X1 g168(.A(new_n369), .B(new_n366), .C1(new_n354), .C2(new_n361), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n291), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n362), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n354), .A2(KEYINPUT77), .A3(new_n361), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n366), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n366), .B1(new_n354), .B2(new_n361), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT30), .ZN(new_n377));
  AND4_X1   g176(.A1(new_n290), .A2(new_n371), .A3(new_n375), .A4(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT35), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n344), .B1(new_n241), .B2(new_n355), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n216), .A2(new_n355), .A3(new_n344), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n217), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(G228gat), .A3(G233gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n385));
  OAI221_X1 g184(.A(new_n382), .B1(new_n250), .B2(new_n240), .C1(new_n380), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n381), .B2(KEYINPUT88), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n389), .A2(G50gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n389), .A2(G50gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393));
  INV_X1    g192(.A(G22gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  OR3_X1    g197(.A1(new_n391), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(new_n391), .B2(new_n392), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT74), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n360), .A2(new_n247), .ZN(new_n403));
  NAND2_X1  g202(.A1(G227gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n335), .A2(new_n238), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT32), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G15gat), .B(G43gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(G71gat), .ZN(new_n412));
  INV_X1    g211(.A(G99gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n408), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n414), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n407), .B(KEYINPUT32), .C1(new_n409), .C2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n402), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n415), .A2(new_n402), .A3(new_n417), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT34), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n335), .A2(new_n238), .ZN(new_n422));
  AOI211_X1 g221(.A(new_n247), .B(new_n311), .C1(new_n333), .C2(new_n334), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n421), .B(new_n404), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT73), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT34), .B1(new_n403), .B2(new_n406), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT73), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n404), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT72), .B1(new_n422), .B2(new_n423), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT72), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n403), .A2(new_n430), .A3(new_n406), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n404), .A3(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n425), .A2(new_n428), .B1(new_n432), .B2(KEYINPUT34), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n419), .A2(new_n420), .A3(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n415), .A2(new_n402), .A3(new_n417), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n425), .A2(new_n428), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(KEYINPUT34), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n435), .B1(new_n418), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n401), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n378), .A2(KEYINPUT90), .A3(new_n379), .A4(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n354), .A2(KEYINPUT77), .A3(new_n361), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT77), .B1(new_n354), .B2(new_n361), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n445), .A2(new_n366), .B1(new_n376), .B2(KEYINPUT30), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n446), .A2(new_n379), .A3(new_n290), .A4(new_n371), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n399), .A2(new_n400), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n435), .A2(new_n418), .A3(new_n438), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n415), .A2(new_n417), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n433), .A2(new_n450), .A3(KEYINPUT74), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n448), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n442), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n441), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n371), .A2(new_n290), .A3(new_n375), .A4(new_n377), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n446), .A2(KEYINPUT86), .A3(new_n290), .A4(new_n371), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n440), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n454), .B1(KEYINPUT35), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n271), .A2(new_n246), .A3(new_n273), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n257), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n462), .B(KEYINPUT39), .C1(new_n257), .C2(new_n263), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT39), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(new_n464), .A3(new_n257), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n465), .A2(new_n466), .A3(new_n281), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n466), .B1(new_n465), .B2(new_n281), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n286), .B1(new_n469), .B2(new_n470), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n362), .A2(new_n367), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n369), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n376), .A2(KEYINPUT78), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT30), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n375), .A2(new_n377), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n471), .B(new_n472), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n448), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n286), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT85), .B1(new_n286), .B2(KEYINPUT6), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n482), .B(new_n289), .C1(new_n368), .C2(new_n370), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n337), .A2(new_n351), .A3(new_n353), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n344), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n350), .A2(new_n356), .ZN(new_n486));
  INV_X1    g285(.A(new_n292), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(new_n335), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n485), .B(KEYINPUT37), .C1(new_n344), .C2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT37), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n362), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n366), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n373), .A2(KEYINPUT37), .A3(new_n374), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n495), .A2(KEYINPUT38), .A3(new_n366), .A4(new_n491), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n483), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n479), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n448), .B1(new_n457), .B2(new_n458), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT75), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT36), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n500), .A2(KEYINPUT36), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n501), .B(new_n502), .C1(new_n449), .C2(new_n451), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n434), .A2(new_n439), .A3(new_n500), .A4(KEYINPUT36), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n498), .A2(new_n499), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n202), .B1(new_n460), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT16), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(G1gat), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(G1gat), .B2(new_n508), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G8gat), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n512), .B(KEYINPUT94), .Z(new_n513));
  INV_X1    g312(.A(KEYINPUT95), .ZN(new_n514));
  AOI21_X1  g313(.A(G8gat), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n510), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT14), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT14), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT93), .ZN(new_n525));
  XOR2_X1   g324(.A(G43gat), .B(G50gat), .Z(new_n526));
  INV_X1    g325(.A(KEYINPUT15), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n526), .A2(new_n527), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n525), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n524), .B2(KEYINPUT92), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(KEYINPUT92), .B2(new_n524), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT17), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n513), .A2(new_n517), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n534), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n537), .B(new_n534), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n540), .B(KEYINPUT13), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n539), .A2(KEYINPUT18), .A3(new_n540), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G197gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT11), .ZN(new_n551));
  INV_X1    g350(.A(G169gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT12), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n548), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n543), .A2(new_n554), .A3(new_n546), .A4(new_n547), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n556), .A2(KEYINPUT96), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT96), .B1(new_n556), .B2(new_n557), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n459), .A2(KEYINPUT35), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(new_n453), .A3(new_n441), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n457), .A2(new_n458), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n401), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n496), .A2(new_n494), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n448), .B(new_n478), .C1(new_n566), .C2(new_n483), .ZN(new_n567));
  INV_X1    g366(.A(new_n505), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(new_n569), .A3(KEYINPUT91), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT100), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(KEYINPUT7), .ZN(new_n572));
  NAND2_X1  g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(G99gat), .A2(G106gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n572), .A2(new_n573), .B1(KEYINPUT8), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(KEYINPUT7), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT100), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n576), .A2(new_n578), .A3(G85gat), .A4(G92gat), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n575), .B(new_n579), .C1(G85gat), .C2(G92gat), .ZN(new_n580));
  XOR2_X1   g379(.A(G99gat), .B(G106gat), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT101), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n580), .A2(new_n581), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n535), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n534), .ZN(new_n588));
  NAND3_X1  g387(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(G190gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(G218gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT102), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT99), .B(G134gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G162gat), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OR3_X1    g399(.A1(new_n594), .A2(new_n595), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n595), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G57gat), .B(G64gat), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G71gat), .B(G78gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT97), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT98), .B(KEYINPUT21), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI211_X1 g410(.A(new_n611), .B(new_n537), .C1(KEYINPUT21), .C2(new_n609), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n537), .A2(new_n611), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n615));
  XNOR2_X1  g414(.A(G155gat), .B(G183gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n614), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(new_n219), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G211gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n603), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT103), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n580), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n581), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n608), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(new_n587), .B2(new_n609), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n632), .A2(KEYINPUT10), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n609), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(G230gat), .ZN(new_n636));
  INV_X1    g435(.A(G233gat), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n632), .A2(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G176gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G204gat), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(KEYINPUT104), .A3(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n627), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n507), .A2(new_n561), .A3(new_n570), .A4(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n290), .B(KEYINPUT105), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g459(.A1(new_n476), .A2(new_n477), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(G8gat), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n656), .B(new_n662), .C1(new_n509), .C2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n509), .B2(new_n663), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n656), .B2(new_n662), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT42), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(KEYINPUT42), .B2(new_n665), .ZN(G1325gat));
  INV_X1    g467(.A(G15gat), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n655), .A2(new_n669), .A3(new_n568), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n449), .A2(new_n451), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n670), .B1(new_n673), .B2(new_n669), .ZN(G1326gat));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n563), .A2(KEYINPUT91), .A3(new_n569), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT91), .B1(new_n563), .B2(new_n569), .ZN(new_n677));
  INV_X1    g476(.A(new_n627), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n652), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n680), .A2(KEYINPUT106), .A3(new_n561), .A4(new_n401), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n655), .B2(new_n448), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n675), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n683), .A3(new_n675), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n685), .A2(G22gat), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(G22gat), .B1(new_n685), .B2(new_n686), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(G1327gat));
  NOR3_X1   g488(.A1(new_n676), .A2(new_n677), .A3(new_n603), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n653), .A2(new_n560), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n690), .A2(new_n625), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n519), .A3(new_n658), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n695), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n603), .A2(KEYINPUT44), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n563), .A2(KEYINPUT110), .A3(new_n569), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT110), .B1(new_n563), .B2(new_n569), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n690), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n625), .B(KEYINPUT108), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n556), .A2(new_n557), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(new_n706), .A3(new_n652), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT109), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n704), .A2(new_n657), .A3(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n696), .B(new_n697), .C1(new_n709), .C2(new_n519), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n690), .A2(new_n625), .A3(new_n691), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n711), .A2(G36gat), .A3(new_n661), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n704), .A2(new_n661), .A3(new_n708), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n714), .B(new_n715), .C1(new_n716), .C2(new_n520), .ZN(G1329gat));
  AND2_X1   g516(.A1(new_n601), .A2(new_n602), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n507), .A2(new_n570), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT44), .ZN(new_n720));
  AOI211_X1 g519(.A(new_n568), .B(new_n708), .C1(new_n720), .C2(new_n701), .ZN(new_n721));
  INV_X1    g520(.A(G43gat), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT111), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n692), .A2(new_n722), .A3(new_n672), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n721), .B2(new_n722), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI221_X1 g526(.A(new_n724), .B1(KEYINPUT111), .B2(KEYINPUT47), .C1(new_n721), .C2(new_n722), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1330gat));
  INV_X1    g528(.A(new_n708), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n703), .A2(G50gat), .A3(new_n401), .A4(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n711), .A2(new_n448), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(G50gat), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT48), .ZN(G1331gat));
  OR2_X1    g533(.A1(new_n699), .A2(new_n700), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n652), .A2(new_n706), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n678), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n658), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  INV_X1    g539(.A(KEYINPUT49), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n661), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT112), .ZN(new_n743));
  OR3_X1    g542(.A1(new_n737), .A2(KEYINPUT113), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT113), .B1(new_n737), .B2(new_n743), .ZN(new_n745));
  AND4_X1   g544(.A1(new_n741), .A2(new_n744), .A3(new_n364), .A4(new_n745), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n744), .A2(new_n745), .B1(new_n741), .B2(new_n364), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(G1333gat));
  OAI21_X1  g547(.A(G71gat), .B1(new_n737), .B2(new_n568), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n671), .A2(G71gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n737), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1334gat));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n401), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G78gat), .ZN(G1335gat));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n441), .A2(new_n453), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n505), .B1(new_n564), .B2(new_n401), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n757), .A2(new_n562), .B1(new_n758), .B2(new_n567), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n756), .B1(new_n759), .B2(new_n603), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n626), .A2(new_n706), .ZN(new_n761));
  OAI211_X1 g560(.A(KEYINPUT114), .B(new_n718), .C1(new_n460), .C2(new_n506), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n760), .A2(new_n762), .A3(KEYINPUT51), .A4(new_n761), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n767), .A2(new_n280), .A3(new_n658), .A4(new_n653), .ZN(new_n768));
  AND4_X1   g567(.A1(new_n658), .A2(new_n703), .A3(new_n653), .A4(new_n761), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n280), .ZN(G1336gat));
  NAND4_X1  g569(.A1(new_n703), .A2(new_n662), .A3(new_n653), .A4(new_n761), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G92gat), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n765), .A2(new_n773), .A3(new_n766), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n763), .A2(KEYINPUT115), .A3(new_n764), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n653), .A2(new_n662), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(G92gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT52), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(new_n767), .B2(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n772), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1337gat));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n413), .A3(new_n672), .A4(new_n653), .ZN(new_n784));
  AND4_X1   g583(.A1(new_n505), .A2(new_n703), .A3(new_n653), .A4(new_n761), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(new_n413), .ZN(G1338gat));
  NAND4_X1  g585(.A1(new_n703), .A2(new_n401), .A3(new_n653), .A4(new_n761), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G106gat), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n652), .A2(G106gat), .A3(new_n448), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n775), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT53), .B1(new_n767), .B2(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1339gat));
  NOR2_X1   g594(.A1(new_n539), .A2(new_n540), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n544), .A2(new_n545), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n553), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n800), .A2(new_n557), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n650), .A2(new_n802), .A3(new_n651), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT54), .B1(new_n635), .B2(new_n639), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n638), .B1(new_n633), .B2(new_n634), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n645), .B1(new_n640), .B2(KEYINPUT54), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n808), .A2(KEYINPUT116), .A3(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n642), .A2(new_n645), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n806), .A2(new_n807), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n816), .B2(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n706), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n803), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n603), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n601), .A2(new_n602), .A3(new_n817), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n812), .A2(new_n802), .A3(new_n813), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n705), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n627), .A2(new_n706), .A3(new_n653), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n657), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(new_n661), .A3(new_n440), .ZN(new_n828));
  OAI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n560), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n706), .A2(new_n226), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n828), .B2(new_n830), .ZN(G1340gat));
  NOR2_X1   g630(.A1(new_n828), .A2(new_n652), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(new_n224), .ZN(G1341gat));
  NOR3_X1   g632(.A1(new_n828), .A2(new_n219), .A3(new_n705), .ZN(new_n834));
  INV_X1    g633(.A(new_n828), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n626), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n834), .B1(new_n219), .B2(new_n836), .ZN(G1342gat));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n835), .A2(new_n838), .A3(new_n221), .A4(new_n718), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n835), .A2(new_n718), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT56), .B1(new_n841), .B2(G134gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(G134gat), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n840), .A2(new_n842), .A3(new_n843), .A4(new_n844), .ZN(G1343gat));
  OAI211_X1 g644(.A(new_n810), .B(new_n817), .C1(new_n558), .C2(new_n559), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n846), .A2(new_n803), .A3(KEYINPUT119), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT119), .B1(new_n846), .B2(new_n803), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n603), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT120), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n821), .A2(new_n822), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n852), .B(new_n603), .C1(new_n847), .C2(new_n848), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n825), .B1(new_n854), .B2(new_n625), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n448), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n824), .A2(new_n826), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n858), .A3(new_n401), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n505), .A2(new_n662), .A3(new_n657), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n856), .A2(new_n561), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(G141gat), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n661), .B1(new_n827), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n819), .A2(new_n603), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n851), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n825), .B1(new_n866), .B2(new_n705), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n867), .A2(KEYINPUT121), .A3(new_n657), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n505), .A2(new_n448), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n864), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n560), .A2(G141gat), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT122), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n862), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n856), .A2(new_n706), .A3(new_n859), .A4(new_n860), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n879), .A2(G141gat), .B1(new_n871), .B2(new_n874), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n877), .B1(new_n878), .B2(new_n880), .ZN(G1344gat));
  NAND3_X1  g680(.A1(new_n871), .A2(new_n206), .A3(new_n653), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n856), .A2(new_n653), .A3(new_n859), .A4(new_n860), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n883), .A2(new_n884), .A3(G148gat), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT57), .B1(new_n867), .B2(new_n448), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n679), .A2(new_n561), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n626), .B1(new_n851), .B2(new_n849), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n858), .B(new_n401), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n886), .A2(new_n889), .A3(new_n653), .A4(new_n860), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n884), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n882), .B1(new_n885), .B2(new_n891), .ZN(G1345gat));
  AOI21_X1  g691(.A(G155gat), .B1(new_n871), .B2(new_n626), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n856), .A2(new_n859), .A3(new_n860), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n705), .A2(new_n209), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(G1346gat));
  AOI21_X1  g695(.A(G162gat), .B1(new_n871), .B2(new_n718), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n603), .A2(new_n210), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n894), .B2(new_n898), .ZN(G1347gat));
  NAND2_X1  g698(.A1(new_n857), .A2(new_n657), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n452), .A2(new_n661), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT124), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n308), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n706), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906));
  INV_X1    g705(.A(new_n901), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n900), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n857), .A2(KEYINPUT125), .A3(new_n657), .A4(new_n901), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(new_n561), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n905), .B1(new_n911), .B2(new_n552), .ZN(G1348gat));
  AOI21_X1  g711(.A(G176gat), .B1(new_n903), .B2(new_n653), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n652), .A2(new_n299), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n910), .B2(new_n914), .ZN(G1349gat));
  INV_X1    g714(.A(new_n705), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n908), .A2(new_n916), .A3(new_n909), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G183gat), .ZN(new_n918));
  INV_X1    g717(.A(new_n327), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n919), .A3(new_n626), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT60), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n918), .A2(new_n923), .A3(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1350gat));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n718), .A3(new_n909), .ZN(new_n926));
  NAND2_X1  g725(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(G190gat), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n929), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n926), .A2(G190gat), .A3(new_n927), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n903), .A2(new_n718), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n930), .B(new_n932), .C1(G190gat), .C2(new_n933), .ZN(G1351gat));
  NOR2_X1   g733(.A1(new_n658), .A2(new_n505), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n662), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n886), .A2(new_n889), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n560), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n867), .A2(new_n448), .A3(new_n936), .ZN(new_n940));
  INV_X1    g739(.A(G197gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(new_n941), .A3(new_n706), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n939), .A2(new_n942), .ZN(G1352gat));
  XNOR2_X1  g742(.A(KEYINPUT127), .B(G204gat), .ZN(new_n944));
  NOR4_X1   g743(.A1(new_n900), .A2(new_n776), .A3(new_n870), .A4(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT62), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n886), .A2(new_n889), .A3(new_n653), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n947), .B2(new_n936), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1353gat));
  NAND3_X1  g748(.A1(new_n940), .A2(new_n339), .A3(new_n626), .ZN(new_n950));
  INV_X1    g749(.A(new_n938), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n626), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n952), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(G1354gat));
  AOI21_X1  g754(.A(G218gat), .B1(new_n940), .B2(new_n718), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n603), .A2(new_n340), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n951), .B2(new_n957), .ZN(G1355gat));
endmodule


