

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783;

  NAND2_X1 U373 ( .A1(n390), .A2(n388), .ZN(n644) );
  BUF_X1 U374 ( .A(n561), .Z(n350) );
  NAND2_X1 U375 ( .A1(n447), .A2(n445), .ZN(n621) );
  XNOR2_X1 U376 ( .A(n536), .B(n481), .ZN(n773) );
  XNOR2_X1 U377 ( .A(G119), .B(G128), .ZN(n493) );
  XNOR2_X1 U378 ( .A(G137), .B(KEYINPUT69), .ZN(n375) );
  BUF_X1 U379 ( .A(n516), .Z(n597) );
  BUF_X1 U380 ( .A(n584), .Z(n638) );
  XNOR2_X1 U381 ( .A(n516), .B(n485), .ZN(n553) );
  XNOR2_X2 U382 ( .A(n513), .B(KEYINPUT101), .ZN(n431) );
  XNOR2_X2 U383 ( .A(n555), .B(KEYINPUT33), .ZN(n728) );
  XNOR2_X2 U384 ( .A(n542), .B(KEYINPUT106), .ZN(n643) );
  AND2_X1 U385 ( .A1(n427), .A2(KEYINPUT107), .ZN(n425) );
  NOR2_X1 U386 ( .A1(n742), .A2(n741), .ZN(n745) );
  XNOR2_X1 U387 ( .A(n393), .B(n588), .ZN(n664) );
  AND2_X1 U388 ( .A1(n372), .A2(n424), .ZN(n371) );
  NAND2_X1 U389 ( .A1(n370), .A2(n425), .ZN(n369) );
  AND2_X1 U390 ( .A1(n552), .A2(n408), .ZN(n407) );
  XNOR2_X1 U391 ( .A(n405), .B(KEYINPUT42), .ZN(n668) );
  NOR2_X1 U392 ( .A1(n718), .A2(n431), .ZN(n430) );
  AND2_X1 U393 ( .A1(n695), .A2(n602), .ZN(n725) );
  XNOR2_X1 U394 ( .A(n638), .B(n585), .ZN(n721) );
  XNOR2_X1 U395 ( .A(n541), .B(n540), .ZN(n545) );
  XNOR2_X1 U396 ( .A(n529), .B(n528), .ZN(n559) );
  XNOR2_X1 U397 ( .A(n433), .B(n432), .ZN(n755) );
  XNOR2_X1 U398 ( .A(n479), .B(n478), .ZN(n536) );
  XNOR2_X1 U399 ( .A(n453), .B(G125), .ZN(n491) );
  XNOR2_X1 U400 ( .A(G143), .B(KEYINPUT102), .ZN(n521) );
  INV_X2 U401 ( .A(G953), .ZN(n465) );
  AND2_X2 U402 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U403 ( .A(n444), .B(n356), .ZN(n613) );
  AND2_X2 U404 ( .A1(n736), .A2(n743), .ZN(n354) );
  XNOR2_X2 U405 ( .A(n764), .B(KEYINPUT72), .ZN(n477) );
  XNOR2_X2 U406 ( .A(n441), .B(n458), .ZN(n764) );
  XNOR2_X2 U407 ( .A(n773), .B(G146), .ZN(n508) );
  XNOR2_X2 U408 ( .A(n579), .B(n380), .ZN(n561) );
  OR2_X2 U409 ( .A1(n683), .A2(n460), .ZN(n428) );
  OR2_X1 U410 ( .A1(n556), .A2(n547), .ZN(n549) );
  XNOR2_X1 U411 ( .A(G902), .B(KEYINPUT94), .ZN(n459) );
  XNOR2_X1 U412 ( .A(n385), .B(n384), .ZN(n525) );
  INV_X1 U413 ( .A(KEYINPUT78), .ZN(n384) );
  NAND2_X1 U414 ( .A1(n387), .A2(n386), .ZN(n385) );
  NAND2_X1 U415 ( .A1(n621), .A2(KEYINPUT39), .ZN(n392) );
  XNOR2_X1 U416 ( .A(n491), .B(n490), .ZN(n771) );
  XNOR2_X1 U417 ( .A(n725), .B(KEYINPUT86), .ZN(n608) );
  NOR2_X1 U418 ( .A1(n359), .A2(n395), .ZN(n394) );
  INV_X1 U419 ( .A(KEYINPUT44), .ZN(n395) );
  XNOR2_X1 U420 ( .A(G101), .B(KEYINPUT5), .ZN(n502) );
  INV_X1 U421 ( .A(KEYINPUT4), .ZN(n480) );
  XNOR2_X1 U422 ( .A(n496), .B(n436), .ZN(n530) );
  INV_X1 U423 ( .A(KEYINPUT8), .ZN(n436) );
  NAND2_X1 U424 ( .A1(n409), .A2(n414), .ZN(n415) );
  NAND2_X1 U425 ( .A1(n440), .A2(n739), .ZN(n411) );
  INV_X1 U426 ( .A(G902), .ZN(n539) );
  XNOR2_X1 U427 ( .A(n419), .B(n417), .ZN(n416) );
  INV_X1 U428 ( .A(G146), .ZN(n453) );
  XNOR2_X1 U429 ( .A(n383), .B(KEYINPUT41), .ZN(n748) );
  NOR2_X1 U430 ( .A1(n721), .A2(n381), .ZN(n383) );
  NOR2_X1 U431 ( .A1(n723), .A2(n720), .ZN(n382) );
  AND2_X1 U432 ( .A1(n392), .A2(n391), .ZN(n390) );
  NOR2_X1 U433 ( .A1(n755), .A2(G902), .ZN(n497) );
  XNOR2_X1 U434 ( .A(n544), .B(n543), .ZN(n602) );
  NAND2_X1 U435 ( .A1(n608), .A2(n426), .ZN(n424) );
  NOR2_X2 U436 ( .A1(n608), .A2(KEYINPUT47), .ZN(n422) );
  NAND2_X1 U437 ( .A1(n406), .A2(KEYINPUT91), .ZN(n400) );
  NOR2_X1 U438 ( .A1(n710), .A2(n377), .ZN(n711) );
  XNOR2_X1 U439 ( .A(n486), .B(KEYINPUT20), .ZN(n499) );
  XOR2_X1 U440 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n522) );
  INV_X1 U441 ( .A(n771), .ZN(n421) );
  XNOR2_X1 U442 ( .A(n418), .B(n526), .ZN(n417) );
  XNOR2_X1 U443 ( .A(G113), .B(G104), .ZN(n526) );
  XNOR2_X1 U444 ( .A(n527), .B(n520), .ZN(n418) );
  INV_X1 U445 ( .A(G122), .ZN(n527) );
  XOR2_X1 U446 ( .A(G140), .B(KEYINPUT82), .Z(n474) );
  OR2_X1 U447 ( .A1(n721), .A2(n720), .ZN(n724) );
  XNOR2_X1 U448 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n577) );
  XNOR2_X1 U449 ( .A(n592), .B(n591), .ZN(n367) );
  NAND2_X1 U450 ( .A1(n721), .A2(KEYINPUT39), .ZN(n391) );
  NOR2_X1 U451 ( .A1(n582), .A2(n579), .ZN(n512) );
  XNOR2_X1 U452 ( .A(n364), .B(KEYINPUT30), .ZN(n447) );
  XNOR2_X1 U453 ( .A(n508), .B(n507), .ZN(n669) );
  BUF_X1 U454 ( .A(n736), .Z(n737) );
  XNOR2_X1 U455 ( .A(n351), .B(G101), .ZN(n441) );
  XOR2_X1 U456 ( .A(G110), .B(KEYINPUT95), .Z(n351) );
  XOR2_X1 U457 ( .A(KEYINPUT104), .B(G107), .Z(n534) );
  XNOR2_X1 U458 ( .A(G116), .B(G122), .ZN(n533) );
  INV_X1 U459 ( .A(G134), .ZN(n478) );
  NAND2_X1 U460 ( .A1(n415), .A2(n411), .ZN(n410) );
  XNOR2_X1 U461 ( .A(n505), .B(n457), .ZN(n763) );
  XNOR2_X1 U462 ( .A(KEYINPUT16), .B(G122), .ZN(n457) );
  NAND2_X1 U463 ( .A1(G234), .A2(G237), .ZN(n464) );
  NOR2_X2 U464 ( .A1(n584), .A2(n720), .ZN(n444) );
  INV_X1 U465 ( .A(n621), .ZN(n624) );
  INV_X1 U466 ( .A(KEYINPUT6), .ZN(n380) );
  XNOR2_X1 U467 ( .A(n669), .B(KEYINPUT62), .ZN(n670) );
  XNOR2_X1 U468 ( .A(n495), .B(n771), .ZN(n432) );
  XNOR2_X1 U469 ( .A(n676), .B(n675), .ZN(n677) );
  AND2_X1 U470 ( .A1(n656), .A2(G953), .ZN(n758) );
  NOR2_X1 U471 ( .A1(n748), .A2(n611), .ZN(n405) );
  NAND2_X1 U472 ( .A1(n644), .A2(n586), .ZN(n393) );
  XNOR2_X1 U473 ( .A(n602), .B(n601), .ZN(n704) );
  OR2_X1 U474 ( .A1(n747), .A2(n352), .ZN(n404) );
  XNOR2_X1 U475 ( .A(n552), .B(n368), .ZN(n688) );
  INV_X1 U476 ( .A(G101), .ZN(n368) );
  XNOR2_X1 U477 ( .A(n459), .B(KEYINPUT15), .ZN(n650) );
  INV_X1 U478 ( .A(n608), .ZN(n427) );
  XOR2_X1 U479 ( .A(n749), .B(KEYINPUT119), .Z(n352) );
  XNOR2_X1 U480 ( .A(n497), .B(n498), .ZN(n713) );
  XOR2_X1 U481 ( .A(n634), .B(n603), .Z(n353) );
  AND2_X1 U482 ( .A1(n379), .A2(n367), .ZN(n355) );
  INV_X1 U483 ( .A(KEYINPUT107), .ZN(n426) );
  XOR2_X1 U484 ( .A(n463), .B(KEYINPUT19), .Z(n356) );
  XNOR2_X1 U485 ( .A(KEYINPUT84), .B(KEYINPUT34), .ZN(n357) );
  XOR2_X1 U486 ( .A(n652), .B(n654), .Z(n358) );
  AND2_X1 U487 ( .A1(KEYINPUT44), .A2(KEYINPUT91), .ZN(n359) );
  AND2_X1 U488 ( .A1(n460), .A2(KEYINPUT88), .ZN(n360) );
  INV_X1 U489 ( .A(G953), .ZN(n386) );
  AND2_X1 U490 ( .A1(n361), .A2(n386), .ZN(n750) );
  NOR2_X1 U491 ( .A1(n746), .A2(n404), .ZN(n361) );
  AND2_X1 U492 ( .A1(n437), .A2(n651), .ZN(n362) );
  NAND2_X1 U493 ( .A1(n736), .A2(n743), .ZN(n363) );
  AND2_X2 U494 ( .A1(n437), .A2(n651), .ZN(n754) );
  NAND2_X1 U495 ( .A1(n624), .A2(n389), .ZN(n388) );
  NOR2_X1 U496 ( .A1(n579), .A2(n720), .ZN(n364) );
  XNOR2_X1 U497 ( .A(n365), .B(KEYINPUT46), .ZN(n607) );
  NAND2_X1 U498 ( .A1(n600), .A2(n403), .ZN(n365) );
  XNOR2_X1 U499 ( .A(n434), .B(n435), .ZN(n433) );
  INV_X1 U500 ( .A(n713), .ZN(n378) );
  NAND2_X1 U501 ( .A1(n399), .A2(n569), .ZN(n571) );
  XNOR2_X1 U502 ( .A(n515), .B(KEYINPUT31), .ZN(n702) );
  XNOR2_X1 U503 ( .A(n366), .B(n492), .ZN(n434) );
  XNOR2_X1 U504 ( .A(n375), .B(KEYINPUT24), .ZN(n366) );
  NAND2_X1 U505 ( .A1(n367), .A2(n565), .ZN(n595) );
  NAND2_X1 U506 ( .A1(n423), .A2(n551), .ZN(n552) );
  NAND2_X1 U507 ( .A1(n371), .A2(n369), .ZN(n376) );
  OR2_X1 U508 ( .A1(n689), .A2(n702), .ZN(n370) );
  NAND2_X1 U509 ( .A1(n374), .A2(n373), .ZN(n372) );
  INV_X1 U510 ( .A(n702), .ZN(n373) );
  NOR2_X1 U511 ( .A1(n689), .A2(KEYINPUT107), .ZN(n374) );
  XNOR2_X1 U512 ( .A(n375), .B(KEYINPUT96), .ZN(n770) );
  NAND2_X1 U513 ( .A1(n376), .A2(n552), .ZN(n406) );
  NAND2_X1 U514 ( .A1(n376), .A2(n407), .ZN(n398) );
  INV_X1 U515 ( .A(n582), .ZN(n377) );
  NOR2_X1 U516 ( .A1(n561), .A2(n582), .ZN(n554) );
  NAND2_X1 U517 ( .A1(n350), .A2(n378), .ZN(n550) );
  INV_X1 U518 ( .A(n561), .ZN(n379) );
  INV_X1 U519 ( .A(n382), .ZN(n381) );
  NAND2_X1 U520 ( .A1(n525), .A2(G210), .ZN(n503) );
  INV_X1 U521 ( .A(G237), .ZN(n387) );
  NOR2_X1 U522 ( .A1(n721), .A2(KEYINPUT39), .ZN(n389) );
  NAND2_X1 U523 ( .A1(n665), .A2(n359), .ZN(n402) );
  NAND2_X1 U524 ( .A1(n665), .A2(n394), .ZN(n396) );
  NAND2_X1 U525 ( .A1(n397), .A2(n396), .ZN(n401) );
  NAND2_X1 U526 ( .A1(n398), .A2(n402), .ZN(n397) );
  NAND2_X1 U527 ( .A1(n401), .A2(n400), .ZN(n399) );
  NAND2_X1 U528 ( .A1(n530), .A2(G221), .ZN(n435) );
  NAND2_X1 U529 ( .A1(n613), .A2(n470), .ZN(n472) );
  INV_X1 U530 ( .A(n668), .ZN(n403) );
  INV_X1 U531 ( .A(KEYINPUT91), .ZN(n408) );
  NAND2_X1 U532 ( .A1(n743), .A2(n360), .ZN(n409) );
  NAND2_X1 U533 ( .A1(n412), .A2(n410), .ZN(n437) );
  NAND2_X1 U534 ( .A1(n413), .A2(n649), .ZN(n412) );
  NAND2_X1 U535 ( .A1(n354), .A2(n460), .ZN(n413) );
  NAND2_X1 U536 ( .A1(n460), .A2(KEYINPUT2), .ZN(n414) );
  XNOR2_X1 U537 ( .A(n420), .B(n416), .ZN(n676) );
  NAND2_X1 U538 ( .A1(n525), .A2(G214), .ZN(n419) );
  XNOR2_X1 U539 ( .A(n524), .B(n421), .ZN(n420) );
  INV_X1 U540 ( .A(n610), .ZN(n618) );
  XNOR2_X2 U541 ( .A(n422), .B(KEYINPUT76), .ZN(n610) );
  NAND2_X1 U542 ( .A1(n423), .A2(n566), .ZN(n567) );
  NAND2_X1 U543 ( .A1(n423), .A2(n563), .ZN(n564) );
  XNOR2_X2 U544 ( .A(n549), .B(n548), .ZN(n423) );
  XNOR2_X1 U545 ( .A(n519), .B(KEYINPUT100), .ZN(n689) );
  XNOR2_X2 U546 ( .A(n428), .B(n461), .ZN(n584) );
  XNOR2_X1 U547 ( .A(n429), .B(n477), .ZN(n683) );
  XNOR2_X1 U548 ( .A(n442), .B(n763), .ZN(n429) );
  NAND2_X1 U549 ( .A1(n514), .A2(n431), .ZN(n515) );
  XNOR2_X2 U550 ( .A(G143), .B(G128), .ZN(n479) );
  XNOR2_X2 U551 ( .A(n438), .B(KEYINPUT35), .ZN(n665) );
  NAND2_X1 U552 ( .A1(n439), .A2(n560), .ZN(n438) );
  XNOR2_X1 U553 ( .A(n557), .B(n357), .ZN(n439) );
  INV_X1 U554 ( .A(n736), .ZN(n440) );
  XNOR2_X1 U555 ( .A(n443), .B(n454), .ZN(n442) );
  XNOR2_X1 U556 ( .A(n452), .B(n451), .ZN(n443) );
  XNOR2_X1 U557 ( .A(n456), .B(n455), .ZN(n505) );
  NAND2_X1 U558 ( .A1(n353), .A2(n444), .ZN(n605) );
  AND2_X1 U559 ( .A1(n583), .A2(n597), .ZN(n445) );
  XOR2_X1 U560 ( .A(n712), .B(n501), .Z(n446) );
  NOR2_X1 U561 ( .A1(n607), .A2(n707), .ZN(n631) );
  INV_X1 U562 ( .A(KEYINPUT48), .ZN(n632) );
  INV_X1 U563 ( .A(n758), .ZN(n657) );
  AND2_X1 U564 ( .A1(n606), .A2(n710), .ZN(n707) );
  XNOR2_X2 U565 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n449) );
  XNOR2_X2 U566 ( .A(KEYINPUT18), .B(KEYINPUT83), .ZN(n448) );
  XNOR2_X1 U567 ( .A(n449), .B(n448), .ZN(n452) );
  NAND2_X1 U568 ( .A1(n465), .A2(G224), .ZN(n450) );
  XNOR2_X1 U569 ( .A(n450), .B(KEYINPUT4), .ZN(n451) );
  XNOR2_X1 U570 ( .A(n479), .B(n491), .ZN(n454) );
  XNOR2_X1 U571 ( .A(G116), .B(G113), .ZN(n456) );
  XNOR2_X1 U572 ( .A(KEYINPUT3), .B(G119), .ZN(n455) );
  XNOR2_X1 U573 ( .A(G104), .B(G107), .ZN(n458) );
  INV_X1 U574 ( .A(n650), .ZN(n460) );
  NAND2_X1 U575 ( .A1(n387), .A2(n539), .ZN(n462) );
  NAND2_X1 U576 ( .A1(n462), .A2(G210), .ZN(n461) );
  AND2_X1 U577 ( .A1(n462), .A2(G214), .ZN(n720) );
  INV_X1 U578 ( .A(KEYINPUT79), .ZN(n463) );
  XNOR2_X1 U579 ( .A(n464), .B(KEYINPUT14), .ZN(n709) );
  BUF_X2 U580 ( .A(n465), .Z(n774) );
  INV_X1 U581 ( .A(G952), .ZN(n656) );
  NAND2_X1 U582 ( .A1(n774), .A2(n656), .ZN(n467) );
  OR2_X1 U583 ( .A1(n774), .A2(G902), .ZN(n466) );
  AND2_X1 U584 ( .A1(n467), .A2(n466), .ZN(n468) );
  AND2_X1 U585 ( .A1(n709), .A2(n468), .ZN(n581) );
  NAND2_X1 U586 ( .A1(G953), .A2(G898), .ZN(n469) );
  AND2_X1 U587 ( .A1(n581), .A2(n469), .ZN(n470) );
  XNOR2_X1 U588 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n471) );
  XNOR2_X2 U589 ( .A(n472), .B(n471), .ZN(n556) );
  INV_X1 U590 ( .A(n556), .ZN(n514) );
  NAND2_X1 U591 ( .A1(G227), .A2(n774), .ZN(n473) );
  XNOR2_X1 U592 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U593 ( .A(n475), .B(n770), .ZN(n476) );
  XNOR2_X1 U594 ( .A(n477), .B(n476), .ZN(n482) );
  XNOR2_X1 U595 ( .A(n480), .B(G131), .ZN(n481) );
  XNOR2_X1 U596 ( .A(n508), .B(n482), .ZN(n652) );
  NAND2_X1 U597 ( .A1(n652), .A2(n539), .ZN(n484) );
  XOR2_X1 U598 ( .A(KEYINPUT71), .B(G469), .Z(n483) );
  XNOR2_X2 U599 ( .A(n484), .B(n483), .ZN(n516) );
  XNOR2_X1 U600 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n485) );
  XOR2_X1 U601 ( .A(KEYINPUT98), .B(KEYINPUT80), .Z(n488) );
  NAND2_X1 U602 ( .A1(G234), .A2(n650), .ZN(n486) );
  NAND2_X1 U603 ( .A1(n499), .A2(G217), .ZN(n487) );
  XNOR2_X1 U604 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U605 ( .A(n489), .B(KEYINPUT25), .ZN(n498) );
  XNOR2_X1 U606 ( .A(KEYINPUT10), .B(G140), .ZN(n490) );
  XOR2_X1 U607 ( .A(KEYINPUT81), .B(KEYINPUT97), .Z(n492) );
  XOR2_X1 U608 ( .A(KEYINPUT23), .B(G110), .Z(n494) );
  XNOR2_X1 U609 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U610 ( .A1(n774), .A2(G234), .ZN(n496) );
  NAND2_X1 U611 ( .A1(G221), .A2(n499), .ZN(n500) );
  XNOR2_X1 U612 ( .A(n500), .B(KEYINPUT21), .ZN(n712) );
  INV_X1 U613 ( .A(KEYINPUT99), .ZN(n501) );
  NAND2_X2 U614 ( .A1(n378), .A2(n446), .ZN(n582) );
  XNOR2_X1 U615 ( .A(n502), .B(G137), .ZN(n504) );
  XNOR2_X1 U616 ( .A(n504), .B(n503), .ZN(n506) );
  XNOR2_X1 U617 ( .A(n506), .B(n505), .ZN(n507) );
  OR2_X2 U618 ( .A1(n669), .A2(G902), .ZN(n511) );
  INV_X1 U619 ( .A(KEYINPUT74), .ZN(n509) );
  XNOR2_X1 U620 ( .A(n509), .B(G472), .ZN(n510) );
  XNOR2_X2 U621 ( .A(n511), .B(n510), .ZN(n579) );
  INV_X1 U622 ( .A(n579), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n553), .A2(n512), .ZN(n513) );
  NOR2_X1 U624 ( .A1(n582), .A2(n565), .ZN(n517) );
  NAND2_X1 U625 ( .A1(n517), .A2(n597), .ZN(n518) );
  NOR2_X1 U626 ( .A1(n556), .A2(n518), .ZN(n519) );
  INV_X1 U627 ( .A(KEYINPUT103), .ZN(n520) );
  XNOR2_X1 U628 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U629 ( .A(G131), .B(n523), .ZN(n524) );
  NAND2_X1 U630 ( .A1(n676), .A2(n539), .ZN(n529) );
  XOR2_X1 U631 ( .A(KEYINPUT13), .B(G475), .Z(n528) );
  XOR2_X1 U632 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n532) );
  NAND2_X1 U633 ( .A1(G217), .A2(n530), .ZN(n531) );
  XNOR2_X1 U634 ( .A(n532), .B(n531), .ZN(n538) );
  XNOR2_X1 U635 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U636 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U637 ( .A(n538), .B(n537), .ZN(n752) );
  NAND2_X1 U638 ( .A1(n752), .A2(n539), .ZN(n541) );
  INV_X1 U639 ( .A(G478), .ZN(n540) );
  NOR2_X1 U640 ( .A1(n559), .A2(n545), .ZN(n542) );
  INV_X1 U641 ( .A(n643), .ZN(n695) );
  NAND2_X1 U642 ( .A1(n559), .A2(n545), .ZN(n544) );
  INV_X1 U643 ( .A(KEYINPUT105), .ZN(n543) );
  INV_X1 U644 ( .A(n545), .ZN(n558) );
  OR2_X1 U645 ( .A1(n559), .A2(n558), .ZN(n723) );
  INV_X1 U646 ( .A(n723), .ZN(n546) );
  NAND2_X1 U647 ( .A1(n546), .A2(n446), .ZN(n547) );
  INV_X1 U648 ( .A(KEYINPUT22), .ZN(n548) );
  BUF_X1 U649 ( .A(n553), .Z(n710) );
  NOR2_X1 U650 ( .A1(n710), .A2(n550), .ZN(n551) );
  NOR2_X1 U651 ( .A1(n728), .A2(n556), .ZN(n557) );
  NAND2_X1 U652 ( .A1(n559), .A2(n558), .ZN(n622) );
  INV_X1 U653 ( .A(n622), .ZN(n560) );
  AND2_X1 U654 ( .A1(n350), .A2(n713), .ZN(n562) );
  AND2_X1 U655 ( .A1(n710), .A2(n562), .ZN(n563) );
  XNOR2_X1 U656 ( .A(n564), .B(KEYINPUT32), .ZN(n662) );
  NOR2_X1 U657 ( .A1(n710), .A2(n565), .ZN(n566) );
  XNOR2_X1 U658 ( .A(n567), .B(KEYINPUT65), .ZN(n568) );
  NAND2_X1 U659 ( .A1(n568), .A2(n713), .ZN(n666) );
  NAND2_X1 U660 ( .A1(n662), .A2(n666), .ZN(n572) );
  NAND2_X1 U661 ( .A1(n572), .A2(KEYINPUT44), .ZN(n569) );
  INV_X1 U662 ( .A(KEYINPUT90), .ZN(n570) );
  XNOR2_X1 U663 ( .A(n571), .B(n570), .ZN(n576) );
  OR2_X1 U664 ( .A1(n665), .A2(KEYINPUT44), .ZN(n573) );
  NOR2_X1 U665 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U666 ( .A(n574), .B(KEYINPUT73), .ZN(n575) );
  NAND2_X1 U667 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X2 U668 ( .A(n578), .B(n577), .ZN(n736) );
  NAND2_X1 U669 ( .A1(G953), .A2(G900), .ZN(n580) );
  NAND2_X1 U670 ( .A1(n581), .A2(n580), .ZN(n589) );
  NOR2_X1 U671 ( .A1(n582), .A2(n589), .ZN(n583) );
  XNOR2_X1 U672 ( .A(KEYINPUT77), .B(KEYINPUT38), .ZN(n585) );
  INV_X1 U673 ( .A(n602), .ZN(n586) );
  XNOR2_X1 U674 ( .A(KEYINPUT112), .B(KEYINPUT40), .ZN(n587) );
  XNOR2_X1 U675 ( .A(n587), .B(KEYINPUT111), .ZN(n588) );
  INV_X1 U676 ( .A(n664), .ZN(n600) );
  NOR2_X1 U677 ( .A1(n712), .A2(n589), .ZN(n590) );
  NAND2_X1 U678 ( .A1(n713), .A2(n590), .ZN(n592) );
  INV_X1 U679 ( .A(KEYINPUT70), .ZN(n591) );
  INV_X1 U680 ( .A(KEYINPUT110), .ZN(n593) );
  XNOR2_X1 U681 ( .A(n593), .B(KEYINPUT28), .ZN(n594) );
  XNOR2_X1 U682 ( .A(n595), .B(n594), .ZN(n599) );
  INV_X1 U683 ( .A(KEYINPUT109), .ZN(n596) );
  XNOR2_X1 U684 ( .A(n597), .B(n596), .ZN(n598) );
  NAND2_X1 U685 ( .A1(n599), .A2(n598), .ZN(n611) );
  INV_X1 U686 ( .A(KEYINPUT108), .ZN(n601) );
  NAND2_X1 U687 ( .A1(n704), .A2(n355), .ZN(n634) );
  INV_X1 U688 ( .A(KEYINPUT113), .ZN(n603) );
  INV_X1 U689 ( .A(KEYINPUT36), .ZN(n604) );
  XNOR2_X1 U690 ( .A(n605), .B(n604), .ZN(n606) );
  INV_X1 U691 ( .A(KEYINPUT75), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n610), .A2(n609), .ZN(n614) );
  INV_X1 U693 ( .A(n611), .ZN(n612) );
  AND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n700) );
  NAND2_X1 U695 ( .A1(n614), .A2(n700), .ZN(n617) );
  INV_X1 U696 ( .A(n700), .ZN(n696) );
  NOR2_X1 U697 ( .A1(KEYINPUT75), .A2(KEYINPUT47), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n696), .A2(n615), .ZN(n616) );
  NAND2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n629) );
  AND2_X1 U700 ( .A1(n618), .A2(KEYINPUT75), .ZN(n627) );
  NAND2_X1 U701 ( .A1(KEYINPUT47), .A2(n725), .ZN(n620) );
  INV_X1 U702 ( .A(KEYINPUT85), .ZN(n619) );
  XNOR2_X1 U703 ( .A(n620), .B(n619), .ZN(n625) );
  NOR2_X1 U704 ( .A1(n622), .A2(n638), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n660) );
  NAND2_X1 U706 ( .A1(n625), .A2(n660), .ZN(n626) );
  NOR2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n628) );
  AND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n633), .B(n632), .ZN(n641) );
  INV_X1 U711 ( .A(n634), .ZN(n636) );
  NOR2_X1 U712 ( .A1(n710), .A2(n720), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U714 ( .A(n637), .B(KEYINPUT43), .ZN(n639) );
  AND2_X1 U715 ( .A1(n638), .A2(n639), .ZN(n661) );
  INV_X1 U716 ( .A(n661), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n642), .B(KEYINPUT89), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n646) );
  INV_X1 U720 ( .A(KEYINPUT114), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(n783) );
  INV_X1 U722 ( .A(n783), .ZN(n647) );
  AND2_X2 U723 ( .A1(n648), .A2(n647), .ZN(n743) );
  INV_X1 U724 ( .A(KEYINPUT88), .ZN(n649) );
  INV_X1 U725 ( .A(KEYINPUT2), .ZN(n739) );
  OR2_X1 U726 ( .A1(n363), .A2(n739), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n362), .A2(G469), .ZN(n655) );
  XNOR2_X1 U728 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n653), .B(KEYINPUT58), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n655), .B(n358), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U733 ( .A(n660), .B(G143), .ZN(G45) );
  XOR2_X1 U734 ( .A(G140), .B(n661), .Z(G42) );
  XNOR2_X1 U735 ( .A(n662), .B(G119), .ZN(G21) );
  XNOR2_X1 U736 ( .A(G131), .B(KEYINPUT127), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(G33) );
  XOR2_X1 U738 ( .A(n665), .B(G122), .Z(G24) );
  XNOR2_X1 U739 ( .A(n666), .B(G110), .ZN(G12) );
  XOR2_X1 U740 ( .A(G137), .B(KEYINPUT126), .Z(n667) );
  XNOR2_X1 U741 ( .A(n668), .B(n667), .ZN(G39) );
  NAND2_X1 U742 ( .A1(n754), .A2(G472), .ZN(n671) );
  XNOR2_X1 U743 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X2 U744 ( .A1(n672), .A2(n758), .ZN(n674) );
  XNOR2_X1 U745 ( .A(KEYINPUT93), .B(KEYINPUT63), .ZN(n673) );
  XNOR2_X1 U746 ( .A(n674), .B(n673), .ZN(G57) );
  NAND2_X1 U747 ( .A1(n754), .A2(G475), .ZN(n678) );
  XOR2_X1 U748 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n675) );
  XNOR2_X1 U749 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X2 U750 ( .A1(n679), .A2(n758), .ZN(n681) );
  XNOR2_X1 U751 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n680) );
  XNOR2_X1 U752 ( .A(n681), .B(n680), .ZN(G60) );
  NAND2_X1 U753 ( .A1(n754), .A2(G210), .ZN(n685) );
  XOR2_X1 U754 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n682) );
  XNOR2_X1 U755 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U756 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X2 U757 ( .A1(n686), .A2(n758), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n687), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT115), .ZN(G3) );
  NAND2_X1 U760 ( .A1(n689), .A2(n704), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n690), .B(G104), .ZN(G6) );
  XNOR2_X1 U762 ( .A(G107), .B(KEYINPUT116), .ZN(n694) );
  XOR2_X1 U763 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n692) );
  NAND2_X1 U764 ( .A1(n689), .A2(n643), .ZN(n691) );
  XNOR2_X1 U765 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U766 ( .A(n694), .B(n693), .ZN(G9) );
  NOR2_X1 U767 ( .A1(n696), .A2(n695), .ZN(n698) );
  XNOR2_X1 U768 ( .A(KEYINPUT29), .B(KEYINPUT117), .ZN(n697) );
  XNOR2_X1 U769 ( .A(n698), .B(n697), .ZN(n699) );
  XOR2_X1 U770 ( .A(G128), .B(n699), .Z(G30) );
  NAND2_X1 U771 ( .A1(n700), .A2(n704), .ZN(n701) );
  XNOR2_X1 U772 ( .A(n701), .B(G146), .ZN(G48) );
  BUF_X1 U773 ( .A(n702), .Z(n703) );
  NAND2_X1 U774 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U775 ( .A(n705), .B(G113), .ZN(G15) );
  NAND2_X1 U776 ( .A1(n643), .A2(n703), .ZN(n706) );
  XNOR2_X1 U777 ( .A(n706), .B(G116), .ZN(G18) );
  XNOR2_X1 U778 ( .A(G125), .B(n707), .ZN(n708) );
  XNOR2_X1 U779 ( .A(n708), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U780 ( .A1(G952), .A2(n709), .ZN(n735) );
  XNOR2_X1 U781 ( .A(n711), .B(KEYINPUT50), .ZN(n717) );
  AND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U783 ( .A(n714), .B(KEYINPUT49), .ZN(n715) );
  NAND2_X1 U784 ( .A1(n715), .A2(n579), .ZN(n716) );
  NOR2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U786 ( .A(KEYINPUT51), .B(n430), .Z(n719) );
  OR2_X1 U787 ( .A1(n719), .A2(n748), .ZN(n731) );
  AND2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n727) );
  NOR2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U791 ( .A1(n727), .A2(n726), .ZN(n729) );
  OR2_X1 U792 ( .A1(n729), .A2(n728), .ZN(n730) );
  AND2_X1 U793 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U794 ( .A(KEYINPUT52), .B(n732), .ZN(n733) );
  XNOR2_X1 U795 ( .A(KEYINPUT118), .B(n733), .ZN(n734) );
  NOR2_X1 U796 ( .A1(n735), .A2(n734), .ZN(n747) );
  XNOR2_X1 U797 ( .A(n737), .B(KEYINPUT87), .ZN(n738) );
  NOR2_X1 U798 ( .A1(n738), .A2(KEYINPUT2), .ZN(n742) );
  NOR2_X1 U799 ( .A1(n739), .A2(KEYINPUT87), .ZN(n740) );
  AND2_X1 U800 ( .A1(n363), .A2(n740), .ZN(n741) );
  NOR2_X1 U801 ( .A1(n743), .A2(KEYINPUT2), .ZN(n744) );
  NOR2_X1 U802 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U803 ( .A1(n728), .A2(n748), .ZN(n749) );
  XNOR2_X1 U804 ( .A(n750), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U805 ( .A1(n362), .A2(G478), .ZN(n751) );
  XOR2_X1 U806 ( .A(n752), .B(n751), .Z(n753) );
  NOR2_X1 U807 ( .A1(n758), .A2(n753), .ZN(G63) );
  NAND2_X1 U808 ( .A1(n362), .A2(G217), .ZN(n756) );
  XNOR2_X1 U809 ( .A(n756), .B(n755), .ZN(n757) );
  NOR2_X1 U810 ( .A1(n758), .A2(n757), .ZN(G66) );
  NAND2_X1 U811 ( .A1(n737), .A2(n774), .ZN(n762) );
  NAND2_X1 U812 ( .A1(G953), .A2(G224), .ZN(n759) );
  XNOR2_X1 U813 ( .A(KEYINPUT61), .B(n759), .ZN(n760) );
  NAND2_X1 U814 ( .A1(n760), .A2(G898), .ZN(n761) );
  NAND2_X1 U815 ( .A1(n762), .A2(n761), .ZN(n768) );
  XNOR2_X1 U816 ( .A(n764), .B(n763), .ZN(n766) );
  NOR2_X1 U817 ( .A1(G898), .A2(n774), .ZN(n765) );
  NOR2_X1 U818 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U819 ( .A(n768), .B(n767), .ZN(n769) );
  XOR2_X1 U820 ( .A(KEYINPUT123), .B(n769), .Z(G69) );
  XNOR2_X1 U821 ( .A(n771), .B(n770), .ZN(n772) );
  XNOR2_X1 U822 ( .A(n773), .B(n772), .ZN(n776) );
  XNOR2_X1 U823 ( .A(n743), .B(n776), .ZN(n775) );
  NAND2_X1 U824 ( .A1(n775), .A2(n774), .ZN(n782) );
  XOR2_X1 U825 ( .A(KEYINPUT124), .B(n776), .Z(n777) );
  XNOR2_X1 U826 ( .A(G227), .B(n777), .ZN(n778) );
  NAND2_X1 U827 ( .A1(G900), .A2(n778), .ZN(n779) );
  NAND2_X1 U828 ( .A1(G953), .A2(n779), .ZN(n780) );
  XOR2_X1 U829 ( .A(KEYINPUT125), .B(n780), .Z(n781) );
  NAND2_X1 U830 ( .A1(n782), .A2(n781), .ZN(G72) );
  XOR2_X1 U831 ( .A(G134), .B(n783), .Z(G36) );
endmodule

