//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  AOI21_X1  g001(.A(new_n202), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR3_X1   g004(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207));
  OAI221_X1 g006(.A(new_n203), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(KEYINPUT15), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n208), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT84), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n208), .B(new_n209), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(KEYINPUT84), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT86), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(G1gat), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n217), .B(KEYINPUT86), .ZN(new_n223));
  INV_X1    g022(.A(G1gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n221), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n222), .B1(new_n221), .B2(new_n225), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT88), .B1(new_n216), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n211), .B(new_n212), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT88), .ZN(new_n232));
  INV_X1    g031(.A(new_n228), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n226), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT87), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n229), .A2(KEYINPUT87), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n213), .B2(new_n215), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n214), .A2(KEYINPUT17), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n239), .A2(new_n240), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n236), .A2(new_n237), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT18), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n216), .A2(new_n229), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n236), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n237), .B(KEYINPUT13), .Z(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n236), .A2(KEYINPUT18), .A3(new_n237), .A4(new_n244), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n247), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT82), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G197gat), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT11), .B(G169gat), .Z(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n258), .B(KEYINPUT12), .Z(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n259), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n253), .A2(KEYINPUT82), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT31), .B(G50gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g065(.A(KEYINPUT3), .ZN(new_n267));
  XNOR2_X1  g066(.A(G197gat), .B(G204gat), .ZN(new_n268));
  INV_X1    g067(.A(G211gat), .ZN(new_n269));
  INV_X1    g068(.A(G218gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n268), .B1(KEYINPUT22), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n273));
  XOR2_X1   g072(.A(G211gat), .B(G218gat), .Z(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n272), .B(new_n274), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(new_n273), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n267), .B1(new_n277), .B2(KEYINPUT29), .ZN(new_n278));
  INV_X1    g077(.A(G141gat), .ZN(new_n279));
  INV_X1    g078(.A(G148gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT68), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT2), .ZN(new_n285));
  NAND2_X1  g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n281), .A2(new_n283), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G155gat), .B(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  INV_X1    g095(.A(G162gat), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT2), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n294), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n291), .A2(KEYINPUT69), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT69), .B1(new_n291), .B2(new_n299), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n278), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n291), .A2(new_n299), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(KEYINPUT3), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n277), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G228gat), .ZN(new_n310));
  INV_X1    g109(.A(G233gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n277), .A2(KEYINPUT75), .A3(new_n306), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n303), .A2(new_n309), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n307), .ZN(new_n315));
  XNOR2_X1  g114(.A(G141gat), .B(G148gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n290), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n317), .A2(new_n298), .B1(new_n290), .B2(new_n287), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n276), .A2(new_n304), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(new_n267), .ZN(new_n320));
  OAI22_X1  g119(.A1(new_n315), .A2(new_n320), .B1(new_n310), .B2(new_n311), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n266), .B1(new_n322), .B2(G22gat), .ZN(new_n323));
  XOR2_X1   g122(.A(KEYINPUT76), .B(G22gat), .Z(new_n324));
  NAND4_X1  g123(.A1(new_n314), .A2(KEYINPUT77), .A3(new_n324), .A4(new_n321), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n314), .A2(new_n324), .A3(new_n321), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n323), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n326), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n324), .B1(new_n314), .B2(new_n321), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n266), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT65), .ZN(new_n337));
  NOR2_X1   g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT26), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT65), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n334), .A2(new_n341), .A3(new_n335), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n337), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G183gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT27), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT27), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G183gat), .ZN(new_n347));
  INV_X1    g146(.A(G190gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n349), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n345), .A2(new_n347), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n348), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n343), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT24), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(G183gat), .A3(G190gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G183gat), .B(G190gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(new_n355), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(G169gat), .B2(G176gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n338), .A2(KEYINPUT23), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT64), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n335), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n358), .A2(new_n361), .A3(new_n366), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n355), .A2(G183gat), .A3(G190gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n344), .A2(G190gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n348), .A2(G183gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n368), .B1(new_n371), .B2(KEYINPUT24), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n362), .A2(new_n335), .A3(new_n360), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT25), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n354), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G113gat), .B(G120gat), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT66), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT1), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G127gat), .B(G134gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n381), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n376), .B2(new_n379), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n375), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n362), .A2(new_n335), .A3(new_n360), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n358), .B2(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n366), .A2(new_n361), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n358), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n382), .A2(new_n384), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n354), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT33), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G15gat), .B(G43gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G71gat), .B(G99gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT34), .B1(new_n394), .B2(new_n396), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT34), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n386), .A2(new_n393), .A3(new_n403), .A4(new_n395), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n394), .A2(new_n396), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT32), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n402), .B(new_n404), .C1(new_n397), .C2(new_n400), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n406), .B2(new_n410), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n333), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n277), .ZN(new_n416));
  INV_X1    g215(.A(G226gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(new_n311), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n375), .B2(new_n304), .ZN(new_n419));
  INV_X1    g218(.A(new_n418), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n391), .B2(new_n354), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n416), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n375), .A2(new_n418), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT29), .B1(new_n391), .B2(new_n354), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n427), .B(new_n277), .C1(new_n428), .C2(new_n418), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n422), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT30), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n426), .B1(new_n422), .B2(new_n429), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI211_X1 g232(.A(KEYINPUT30), .B(new_n426), .C1(new_n422), .C2(new_n429), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G1gat), .B(G29gat), .Z(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G57gat), .B(G85gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n392), .A2(new_n318), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n444), .B(KEYINPUT72), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n392), .A2(KEYINPUT4), .A3(new_n318), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT71), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT70), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n318), .B2(new_n267), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n302), .B2(KEYINPUT3), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT69), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n294), .A2(new_n295), .A3(new_n298), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n295), .B1(new_n294), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n291), .A2(KEYINPUT69), .A3(new_n299), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n457), .A2(KEYINPUT70), .A3(KEYINPUT3), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n385), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n449), .B1(new_n452), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(KEYINPUT3), .A3(new_n458), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT70), .B1(new_n305), .B2(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n464), .A2(KEYINPUT71), .A3(new_n385), .A4(new_n459), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n448), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT73), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n457), .A2(new_n458), .A3(new_n385), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n441), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n469), .B2(new_n446), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n441), .A2(new_n468), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(KEYINPUT73), .A3(new_n445), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(KEYINPUT5), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  AOI211_X1 g273(.A(KEYINPUT5), .B(new_n448), .C1(new_n461), .C2(new_n465), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n440), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n466), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n440), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n478), .B(new_n479), .C1(new_n466), .C2(new_n473), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(KEYINPUT6), .B(new_n440), .C1(new_n474), .C2(new_n475), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n435), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n415), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT35), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n333), .A2(new_n414), .A3(KEYINPUT81), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n415), .B(new_n484), .C1(KEYINPUT81), .C2(KEYINPUT35), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT80), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT37), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n422), .A2(new_n493), .A3(new_n429), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n422), .B2(new_n429), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n426), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n496), .A2(KEYINPUT38), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n432), .B1(new_n496), .B2(KEYINPUT38), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n333), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n443), .A2(new_n447), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n460), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT71), .B1(new_n503), .B2(new_n464), .ZN(new_n504));
  AND4_X1   g303(.A1(KEYINPUT71), .A2(new_n464), .A3(new_n385), .A4(new_n459), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT39), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n507), .A3(new_n445), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n469), .B2(new_n446), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n501), .B1(new_n461), .B2(new_n465), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(new_n446), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n508), .A2(new_n511), .A3(KEYINPUT40), .A4(new_n479), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n435), .A2(new_n512), .A3(new_n476), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n508), .A2(new_n511), .A3(KEYINPUT78), .A4(new_n479), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT79), .B(KEYINPUT40), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n508), .A2(new_n511), .A3(new_n479), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT78), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n513), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n492), .B1(new_n500), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n517), .ZN(new_n521));
  INV_X1    g320(.A(new_n515), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n514), .A3(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n435), .A2(new_n512), .A3(new_n476), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n525), .A2(KEYINPUT80), .A3(new_n333), .A4(new_n499), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(new_n412), .B2(new_n413), .ZN(new_n529));
  INV_X1    g328(.A(new_n413), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(KEYINPUT36), .A3(new_n411), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(new_n484), .B2(new_n333), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n263), .B1(new_n491), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT8), .ZN(new_n537));
  NAND2_X1  g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(KEYINPUT96), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(KEYINPUT96), .B2(new_n538), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT97), .B(G85gat), .ZN(new_n541));
  INV_X1    g340(.A(G92gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G85gat), .A2(G92gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G99gat), .B(G106gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n242), .A2(new_n243), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT41), .ZN(new_n550));
  INV_X1    g349(.A(G232gat), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n550), .A2(new_n551), .A3(new_n311), .ZN(new_n552));
  INV_X1    g351(.A(new_n548), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n552), .B1(new_n231), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT98), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n549), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(new_n549), .B2(new_n554), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT95), .ZN(new_n560));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n550), .B1(new_n551), .B2(new_n311), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT99), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n559), .A2(KEYINPUT95), .A3(new_n566), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n568), .B(new_n569), .C1(KEYINPUT99), .C2(new_n559), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G57gat), .B(G64gat), .Z(new_n572));
  NAND2_X1  g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(G71gat), .A2(G78gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(KEYINPUT89), .A2(new_n575), .B1(new_n577), .B2(new_n573), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n234), .B1(KEYINPUT21), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n582), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G127gat), .B(G155gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT20), .ZN(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT90), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n588), .B(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G183gat), .B(G211gat), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT92), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n591), .B(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n586), .B(new_n594), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n571), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(G176gat), .B(G204gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n597), .B(new_n598), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT103), .ZN(new_n602));
  INV_X1    g401(.A(new_n547), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n546), .A2(KEYINPUT100), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT100), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n547), .B2(KEYINPUT101), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n546), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n581), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n548), .A2(new_n579), .A3(new_n580), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n553), .A2(KEYINPUT10), .A3(new_n581), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n602), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n602), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n616), .B1(new_n610), .B2(new_n612), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n600), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT104), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT104), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n620), .B(new_n600), .C1(new_n615), .C2(new_n617), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT102), .B1(new_n613), .B2(new_n614), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(new_n602), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n613), .A2(KEYINPUT102), .A3(new_n614), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n617), .A2(new_n600), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n619), .A2(new_n621), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n596), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n536), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n482), .A2(new_n483), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n224), .ZN(G1324gat));
  INV_X1    g432(.A(new_n435), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  AOI21_X1  g435(.A(KEYINPUT42), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  OAI21_X1  g437(.A(G8gat), .B1(new_n630), .B2(new_n634), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n640), .B2(KEYINPUT42), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT105), .Z(G1325gat));
  INV_X1    g441(.A(new_n630), .ZN(new_n643));
  AOI21_X1  g442(.A(G15gat), .B1(new_n643), .B2(new_n414), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n532), .B(KEYINPUT106), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(G15gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(KEYINPUT107), .Z(new_n647));
  AOI21_X1  g446(.A(new_n644), .B1(new_n643), .B2(new_n647), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n630), .A2(new_n333), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT43), .B(G22gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  INV_X1    g450(.A(new_n595), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n570), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n627), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT108), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n536), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n657), .A2(G29gat), .A3(new_n631), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT45), .Z(new_n659));
  NOR3_X1   g458(.A1(new_n263), .A2(new_n595), .A3(new_n628), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n571), .A2(KEYINPUT44), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n535), .A2(KEYINPUT109), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n533), .B1(new_n520), .B2(new_n526), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT109), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n662), .B1(new_n667), .B2(new_n491), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n570), .B1(new_n490), .B2(new_n664), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n669), .A2(KEYINPUT44), .ZN(new_n670));
  OAI211_X1 g469(.A(KEYINPUT110), .B(new_n660), .C1(new_n668), .C2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT110), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n665), .B1(new_n527), .B2(new_n534), .ZN(new_n673));
  AOI211_X1 g472(.A(KEYINPUT109), .B(new_n533), .C1(new_n520), .C2(new_n526), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n491), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n675), .A2(new_n661), .B1(KEYINPUT44), .B2(new_n669), .ZN(new_n676));
  INV_X1    g475(.A(new_n660), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n631), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n671), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(G29gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n659), .A2(new_n681), .ZN(G1328gat));
  NOR3_X1   g481(.A1(new_n657), .A2(G36gat), .A3(new_n634), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT46), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n671), .A2(new_n678), .A3(new_n435), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT111), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(G36gat), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n685), .A2(KEYINPUT111), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n684), .B1(new_n687), .B2(new_n688), .ZN(G1329gat));
  NOR4_X1   g488(.A1(new_n657), .A2(G43gat), .A3(new_n412), .A4(new_n413), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(G43gat), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n676), .A2(new_n532), .A3(new_n677), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n691), .B(KEYINPUT47), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n671), .A2(new_n678), .A3(new_n645), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n690), .B1(new_n695), .B2(G43gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n696), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g496(.A(new_n333), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n671), .A2(new_n678), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G50gat), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n333), .A2(G50gat), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n657), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT48), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n698), .B(new_n660), .C1(new_n668), .C2(new_n670), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G50gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n702), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT48), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n706), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n704), .B1(new_n699), .B2(G50gat), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n703), .B1(new_n709), .B2(new_n702), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT112), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(G1331gat));
  INV_X1    g515(.A(new_n675), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n263), .A2(new_n628), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n717), .A2(new_n596), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n679), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g520(.A(new_n435), .B(KEYINPUT113), .Z(new_n722));
  OR3_X1    g521(.A1(new_n717), .A2(new_n596), .A3(new_n718), .ZN(new_n723));
  AOI211_X1 g522(.A(new_n722), .B(new_n723), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1333gat));
  INV_X1    g525(.A(new_n645), .ZN(new_n727));
  OAI21_X1  g526(.A(G71gat), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(G71gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n719), .A2(new_n729), .A3(new_n414), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g531(.A1(new_n719), .A2(new_n698), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g533(.A1(new_n263), .A2(new_n652), .A3(new_n628), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n668), .B2(new_n670), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n631), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n654), .A2(new_n263), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT51), .B1(new_n717), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n675), .A2(new_n741), .A3(new_n263), .A4(new_n654), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n628), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n679), .A2(new_n541), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n738), .A2(new_n541), .B1(new_n743), .B2(new_n744), .ZN(G1336gat));
  OAI21_X1  g544(.A(G92gat), .B1(new_n737), .B2(new_n722), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n747));
  NOR2_X1   g546(.A1(new_n722), .A2(G92gat), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n746), .B(new_n747), .C1(new_n743), .C2(new_n749), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n676), .A2(new_n634), .A3(new_n735), .ZN(new_n751));
  OAI22_X1  g550(.A1(new_n743), .A2(new_n749), .B1(new_n751), .B2(new_n542), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n752), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT114), .B1(new_n752), .B2(KEYINPUT52), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(G1337gat));
  NAND2_X1  g554(.A1(new_n645), .A2(G99gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n737), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(G99gat), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n740), .A2(new_n414), .A3(new_n628), .A4(new_n742), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT116), .ZN(G1338gat));
  OAI211_X1 g560(.A(new_n698), .B(new_n736), .C1(new_n668), .C2(new_n670), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G106gat), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n333), .A2(G106gat), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n740), .A2(new_n628), .A3(new_n742), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n763), .A2(KEYINPUT118), .A3(new_n764), .A4(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n763), .A2(new_n766), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT117), .B1(new_n772), .B2(KEYINPUT53), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n772), .A2(KEYINPUT117), .A3(KEYINPUT53), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(G1339gat));
  NAND2_X1  g574(.A1(new_n629), .A2(new_n263), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n247), .A2(new_n251), .A3(new_n252), .A4(new_n261), .ZN(new_n777));
  INV_X1    g576(.A(new_n250), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n236), .A2(new_n248), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n237), .B1(new_n236), .B2(new_n244), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n258), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n599), .B1(new_n615), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n624), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n786), .A2(new_n602), .A3(new_n622), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n613), .A2(new_n614), .A3(new_n602), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT54), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT55), .B(new_n785), .C1(new_n787), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n625), .A2(new_n626), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n789), .B1(new_n623), .B2(new_n624), .ZN(new_n794));
  INV_X1    g593(.A(new_n785), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n570), .A2(new_n783), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n782), .B2(new_n627), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n628), .A2(KEYINPUT119), .A3(new_n781), .A4(new_n777), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n796), .A2(new_n790), .A3(new_n791), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n800), .B(new_n801), .C1(new_n263), .C2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n798), .B1(new_n803), .B2(new_n571), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n652), .B1(new_n804), .B2(KEYINPUT120), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n800), .A2(new_n801), .ZN(new_n806));
  INV_X1    g605(.A(new_n262), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n261), .B1(new_n253), .B2(KEYINPUT82), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n807), .A2(new_n802), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n571), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n797), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n776), .B1(new_n805), .B2(new_n813), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n814), .A2(new_n679), .A3(new_n415), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n815), .A2(new_n722), .ZN(new_n816));
  INV_X1    g615(.A(new_n263), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n628), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g620(.A1(new_n816), .A2(new_n595), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(G127gat), .ZN(G1342gat));
  INV_X1    g622(.A(G134gat), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n571), .A2(new_n435), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n815), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n816), .A2(new_n570), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n824), .ZN(G1343gat));
  NAND3_X1  g629(.A1(new_n722), .A2(new_n679), .A3(new_n532), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  INV_X1    g631(.A(new_n776), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n595), .B1(new_n811), .B2(new_n812), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n804), .A2(KEYINPUT120), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n836), .B2(new_n333), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n333), .A2(new_n832), .ZN(new_n838));
  OR3_X1    g637(.A1(new_n794), .A2(KEYINPUT121), .A3(new_n795), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT121), .B1(new_n794), .B2(new_n795), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n793), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n841), .A2(new_n260), .A3(new_n262), .A4(new_n792), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n783), .A2(new_n628), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n571), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n798), .B1(new_n845), .B2(KEYINPUT122), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n570), .B1(new_n842), .B2(new_n843), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n595), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n838), .B1(new_n850), .B2(new_n833), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n831), .B1(new_n837), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n279), .B1(new_n852), .B2(new_n817), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n836), .A2(new_n333), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n645), .A2(new_n631), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n722), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n817), .A2(new_n279), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT123), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT58), .B1(new_n853), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n831), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT57), .B1(new_n814), .B2(new_n698), .ZN(new_n863));
  INV_X1    g662(.A(new_n838), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n849), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n652), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n866), .B2(new_n776), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n862), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G141gat), .B1(new_n868), .B2(new_n263), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n856), .A2(new_n859), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n861), .A2(new_n872), .ZN(G1344gat));
  OAI21_X1  g672(.A(KEYINPUT59), .B1(new_n856), .B2(new_n627), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n280), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n862), .A2(new_n628), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(KEYINPUT59), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n863), .B2(new_n867), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n776), .A2(KEYINPUT124), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n652), .B1(new_n847), .B2(new_n798), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n776), .A2(KEYINPUT124), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(new_n882), .B2(new_n698), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n836), .A2(new_n864), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT59), .B(G148gat), .C1(new_n885), .C2(new_n876), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n875), .A2(new_n878), .A3(new_n886), .ZN(G1345gat));
  AOI21_X1  g686(.A(new_n296), .B1(new_n852), .B2(new_n595), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n652), .A2(G155gat), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n856), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT125), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G155gat), .B1(new_n868), .B2(new_n652), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n856), .A2(new_n890), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n892), .A2(new_n896), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n868), .B2(new_n571), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n854), .A2(new_n297), .A3(new_n825), .A4(new_n855), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1347gat));
  NAND4_X1  g699(.A1(new_n814), .A2(new_n631), .A3(new_n435), .A4(new_n415), .ZN(new_n901));
  INV_X1    g700(.A(G169gat), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(new_n263), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n836), .A2(new_n679), .ZN(new_n904));
  INV_X1    g703(.A(new_n722), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n415), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n817), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n903), .B1(new_n908), .B2(new_n902), .ZN(G1348gat));
  OR3_X1    g708(.A1(new_n906), .A2(G176gat), .A3(new_n627), .ZN(new_n910));
  OAI21_X1  g709(.A(G176gat), .B1(new_n901), .B2(new_n627), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1349gat));
  OAI21_X1  g711(.A(G183gat), .B1(new_n901), .B2(new_n652), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n595), .A2(new_n351), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n906), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(KEYINPUT126), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n915), .B(new_n917), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n907), .A2(new_n348), .A3(new_n570), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n901), .A2(new_n571), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n921), .A3(G190gat), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n920), .B2(G190gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(G1351gat));
  NOR3_X1   g724(.A1(new_n645), .A2(new_n333), .A3(new_n722), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n904), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(G197gat), .B1(new_n928), .B2(new_n817), .ZN(new_n929));
  INV_X1    g728(.A(new_n885), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n645), .A2(new_n679), .A3(new_n634), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n817), .A2(G197gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(G1352gat));
  NAND3_X1  g733(.A1(new_n930), .A2(new_n628), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G204gat), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n627), .A2(G204gat), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT62), .B1(new_n927), .B2(new_n937), .ZN(new_n938));
  OR3_X1    g737(.A1(new_n927), .A2(KEYINPUT62), .A3(new_n937), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(G1353gat));
  NAND3_X1  g739(.A1(new_n928), .A2(new_n269), .A3(new_n595), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n595), .B(new_n931), .C1(new_n883), .C2(new_n884), .ZN(new_n942));
  AND2_X1   g741(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n943));
  OAI21_X1  g742(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n943), .B1(new_n942), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n941), .B1(new_n946), .B2(new_n947), .ZN(G1354gat));
  NAND3_X1  g747(.A1(new_n930), .A2(new_n570), .A3(new_n931), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G218gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n928), .A2(new_n270), .A3(new_n570), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1355gat));
endmodule


