//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n597, new_n598, new_n600, new_n601, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n202));
  XOR2_X1   g001(.A(G1gat), .B(G29gat), .Z(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT73), .B(KEYINPUT0), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G57gat), .B(G85gat), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  XOR2_X1   g006(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n208));
  XNOR2_X1  g007(.A(G113gat), .B(G120gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT1), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n210), .B2(new_n209), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G134gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G127gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n212), .B(new_n214), .C1(G127gat), .C2(G134gat), .ZN(new_n215));
  INV_X1    g014(.A(G113gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G120gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT68), .B(G120gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(new_n216), .ZN(new_n219));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT1), .B1(new_n220), .B2(KEYINPUT69), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n219), .B(new_n221), .C1(KEYINPUT69), .C2(new_n220), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n215), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G141gat), .B(G148gat), .Z(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT2), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G155gat), .B(G162gat), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n228), .B(new_n229), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n228), .B(new_n229), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n222), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G225gat), .A2(G233gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n208), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n230), .A2(KEYINPUT3), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n232), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n223), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n237), .B1(new_n244), .B2(new_n236), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n236), .B1(new_n242), .B2(new_n243), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT74), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n208), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n246), .B2(new_n208), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n207), .B(new_n245), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n250), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n248), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n207), .B1(new_n255), .B2(new_n245), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n202), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n245), .B1(new_n249), .B2(new_n250), .ZN(new_n258));
  INV_X1    g057(.A(new_n207), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n260), .A2(KEYINPUT76), .A3(new_n252), .A4(new_n251), .ZN(new_n261));
  INV_X1    g060(.A(new_n252), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n257), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G8gat), .B(G36gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n265), .B(new_n266), .Z(new_n267));
  NAND2_X1  g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n268), .B(KEYINPUT64), .Z(new_n269));
  NOR2_X1   g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT23), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(G183gat), .B2(G190gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT65), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(KEYINPUT24), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT24), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(KEYINPUT65), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n272), .B(KEYINPUT25), .C1(new_n274), .C2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n274), .B1(new_n278), .B2(new_n275), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n282), .A2(new_n269), .A3(new_n271), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n283), .B2(KEYINPUT25), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT27), .B(G183gat), .ZN(new_n285));
  INV_X1    g084(.A(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n270), .B(KEYINPUT26), .Z(new_n290));
  OAI211_X1 g089(.A(new_n289), .B(new_n275), .C1(new_n269), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n292), .A2(new_n293), .B1(G226gat), .B2(G233gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G197gat), .B(G204gat), .ZN(new_n296));
  INV_X1    g095(.A(G211gat), .ZN(new_n297));
  INV_X1    g096(.A(G218gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n296), .B1(KEYINPUT22), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G211gat), .B(G218gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n292), .A2(G226gat), .A3(G233gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n295), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n304), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n302), .B1(new_n306), .B2(new_n294), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n267), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT30), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n307), .A3(new_n267), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT30), .A4(new_n267), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n312), .A2(new_n313), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n240), .A2(new_n293), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n302), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n239), .B1(new_n302), .B2(KEYINPUT29), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n230), .ZN(new_n321));
  AND2_X1   g120(.A1(G228gat), .A2(G233gat), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n322), .A2(KEYINPUT78), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(KEYINPUT78), .A3(new_n322), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(KEYINPUT78), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n319), .A2(new_n326), .A3(new_n321), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330));
  INV_X1    g129(.A(G50gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(KEYINPUT77), .B(KEYINPUT31), .Z(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n329), .A2(G22gat), .A3(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(KEYINPUT79), .B(G22gat), .Z(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n325), .B2(new_n327), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n329), .A2(new_n338), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n335), .A2(KEYINPUT80), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n328), .A2(new_n337), .A3(new_n341), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n336), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G15gat), .B(G43gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G71gat), .B(G99gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n292), .B(new_n223), .ZN(new_n348));
  INV_X1    g147(.A(G227gat), .ZN(new_n349));
  INV_X1    g148(.A(G233gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT33), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n347), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(KEYINPUT32), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT34), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n292), .B(new_n223), .Z(new_n358));
  INV_X1    g157(.A(new_n351), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n348), .A2(KEYINPUT34), .A3(new_n351), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n352), .B(KEYINPUT32), .C1(new_n353), .C2(new_n347), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n356), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n356), .B2(new_n363), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n344), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n264), .A2(new_n317), .A3(new_n366), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n367), .A2(KEYINPUT84), .A3(KEYINPUT35), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT84), .B1(new_n367), .B2(KEYINPUT35), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n207), .B(KEYINPUT81), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n255), .B2(new_n245), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n263), .B1(new_n371), .B2(new_n253), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n344), .A2(KEYINPUT35), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n364), .B2(new_n365), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n363), .ZN(new_n377));
  INV_X1    g176(.A(new_n362), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT70), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n374), .A2(new_n380), .A3(new_n316), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n368), .A2(new_n369), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n344), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n383), .B1(new_n264), .B2(new_n317), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n364), .A2(new_n365), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT36), .ZN(new_n387));
  INV_X1    g186(.A(new_n380), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(KEYINPUT36), .ZN(new_n389));
  NOR2_X1   g188(.A1(KEYINPUT82), .A2(KEYINPUT40), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n244), .A2(new_n236), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT39), .ZN(new_n392));
  INV_X1    g191(.A(new_n234), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(new_n235), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n244), .A2(new_n392), .A3(new_n236), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n370), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n390), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n391), .A2(new_n394), .ZN(new_n399));
  INV_X1    g198(.A(new_n390), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n399), .A2(new_n370), .A3(new_n400), .A4(new_n396), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n371), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(new_n316), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT83), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n305), .A2(new_n307), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n267), .B1(new_n406), .B2(KEYINPUT37), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(KEYINPUT37), .B2(new_n406), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n408), .A2(KEYINPUT38), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(KEYINPUT38), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n310), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n383), .B1(new_n411), .B2(new_n372), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n385), .B(new_n389), .C1(new_n405), .C2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n382), .A2(new_n414), .A3(KEYINPUT85), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n369), .A2(new_n381), .ZN(new_n417));
  INV_X1    g216(.A(new_n368), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n416), .B1(new_n419), .B2(new_n413), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(G43gat), .B(G50gat), .Z(new_n422));
  INV_X1    g221(.A(KEYINPUT15), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(G29gat), .A2(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT14), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n426), .A2(KEYINPUT87), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT88), .B(G29gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(G36gat), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n426), .B2(KEYINPUT87), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n424), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n424), .A2(new_n426), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n422), .A2(new_n423), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G15gat), .B(G22gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT16), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(G1gat), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(G1gat), .B2(new_n437), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n440), .B(G8gat), .Z(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT90), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n441), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n435), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n444), .B(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G229gat), .A2(G233gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n448), .B(KEYINPUT89), .Z(new_n449));
  XOR2_X1   g248(.A(new_n449), .B(KEYINPUT13), .Z(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT17), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n441), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n449), .A3(new_n446), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT18), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n457), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n461));
  XNOR2_X1  g260(.A(G113gat), .B(G141gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(G197gat), .ZN(new_n463));
  XOR2_X1   g262(.A(KEYINPUT11), .B(G169gat), .Z(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n465), .B(KEYINPUT12), .Z(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n460), .A2(new_n461), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n460), .B2(new_n461), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n421), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT95), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(G85gat), .A3(G92gat), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT7), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478));
  INV_X1    g277(.A(G85gat), .ZN(new_n479));
  INV_X1    g278(.A(G92gat), .ZN(new_n480));
  AOI22_X1  g279(.A1(KEYINPUT8), .A2(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n474), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(G99gat), .B(G106gat), .Z(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n484), .A2(new_n477), .A3(new_n481), .A4(new_n482), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n473), .B1(new_n436), .B2(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n489), .B(KEYINPUT96), .Z(new_n490));
  NAND3_X1  g289(.A1(new_n452), .A2(new_n454), .A3(new_n488), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XOR2_X1   g291(.A(G190gat), .B(G218gat), .Z(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT94), .ZN(new_n496));
  XNOR2_X1  g295(.A(G134gat), .B(G162gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n494), .A2(new_n499), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n504));
  NAND2_X1  g303(.A1(G71gat), .A2(G78gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT9), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G57gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n508), .A2(G64gat), .ZN(new_n509));
  INV_X1    g308(.A(G64gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(G57gat), .ZN(new_n511));
  OAI211_X1 g310(.A(KEYINPUT91), .B(new_n507), .C1(new_n509), .C2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G71gat), .B(G78gat), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(G57gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n508), .A2(G64gat), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n513), .B1(new_n519), .B2(new_n507), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n504), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n512), .A2(new_n514), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n513), .A3(new_n507), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT92), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT21), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(G127gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n441), .B1(new_n526), .B2(new_n525), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G183gat), .B(G211gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT93), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(new_n225), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n534), .B(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n532), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT10), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n525), .A2(new_n543), .A3(new_n488), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n484), .A2(KEYINPUT98), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n545), .A2(new_n483), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n515), .A2(new_n520), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n483), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n522), .A2(KEYINPUT92), .A3(new_n523), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT92), .B1(new_n522), .B2(new_n523), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n488), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n525), .A2(KEYINPUT97), .A3(new_n488), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n550), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n544), .B1(new_n557), .B2(new_n543), .ZN(new_n558));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT99), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n486), .A2(new_n487), .ZN(new_n562));
  AOI211_X1 g361(.A(new_n554), .B(new_n562), .C1(new_n524), .C2(new_n521), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT97), .B1(new_n525), .B2(new_n488), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n543), .B(new_n549), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n544), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT99), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n559), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n557), .A2(new_n559), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G120gat), .B(G148gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n567), .A2(new_n559), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(new_n571), .A3(new_n575), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n503), .A2(new_n542), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n472), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(new_n264), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(G1gat), .Z(G1324gat));
  NAND3_X1  g383(.A1(new_n472), .A2(new_n316), .A3(new_n581), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT100), .B(KEYINPUT16), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(G8gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT42), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(KEYINPUT42), .A3(new_n588), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n593), .B1(new_n585), .B2(G8gat), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n585), .A2(new_n593), .A3(G8gat), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n591), .B(new_n592), .C1(new_n594), .C2(new_n595), .ZN(G1325gat));
  OAI21_X1  g395(.A(G15gat), .B1(new_n582), .B2(new_n389), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n380), .A2(G15gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n582), .B2(new_n598), .ZN(G1326gat));
  NOR2_X1   g398(.A1(new_n582), .A2(new_n383), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT43), .B(G22gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(G1327gat));
  OAI21_X1  g401(.A(KEYINPUT85), .B1(new_n382), .B2(new_n414), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n419), .A2(new_n416), .A3(new_n413), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n580), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n542), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(new_n471), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n503), .A3(new_n608), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n609), .A2(new_n264), .A3(new_n428), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT45), .Z(new_n611));
  INV_X1    g410(.A(new_n608), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n503), .B1(new_n415), .B2(new_n420), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT44), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n382), .A2(new_n414), .A3(KEYINPUT102), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n616), .B1(new_n419), .B2(new_n413), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n502), .A2(KEYINPUT44), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n612), .B1(new_n614), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n428), .B1(new_n622), .B2(new_n264), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n611), .A2(new_n623), .ZN(G1328gat));
  OAI21_X1  g423(.A(G36gat), .B1(new_n622), .B2(new_n317), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n609), .A2(G36gat), .A3(new_n317), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT46), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(G1329gat));
  INV_X1    g427(.A(new_n389), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n621), .A2(G43gat), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G43gat), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(new_n609), .B2(new_n380), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT47), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT47), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n630), .A2(new_n635), .A3(new_n632), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(G1330gat));
  NAND3_X1  g436(.A1(new_n503), .A2(new_n331), .A3(new_n344), .ZN(new_n638));
  NOR4_X1   g437(.A1(new_n421), .A2(new_n471), .A3(new_n607), .A4(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT48), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n605), .B2(new_n503), .ZN(new_n643));
  INV_X1    g442(.A(new_n619), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n615), .A2(new_n617), .A3(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n344), .B(new_n608), .C1(new_n643), .C2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT103), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(G50gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n646), .A2(KEYINPUT103), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n641), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n331), .B1(new_n621), .B2(new_n344), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n640), .B1(new_n651), .B2(new_n639), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(G1331gat));
  NAND3_X1  g452(.A1(new_n502), .A2(new_n471), .A3(new_n541), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n606), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n618), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n264), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n508), .ZN(G1332gat));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n317), .ZN(new_n659));
  NOR2_X1   g458(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n660));
  AND2_X1   g459(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n659), .B2(new_n660), .ZN(G1333gat));
  OAI21_X1  g462(.A(G71gat), .B1(new_n656), .B2(new_n389), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n380), .A2(G71gat), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n656), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT104), .B(KEYINPUT50), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(G1334gat));
  NOR2_X1   g467(.A1(new_n656), .A2(new_n383), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g469(.A1(new_n541), .A2(new_n470), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n503), .B(new_n671), .C1(new_n382), .C2(new_n414), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT51), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT105), .ZN(new_n674));
  INV_X1    g473(.A(new_n264), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n674), .A2(new_n479), .A3(new_n675), .A4(new_n580), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n580), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n614), .B2(new_n620), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n678), .A2(new_n675), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n676), .B1(new_n479), .B2(new_n679), .ZN(G1336gat));
  INV_X1    g479(.A(new_n677), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n316), .B(new_n681), .C1(new_n643), .C2(new_n645), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(G92gat), .ZN(new_n683));
  INV_X1    g482(.A(new_n673), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n684), .A2(new_n480), .A3(new_n316), .A4(new_n580), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT106), .B(KEYINPUT52), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT107), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n683), .A2(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT52), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n683), .A2(new_n685), .A3(new_n691), .A4(new_n686), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n688), .A2(new_n690), .A3(new_n692), .ZN(G1337gat));
  XOR2_X1   g492(.A(KEYINPUT108), .B(G99gat), .Z(new_n694));
  NAND4_X1  g493(.A1(new_n674), .A2(new_n388), .A3(new_n580), .A4(new_n694), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n678), .A2(new_n629), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(G1338gat));
  NOR4_X1   g496(.A1(new_n673), .A2(G106gat), .A3(new_n383), .A4(new_n606), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n678), .A2(new_n344), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT109), .B(G106gat), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n699), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n700), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n678), .B2(new_n344), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(new_n698), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(G1339gat));
  NAND3_X1  g506(.A1(new_n675), .A2(new_n317), .A3(new_n366), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n561), .A2(new_n569), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT54), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n567), .B2(new_n559), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n558), .A2(new_n560), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n710), .A2(new_n576), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT55), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n712), .B2(new_n713), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n710), .A3(new_n576), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n718), .A2(new_n710), .A3(KEYINPUT112), .A4(new_n576), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT113), .B1(new_n723), .B2(new_n579), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT113), .ZN(new_n725));
  INV_X1    g524(.A(new_n579), .ZN(new_n726));
  AOI211_X1 g525(.A(new_n725), .B(new_n726), .C1(new_n721), .C2(new_n722), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n470), .B(new_n717), .C1(new_n724), .C2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n460), .A2(new_n466), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n447), .A2(new_n450), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n449), .B1(new_n455), .B2(new_n446), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n729), .B1(new_n465), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n580), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n728), .A2(KEYINPUT114), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT114), .B1(new_n728), .B2(new_n734), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n735), .A2(new_n736), .A3(new_n503), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n724), .A2(new_n727), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(new_n716), .B2(new_n715), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n503), .A2(new_n733), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n542), .B1(new_n737), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n654), .A2(new_n580), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n708), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT115), .Z(new_n747));
  NAND2_X1  g546(.A1(new_n470), .A2(new_n216), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(KEYINPUT116), .Z(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n344), .B1(new_n743), .B2(new_n745), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n264), .A2(new_n380), .A3(new_n316), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G113gat), .B1(new_n753), .B2(new_n471), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(new_n754), .ZN(G1340gat));
  INV_X1    g554(.A(new_n218), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n747), .A2(new_n756), .A3(new_n580), .ZN(new_n757));
  OAI21_X1  g556(.A(G120gat), .B1(new_n753), .B2(new_n606), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1341gat));
  OAI21_X1  g558(.A(G127gat), .B1(new_n753), .B2(new_n542), .ZN(new_n760));
  INV_X1    g559(.A(G127gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n761), .A3(new_n541), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT117), .ZN(G1342gat));
  INV_X1    g563(.A(new_n213), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n746), .A2(new_n765), .A3(new_n503), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n503), .A3(new_n752), .ZN(new_n767));
  AOI22_X1  g566(.A1(KEYINPUT56), .A2(new_n766), .B1(new_n767), .B2(G134gat), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n766), .A2(KEYINPUT56), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(KEYINPUT118), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(KEYINPUT118), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(G1343gat));
  INV_X1    g571(.A(G141gat), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n743), .A2(new_n745), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n629), .A2(new_n264), .A3(new_n316), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n344), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n773), .B1(new_n776), .B2(new_n471), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n775), .B(KEYINPUT119), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n728), .A2(new_n734), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n728), .A2(KEYINPUT114), .A3(new_n734), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n502), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n541), .B1(new_n784), .B2(new_n741), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n344), .B1(new_n785), .B2(new_n744), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT120), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n470), .A2(new_n717), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n723), .A2(new_n579), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n734), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT121), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n503), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n794), .A2(new_n795), .B1(new_n739), .B2(new_n740), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n745), .B1(new_n796), .B2(new_n541), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n383), .A2(new_n788), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n789), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n787), .B1(new_n786), .B2(new_n788), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n779), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n470), .A2(G141gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n777), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT58), .B(new_n777), .C1(new_n802), .C2(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1344gat));
  NOR3_X1   g607(.A1(new_n776), .A2(G148gat), .A3(new_n606), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT122), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G148gat), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n789), .A2(new_n799), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n786), .A2(new_n788), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT120), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n778), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n812), .B1(new_n816), .B2(new_n580), .ZN(new_n817));
  INV_X1    g616(.A(new_n798), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n743), .B2(new_n745), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT57), .B1(new_n797), .B2(new_n344), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n580), .B(new_n779), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n811), .B1(new_n821), .B2(G148gat), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n810), .B1(new_n817), .B2(new_n822), .ZN(G1345gat));
  OAI21_X1  g622(.A(G155gat), .B1(new_n802), .B2(new_n542), .ZN(new_n824));
  INV_X1    g623(.A(new_n776), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n225), .A3(new_n541), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(G1346gat));
  OAI211_X1 g626(.A(new_n503), .B(new_n779), .C1(new_n800), .C2(new_n801), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n799), .A3(new_n789), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n831), .A2(KEYINPUT123), .A3(new_n503), .A4(new_n779), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(G162gat), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n825), .A2(new_n226), .A3(new_n503), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1347gat));
  AOI21_X1  g634(.A(new_n675), .B1(new_n743), .B2(new_n745), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n366), .A2(new_n316), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(G169gat), .B1(new_n839), .B2(new_n470), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n675), .A2(new_n317), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n751), .A2(new_n388), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(G169gat), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n842), .A2(new_n843), .A3(new_n471), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n840), .A2(new_n844), .ZN(G1348gat));
  OAI21_X1  g644(.A(G176gat), .B1(new_n842), .B2(new_n606), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n606), .A2(G176gat), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n838), .B2(new_n847), .ZN(G1349gat));
  OAI21_X1  g647(.A(G183gat), .B1(new_n842), .B2(new_n542), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n541), .A2(new_n285), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT124), .B1(new_n839), .B2(new_n850), .ZN(new_n851));
  AND4_X1   g650(.A1(KEYINPUT124), .A2(new_n836), .A3(new_n837), .A4(new_n850), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT60), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT60), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n849), .B(new_n855), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1350gat));
  NAND3_X1  g656(.A1(new_n839), .A2(new_n286), .A3(new_n503), .ZN(new_n858));
  OAI21_X1  g657(.A(G190gat), .B1(new_n842), .B2(new_n502), .ZN(new_n859));
  XOR2_X1   g658(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n860));
  AND2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(G1351gat));
  NOR3_X1   g662(.A1(new_n629), .A2(new_n383), .A3(new_n317), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n836), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(G197gat), .B1(new_n866), .B2(new_n470), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n389), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n819), .B2(new_n820), .ZN(new_n870));
  INV_X1    g669(.A(G197gat), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n870), .A2(new_n871), .A3(new_n471), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n867), .A2(new_n872), .ZN(G1352gat));
  NOR3_X1   g672(.A1(new_n865), .A2(G204gat), .A3(new_n606), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G204gat), .B1(new_n870), .B2(new_n606), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G1353gat));
  NAND3_X1  g678(.A1(new_n866), .A2(new_n297), .A3(new_n541), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n541), .B(new_n869), .C1(new_n819), .C2(new_n820), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n881), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT63), .B1(new_n881), .B2(G211gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT126), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n886), .B(new_n880), .C1(new_n882), .C2(new_n883), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1354gat));
  OAI21_X1  g687(.A(G218gat), .B1(new_n870), .B2(new_n502), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n503), .A2(new_n298), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n865), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


