//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  AND2_X1   g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(KEYINPUT24), .ZN(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n208), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT23), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G169gat), .B2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT25), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G183gat), .B2(G190gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(new_n214), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT66), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n211), .B(new_n224), .C1(G183gat), .C2(G190gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n222), .A2(KEYINPUT25), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT65), .B1(new_n209), .B2(new_n210), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n227), .B1(new_n235), .B2(new_n215), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n231), .B(new_n233), .C1(new_n236), .C2(KEYINPUT25), .ZN(new_n237));
  XOR2_X1   g036(.A(G113gat), .B(G120gat), .Z(new_n238));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n239));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT68), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n238), .A2(new_n243), .A3(new_n239), .A4(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n239), .ZN(new_n245));
  INV_X1    g044(.A(new_n240), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n242), .A2(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n217), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n248), .A2(KEYINPUT26), .ZN(new_n249));
  INV_X1    g048(.A(new_n221), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n250), .B2(KEYINPUT26), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n207), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253));
  INV_X1    g052(.A(G183gat), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n254), .A2(KEYINPUT27), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(KEYINPUT27), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(KEYINPUT27), .ZN(new_n258));
  AOI21_X1  g057(.A(G190gat), .B1(new_n258), .B2(KEYINPUT67), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT28), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT27), .B(G183gat), .Z(new_n261));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n261), .A2(new_n262), .A3(G190gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n252), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n230), .A2(new_n237), .A3(new_n247), .A4(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n230), .A2(new_n237), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n242), .A2(new_n244), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n245), .A2(new_n246), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n266), .A3(new_n271), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n205), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G15gat), .B(G43gat), .Z(new_n276));
  XNOR2_X1  g075(.A(G71gat), .B(G99gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT33), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT32), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT33), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(KEYINPUT32), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n268), .A2(new_n266), .A3(new_n271), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n272), .B2(new_n267), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n288), .B2(new_n205), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n283), .B1(new_n289), .B2(new_n278), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n283), .B(new_n278), .C1(new_n275), .C2(new_n285), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n282), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n203), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT34), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n204), .A2(KEYINPUT34), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n293), .A2(KEYINPUT71), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n278), .B1(new_n275), .B2(new_n285), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT70), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n281), .B1(new_n302), .B2(new_n291), .ZN(new_n303));
  INV_X1    g102(.A(new_n298), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n304), .ZN(new_n306));
  AND4_X1   g105(.A1(KEYINPUT36), .A2(new_n299), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n308), .A3(new_n298), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT72), .B1(new_n303), .B2(new_n304), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(new_n306), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT36), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n307), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT30), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n264), .B1(new_n223), .B2(new_n229), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(KEYINPUT74), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT22), .ZN(new_n328));
  XNOR2_X1  g127(.A(G211gat), .B(G218gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G211gat), .ZN(new_n332));
  INV_X1    g131(.A(G218gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n329), .B(new_n327), .C1(KEYINPUT22), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n322), .A2(KEYINPUT75), .A3(new_n323), .ZN(new_n337));
  INV_X1    g136(.A(new_n323), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n268), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n326), .A2(new_n336), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n320), .A2(new_n323), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n338), .A2(KEYINPUT29), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n341), .B1(new_n268), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n336), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT76), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n318), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n349), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n340), .A2(new_n345), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(KEYINPUT30), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT5), .ZN(new_n358));
  XOR2_X1   g157(.A(G155gat), .B(G162gat), .Z(new_n359));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G148gat), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT77), .B1(new_n362), .B2(G141gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n364));
  INV_X1    g163(.A(G141gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(G148gat), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n363), .B(new_n366), .C1(new_n365), .C2(G148gat), .ZN(new_n367));
  INV_X1    g166(.A(G155gat), .ZN(new_n368));
  INV_X1    g167(.A(G162gat), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT2), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G155gat), .B(G162gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT78), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n361), .A2(new_n367), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G141gat), .B(G148gat), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n359), .B1(KEYINPUT2), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n247), .B(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n271), .B2(new_n376), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n373), .A2(new_n383), .A3(new_n375), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n271), .A3(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n247), .A2(KEYINPUT4), .A3(new_n373), .A4(new_n375), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n381), .A2(new_n385), .A3(new_n378), .A4(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n358), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT0), .ZN(new_n390));
  XOR2_X1   g189(.A(G57gat), .B(G85gat), .Z(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n387), .A2(new_n358), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n388), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT6), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n392), .B1(new_n388), .B2(new_n393), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(KEYINPUT79), .B(new_n392), .C1(new_n388), .C2(new_n393), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT6), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n396), .B1(new_n401), .B2(new_n394), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n357), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G78gat), .B(G106gat), .Z(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT31), .B(G50gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n335), .B(KEYINPUT80), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n410), .A2(new_n331), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n383), .B1(new_n411), .B2(KEYINPUT29), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n376), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n336), .B1(new_n384), .B2(new_n321), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n414), .B1(G228gat), .B2(G233gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n383), .B1(new_n344), .B2(KEYINPUT29), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n376), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n414), .B2(KEYINPUT81), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n414), .A2(KEYINPUT81), .ZN(new_n420));
  OAI211_X1 g219(.A(G228gat), .B(G233gat), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G22gat), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n416), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n416), .B2(new_n421), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n409), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT83), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n407), .A2(new_n408), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n428), .B(new_n409), .C1(new_n423), .C2(new_n424), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n426), .B2(new_n429), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n404), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n202), .B1(new_n317), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n307), .ZN(new_n437));
  INV_X1    g236(.A(new_n316), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n315), .B1(new_n311), .B2(new_n312), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(KEYINPUT84), .A3(new_n434), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n355), .B1(new_n353), .B2(new_n351), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n377), .A2(new_n378), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT39), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n444), .A2(KEYINPUT85), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(KEYINPUT85), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n381), .A2(new_n386), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n378), .B1(new_n447), .B2(new_n385), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT39), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n392), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(KEYINPUT40), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n454), .A2(KEYINPUT86), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(KEYINPUT86), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n394), .B1(new_n453), .B2(KEYINPUT40), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n442), .A2(new_n455), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n340), .A2(new_n345), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n343), .B2(new_n336), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n326), .A2(new_n337), .A3(new_n339), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(new_n336), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT87), .B(KEYINPUT38), .Z(new_n465));
  AND2_X1   g264(.A1(new_n350), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT88), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n461), .A2(new_n469), .A3(new_n464), .A4(new_n466), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n468), .A2(new_n402), .A3(new_n353), .A4(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n352), .B1(new_n459), .B2(new_n460), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n346), .A2(KEYINPUT37), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n432), .B(new_n458), .C1(new_n471), .C2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n436), .A2(new_n441), .A3(new_n475), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n433), .A2(KEYINPUT35), .A3(new_n311), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n404), .A2(KEYINPUT89), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n357), .B2(new_n403), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n305), .A2(new_n306), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n432), .A2(new_n482), .A3(new_n299), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT35), .B1(new_n483), .B2(new_n404), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT104), .ZN(new_n487));
  XNOR2_X1  g286(.A(G190gat), .B(G218gat), .ZN(new_n488));
  XOR2_X1   g287(.A(G43gat), .B(G50gat), .Z(new_n489));
  NOR2_X1   g288(.A1(G29gat), .A2(G36gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT14), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G36gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT91), .B(G29gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT15), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n489), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n490), .B(KEYINPUT14), .ZN(new_n498));
  INV_X1    g297(.A(new_n494), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(G36gat), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT15), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(KEYINPUT15), .A3(new_n489), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT17), .ZN(new_n505));
  NAND2_X1  g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT8), .ZN(new_n507));
  XOR2_X1   g306(.A(KEYINPUT101), .B(G85gat), .Z(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(G92gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT102), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G85gat), .A2(G92gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G99gat), .B(G106gat), .Z(new_n515));
  OR2_X1    g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n505), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n517), .A3(new_n504), .ZN(new_n520));
  NAND3_X1  g319(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n488), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n518), .ZN(new_n524));
  INV_X1    g323(.A(new_n488), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n524), .A2(new_n520), .A3(new_n521), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT100), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT99), .ZN(new_n530));
  XNOR2_X1  g329(.A(G134gat), .B(G162gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT103), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n527), .A2(KEYINPUT100), .A3(new_n532), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n532), .B1(new_n527), .B2(KEYINPUT100), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT100), .ZN(new_n540));
  AOI211_X1 g339(.A(new_n540), .B(new_n533), .C1(new_n523), .C2(new_n526), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n535), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT16), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(G1gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546));
  MUX2_X1   g345(.A(G1gat), .B(new_n545), .S(new_n546), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G8gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT21), .ZN(new_n549));
  XNOR2_X1  g348(.A(G71gat), .B(G78gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT95), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552));
  INV_X1    g351(.A(G71gat), .ZN(new_n553));
  INV_X1    g352(.A(G78gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G57gat), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n556), .A2(G64gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(G64gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(KEYINPUT96), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT96), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n563), .B2(new_n557), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(new_n555), .A3(new_n550), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n548), .B1(new_n549), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT98), .ZN(new_n568));
  XNOR2_X1  g367(.A(G127gat), .B(G155gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(KEYINPUT20), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n549), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(G231gat), .A3(G233gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n566), .A2(new_n549), .A3(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n576), .B1(new_n573), .B2(new_n575), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n571), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n578), .A2(new_n579), .A3(new_n571), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n568), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  INV_X1    g383(.A(new_n568), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n585), .A3(new_n580), .ZN(new_n586));
  XOR2_X1   g385(.A(G183gat), .B(G211gat), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n583), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n583), .B2(new_n586), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n487), .B1(new_n543), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n538), .A2(new_n542), .A3(new_n591), .A4(KEYINPUT104), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n504), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(new_n548), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n548), .B(KEYINPUT92), .Z(new_n598));
  AOI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(new_n505), .ZN(new_n599));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n600), .B(KEYINPUT93), .Z(new_n601));
  AND2_X1   g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n602), .A2(KEYINPUT18), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(KEYINPUT18), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n596), .A2(new_n548), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT94), .ZN(new_n606));
  MUX2_X1   g405(.A(new_n606), .B(KEYINPUT94), .S(new_n597), .Z(new_n607));
  XOR2_X1   g406(.A(new_n601), .B(KEYINPUT13), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n603), .A2(new_n604), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT11), .ZN(new_n612));
  INV_X1    g411(.A(G169gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT90), .B(G197gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n603), .A2(new_n604), .A3(new_n609), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n566), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n516), .A2(new_n623), .A3(new_n517), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT10), .B1(new_n624), .B2(KEYINPUT105), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n624), .A2(KEYINPUT105), .A3(KEYINPUT10), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n518), .A2(new_n566), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n629), .A2(new_n624), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n630), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT106), .ZN(new_n634));
  XOR2_X1   g433(.A(G176gat), .B(G204gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n632), .A2(KEYINPUT107), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n632), .B2(KEYINPUT107), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n595), .A2(new_n622), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT108), .B1(new_n486), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n486), .A2(KEYINPUT108), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n402), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g446(.A(KEYINPUT16), .B(G8gat), .Z(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n442), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(KEYINPUT42), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n645), .A2(new_n442), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n652), .B2(G8gat), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n650), .B1(new_n649), .B2(new_n653), .ZN(G1325gat));
  INV_X1    g453(.A(G15gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n644), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n642), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n655), .B1(new_n657), .B2(new_n311), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT109), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT109), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n660), .B(new_n655), .C1(new_n657), .C2(new_n311), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n317), .A2(G15gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT110), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n659), .A2(new_n661), .B1(new_n645), .B2(new_n663), .ZN(G1326gat));
  NAND2_X1  g463(.A1(new_n645), .A2(new_n433), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT43), .B(G22gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  INV_X1    g466(.A(new_n543), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n476), .B2(new_n485), .ZN(new_n669));
  INV_X1    g468(.A(new_n640), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n621), .A2(new_n592), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n402), .A3(new_n494), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT45), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n486), .A2(KEYINPUT44), .A3(new_n543), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n475), .A2(new_n434), .A3(new_n440), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n485), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n543), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n676), .A2(new_n681), .A3(new_n672), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT111), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n676), .A2(KEYINPUT111), .A3(new_n681), .A4(new_n672), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n684), .A2(new_n402), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n675), .B1(new_n494), .B2(new_n686), .ZN(G1328gat));
  NAND3_X1  g486(.A1(new_n673), .A2(new_n493), .A3(new_n442), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT46), .Z(new_n689));
  NAND3_X1  g488(.A1(new_n684), .A2(new_n442), .A3(new_n685), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G36gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(G1329gat));
  INV_X1    g491(.A(KEYINPUT113), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n682), .B2(new_n440), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n668), .B1(new_n677), .B2(new_n485), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(KEYINPUT44), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(KEYINPUT44), .B2(new_n669), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n697), .A2(KEYINPUT113), .A3(new_n317), .A4(new_n672), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n694), .A2(new_n698), .A3(G43gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n311), .A2(G43gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n669), .A2(new_n672), .A3(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(KEYINPUT47), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n701), .B(KEYINPUT112), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n684), .A2(new_n317), .A3(new_n685), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(G43gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n703), .B1(new_n706), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g506(.A(G50gat), .B1(new_n682), .B2(new_n432), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n432), .A2(G50gat), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT114), .Z(new_n710));
  NAND2_X1  g509(.A1(new_n673), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n708), .A2(KEYINPUT48), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n711), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n684), .A2(new_n433), .A3(new_n685), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(G50gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n712), .B1(new_n715), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g515(.A1(new_n595), .A2(new_n621), .A3(new_n670), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n678), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n403), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(new_n556), .ZN(G1332gat));
  NOR2_X1   g519(.A1(new_n718), .A2(KEYINPUT115), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT115), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n678), .B2(new_n717), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n442), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  AND2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n726), .B2(new_n725), .ZN(G1333gat));
  NOR3_X1   g528(.A1(new_n718), .A2(G71gat), .A3(new_n311), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n724), .A2(new_n317), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(G71gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g532(.A1(new_n724), .A2(new_n433), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT116), .B(G78gat), .Z(new_n735));
  XOR2_X1   g534(.A(new_n734), .B(new_n735), .Z(G1335gat));
  NOR2_X1   g535(.A1(new_n621), .A2(new_n591), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n695), .A2(KEYINPUT51), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT51), .B1(new_n695), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OR4_X1    g539(.A1(new_n403), .A2(new_n740), .A3(new_n508), .A4(new_n670), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n621), .A2(new_n670), .A3(new_n591), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n697), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n508), .B1(new_n743), .B2(new_n403), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(G1336gat));
  NOR3_X1   g544(.A1(new_n670), .A2(G92gat), .A3(new_n357), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n738), .B2(new_n739), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT118), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n676), .A2(new_n442), .A3(new_n681), .A4(new_n742), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G92gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n747), .A2(KEYINPUT117), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n754), .B(new_n746), .C1(new_n738), .C2(new_n739), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT52), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n752), .A2(new_n757), .ZN(G1337gat));
  OAI21_X1  g557(.A(G99gat), .B1(new_n743), .B2(new_n440), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n670), .A2(new_n311), .A3(G99gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n740), .B2(new_n760), .ZN(G1338gat));
  NAND4_X1  g560(.A1(new_n676), .A2(new_n433), .A3(new_n681), .A4(new_n742), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G106gat), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n432), .A2(G106gat), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n640), .B(new_n764), .C1(new_n738), .C2(new_n739), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g566(.A1(new_n593), .A2(new_n594), .A3(new_n622), .A4(new_n670), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT119), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n768), .A2(KEYINPUT119), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n628), .A2(new_n629), .ZN(new_n771));
  INV_X1    g570(.A(new_n627), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n771), .A2(new_n772), .A3(new_n625), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n637), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n772), .B1(new_n771), .B2(new_n625), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n630), .A3(KEYINPUT54), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT121), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT121), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n776), .A2(new_n778), .A3(new_n782), .A4(KEYINPUT55), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n632), .A2(new_n636), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n779), .B2(new_n780), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n621), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n607), .A2(new_n608), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n599), .A2(new_n601), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n616), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n640), .A2(new_n620), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n543), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n620), .A2(new_n790), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n538), .B2(new_n542), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n784), .A3(new_n786), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT122), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT122), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n794), .A2(new_n797), .A3(new_n784), .A4(new_n786), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n792), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n769), .B(new_n770), .C1(new_n799), .C2(new_n591), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n442), .A2(new_n403), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n433), .A2(new_n311), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(G113gat), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n804), .A2(new_n805), .A3(new_n622), .ZN(new_n806));
  INV_X1    g605(.A(new_n483), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n621), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n806), .B1(new_n805), .B2(new_n810), .ZN(G1340gat));
  INV_X1    g610(.A(G120gat), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n804), .A2(new_n812), .A3(new_n670), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n640), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n812), .B2(new_n814), .ZN(G1341gat));
  OAI21_X1  g614(.A(G127gat), .B1(new_n804), .B2(new_n592), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n592), .A2(G127gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n808), .B2(new_n817), .ZN(G1342gat));
  NOR3_X1   g617(.A1(new_n483), .A2(new_n668), .A3(G134gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT56), .Z(new_n821));
  OAI21_X1  g620(.A(G134gat), .B1(new_n804), .B2(new_n668), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1343gat));
  INV_X1    g622(.A(KEYINPUT123), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n440), .A2(new_n801), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n622), .A2(new_n365), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n796), .A2(new_n798), .ZN(new_n828));
  INV_X1    g627(.A(new_n792), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n591), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n768), .B(KEYINPUT119), .ZN(new_n831));
  OAI211_X1 g630(.A(KEYINPUT57), .B(new_n433), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT57), .B1(new_n800), .B2(new_n433), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n826), .B(new_n827), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n317), .A2(new_n432), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n800), .A2(new_n801), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n365), .B1(new_n837), .B2(new_n622), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n824), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI211_X1 g640(.A(KEYINPUT123), .B(KEYINPUT58), .C1(new_n835), .C2(new_n838), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n841), .A2(new_n842), .B1(new_n840), .B2(new_n839), .ZN(G1344gat));
  INV_X1    g642(.A(new_n837), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n362), .A3(new_n640), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(G148gat), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n833), .A2(new_n834), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n825), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n847), .B1(new_n849), .B2(new_n640), .ZN(new_n850));
  INV_X1    g649(.A(new_n795), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n592), .B1(new_n792), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n768), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n433), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n832), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n825), .B(KEYINPUT124), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n640), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n846), .B1(new_n859), .B2(G148gat), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n845), .B1(new_n850), .B2(new_n860), .ZN(G1345gat));
  AOI21_X1  g660(.A(G155gat), .B1(new_n844), .B2(new_n591), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n591), .A2(G155gat), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT125), .Z(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n849), .B2(new_n864), .ZN(G1346gat));
  NAND3_X1  g664(.A1(new_n844), .A2(new_n369), .A3(new_n543), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n848), .A2(new_n668), .A3(new_n825), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n369), .ZN(G1347gat));
  NOR2_X1   g667(.A1(new_n357), .A2(new_n402), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n800), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n803), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(new_n613), .A3(new_n622), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n807), .A3(new_n621), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n613), .B2(new_n873), .ZN(G1348gat));
  OAI21_X1  g673(.A(G176gat), .B1(new_n871), .B2(new_n670), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n870), .A2(new_n807), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n670), .A2(G176gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(G1349gat));
  OR3_X1    g677(.A1(new_n876), .A2(new_n261), .A3(new_n592), .ZN(new_n879));
  OAI21_X1  g678(.A(G183gat), .B1(new_n871), .B2(new_n592), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT60), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT60), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n879), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1350gat));
  OR3_X1    g684(.A1(new_n876), .A2(G190gat), .A3(new_n668), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n543), .A3(new_n803), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(G190gat), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n889), .A2(KEYINPUT126), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n887), .A3(G190gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n891), .B1(new_n889), .B2(KEYINPUT126), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n886), .B1(new_n890), .B2(new_n892), .ZN(G1351gat));
  INV_X1    g692(.A(new_n869), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n317), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n857), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G197gat), .B1(new_n896), .B2(new_n622), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n870), .A2(new_n836), .ZN(new_n898));
  INV_X1    g697(.A(G197gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n899), .A3(new_n621), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(G1352gat));
  INV_X1    g700(.A(G204gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n898), .A2(new_n902), .A3(new_n640), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n857), .A2(new_n640), .A3(new_n895), .ZN(new_n907));
  OAI22_X1  g706(.A1(new_n905), .A2(new_n906), .B1(new_n902), .B2(new_n907), .ZN(G1353gat));
  NAND3_X1  g707(.A1(new_n857), .A2(new_n591), .A3(new_n895), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT127), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n909), .A2(new_n912), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(G211gat), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT63), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n911), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n898), .A2(new_n332), .A3(new_n591), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1354gat));
  OAI21_X1  g718(.A(G218gat), .B1(new_n896), .B2(new_n668), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n898), .A2(new_n333), .A3(new_n543), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1355gat));
endmodule


