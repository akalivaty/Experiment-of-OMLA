//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT26), .B(G101), .Z(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n191), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT2), .B(G113), .Z(new_n195));
  OR2_X1    g009(.A1(new_n195), .A2(KEYINPUT68), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(KEYINPUT68), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G116), .ZN(new_n200));
  INV_X1    g014(.A(G116), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G119), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n198), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n200), .A2(new_n202), .A3(new_n198), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n196), .B(new_n197), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G116), .B(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n195), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT65), .A3(G146), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n213), .B2(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n211), .A2(KEYINPUT64), .A3(G143), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n215), .A2(new_n219), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n212), .A2(new_n217), .A3(new_n214), .A4(new_n218), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT66), .B1(new_n224), .B2(new_n221), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n211), .A2(G143), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n213), .A2(G146), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n229), .A2(new_n222), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n233));
  INV_X1    g047(.A(G134), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(G137), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(G137), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT11), .A3(G134), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  INV_X1    g054(.A(G131), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n235), .A2(new_n238), .A3(new_n241), .A4(new_n236), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n226), .A2(new_n232), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT67), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n231), .B1(new_n223), .B2(new_n225), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n243), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n242), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n237), .A2(G134), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n241), .B1(new_n236), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n215), .A2(new_n219), .A3(new_n253), .A4(G128), .ZN(new_n254));
  OAI21_X1  g068(.A(G128), .B1(new_n228), .B2(new_n253), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n227), .B2(new_n228), .ZN(new_n256));
  AOI211_X1 g070(.A(new_n250), .B(new_n252), .C1(new_n254), .C2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n209), .B1(new_n249), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n244), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n246), .A2(KEYINPUT70), .A3(new_n243), .ZN(new_n262));
  AOI211_X1 g076(.A(new_n208), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT28), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n257), .B1(new_n246), .B2(new_n243), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT28), .B1(new_n265), .B2(new_n209), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n194), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT30), .ZN(new_n269));
  AND4_X1   g083(.A1(new_n247), .A2(new_n226), .A3(new_n232), .A4(new_n243), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n247), .B1(new_n246), .B2(new_n243), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n269), .B(new_n258), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(new_n269), .ZN(new_n274));
  AOI211_X1 g088(.A(new_n263), .B(new_n193), .C1(new_n274), .C2(new_n208), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n187), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n273), .A2(new_n209), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT28), .B1(new_n278), .B2(new_n263), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n279), .A2(KEYINPUT29), .A3(new_n267), .A4(new_n193), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT72), .ZN(new_n281));
  INV_X1    g095(.A(new_n262), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT70), .B1(new_n246), .B2(new_n243), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n258), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n208), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n273), .A2(new_n209), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n266), .B1(new_n287), .B2(KEYINPUT28), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT29), .A4(new_n193), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n276), .A2(new_n277), .A3(new_n281), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G472), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n261), .A2(new_n262), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n269), .B1(new_n293), .B2(new_n258), .ZN(new_n294));
  AOI211_X1 g108(.A(KEYINPUT30), .B(new_n257), .C1(new_n245), .C2(new_n248), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n208), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n286), .A3(new_n193), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT31), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n264), .A2(new_n267), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n194), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n263), .B1(new_n274), .B2(new_n208), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT31), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n193), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n305), .B1(new_n304), .B2(new_n306), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n292), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT16), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(G125), .A2(G140), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n211), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n314), .ZN(new_n318));
  NOR2_X1   g132(.A1(G125), .A2(G140), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT16), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n316), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G146), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT24), .B(G110), .Z(new_n324));
  XNOR2_X1  g138(.A(G119), .B(G128), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n199), .B2(G128), .ZN(new_n328));
  INV_X1    g142(.A(G128), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT23), .A3(G119), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n328), .B(new_n330), .C1(G119), .C2(new_n329), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT73), .ZN(new_n332));
  INV_X1    g146(.A(G110), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n323), .B(new_n326), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(G146), .B1(new_n313), .B2(new_n314), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT74), .ZN(new_n336));
  OAI22_X1  g150(.A1(new_n331), .A2(G110), .B1(new_n325), .B2(new_n324), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n322), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G953), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(G221), .A3(G234), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT22), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(G137), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n344), .B(KEYINPUT75), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n345), .B(new_n346), .C1(new_n340), .C2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n340), .A2(KEYINPUT76), .A3(new_n344), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(KEYINPUT77), .B(KEYINPUT25), .C1(new_n350), .C2(G902), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  AOI21_X1  g166(.A(G902), .B1(new_n348), .B2(new_n349), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n277), .A2(G234), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n351), .A2(G217), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n350), .ZN(new_n358));
  AOI21_X1  g172(.A(G902), .B1(new_n356), .B2(G217), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n309), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G469), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(G107), .ZN(new_n366));
  INV_X1    g180(.A(G107), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(G104), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(KEYINPUT79), .A3(G104), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G101), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT80), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT3), .B1(new_n365), .B2(G107), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n367), .A3(G104), .ZN(new_n375));
  INV_X1    g189(.A(G101), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n365), .A2(G107), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n373), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n367), .A2(G104), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n379), .A3(new_n364), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT80), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G101), .A4(new_n370), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n372), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n224), .A2(new_n255), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n254), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n372), .A2(new_n378), .A3(new_n382), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n256), .A3(new_n254), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT12), .B1(new_n389), .B2(new_n243), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT12), .ZN(new_n391));
  INV_X1    g205(.A(new_n243), .ZN(new_n392));
  AOI211_X1 g206(.A(new_n391), .B(new_n392), .C1(new_n386), .C2(new_n388), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n373), .A2(new_n375), .A3(new_n377), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT78), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT78), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n373), .A2(new_n375), .A3(new_n397), .A4(new_n377), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(G101), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n378), .A2(KEYINPUT4), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n396), .A2(KEYINPUT4), .A3(G101), .A4(new_n398), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n246), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT10), .ZN(new_n405));
  INV_X1    g219(.A(new_n385), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(new_n387), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n254), .A2(new_n256), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n383), .A2(new_n408), .A3(KEYINPUT10), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n404), .A2(new_n407), .A3(new_n392), .A4(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G140), .ZN(new_n411));
  INV_X1    g225(.A(G227), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(G953), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n411), .B(new_n413), .Z(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n394), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n404), .A2(new_n407), .A3(new_n409), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n243), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n414), .B1(new_n418), .B2(new_n410), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n363), .B(new_n277), .C1(new_n416), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(G469), .A2(G902), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n410), .B1(new_n390), .B2(new_n393), .ZN(new_n422));
  INV_X1    g236(.A(new_n414), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n418), .A2(new_n410), .A3(new_n414), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(G469), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n420), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT9), .B(G234), .Z(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G221), .B1(new_n430), .B2(G902), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n427), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n428), .B1(new_n427), .B2(new_n431), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n362), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT89), .ZN(new_n437));
  XNOR2_X1  g251(.A(G113), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(new_n365), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n441));
  AOI21_X1  g255(.A(G143), .B1(new_n189), .B2(G214), .ZN(new_n442));
  OAI211_X1 g256(.A(KEYINPUT17), .B(G131), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n317), .A3(new_n322), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G237), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n341), .A3(G214), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n213), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G131), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n441), .A2(new_n442), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n241), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT17), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n443), .A2(new_n317), .A3(KEYINPUT86), .A4(new_n322), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n446), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT18), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n449), .B1(new_n457), .B2(new_n241), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n451), .A2(KEYINPUT18), .A3(G131), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n313), .A2(G146), .A3(new_n314), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n336), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n456), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n464), .B1(new_n456), .B2(new_n463), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n437), .B(new_n440), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n456), .A2(new_n463), .A3(new_n439), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n456), .A2(new_n463), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT88), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n465), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n437), .B1(new_n473), .B2(new_n440), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n277), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n341), .A2(G952), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(G234), .B2(G237), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT21), .B(G898), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT93), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n277), .B(new_n341), .C1(G234), .C2(G237), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G128), .B(G143), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT13), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n213), .A2(G128), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n486), .B(G134), .C1(KEYINPUT13), .C2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(G116), .B(G122), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(new_n367), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n234), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n485), .B(new_n234), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n367), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT14), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n201), .A2(KEYINPUT14), .A3(G122), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(G107), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n429), .A2(G217), .A3(new_n341), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(KEYINPUT91), .A3(new_n501), .ZN(new_n505));
  INV_X1    g319(.A(new_n500), .ZN(new_n506));
  INV_X1    g320(.A(new_n501), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT90), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n500), .A2(new_n509), .A3(new_n501), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n504), .B(new_n505), .C1(new_n508), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n277), .ZN(new_n512));
  AND2_X1   g326(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n513));
  NOR2_X1   g327(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n514));
  OAI21_X1  g328(.A(G478), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n512), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n313), .A2(new_n314), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT19), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n322), .B1(new_n519), .B2(G146), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n450), .B2(new_n452), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n458), .A2(new_n459), .B1(new_n336), .B2(new_n461), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n440), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n469), .ZN(new_n524));
  NOR2_X1   g338(.A1(G475), .A2(G902), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n525), .B(KEYINPUT87), .Z(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT20), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n476), .A2(new_n484), .A3(new_n516), .A4(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT20), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n527), .B(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n475), .B2(G475), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n534), .A2(KEYINPUT94), .A3(new_n484), .A4(new_n516), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G214), .B1(G237), .B2(G902), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  MUX2_X1   g352(.A(new_n408), .B(new_n246), .S(G125), .Z(new_n539));
  INV_X1    g353(.A(G224), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT7), .B1(new_n540), .B2(G953), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n539), .B(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G113), .B1(new_n200), .B2(KEYINPUT5), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n543), .B(KEYINPUT85), .Z(new_n544));
  AND2_X1   g358(.A1(new_n206), .A2(KEYINPUT5), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n207), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n383), .ZN(new_n547));
  XOR2_X1   g361(.A(G110), .B(G122), .Z(new_n548));
  XOR2_X1   g362(.A(new_n548), .B(KEYINPUT8), .Z(new_n549));
  INV_X1    g363(.A(KEYINPUT5), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n204), .A2(new_n203), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n207), .B1(new_n551), .B2(new_n543), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n547), .B(new_n549), .C1(new_n552), .C2(new_n383), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n403), .A2(new_n208), .ZN(new_n554));
  INV_X1    g368(.A(new_n548), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT82), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n552), .B2(new_n387), .ZN(new_n557));
  INV_X1    g371(.A(new_n203), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n206), .A2(new_n198), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(KEYINPUT5), .ZN(new_n560));
  INV_X1    g374(.A(new_n543), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n383), .A2(KEYINPUT82), .A3(new_n207), .A4(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n554), .A2(new_n555), .A3(new_n557), .A4(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT83), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n542), .B(new_n553), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n557), .A2(new_n563), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n555), .B1(new_n569), .B2(new_n554), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(KEYINPUT6), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n554), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n548), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n566), .B2(new_n567), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n571), .B1(new_n574), .B2(KEYINPUT6), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n540), .A2(G953), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT84), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n539), .B(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n277), .B(new_n568), .C1(new_n575), .C2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G210), .B1(G237), .B2(G902), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n571), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n564), .A2(new_n565), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n569), .A2(KEYINPUT83), .A3(new_n555), .A4(new_n554), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n570), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT6), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n578), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n590), .A2(new_n277), .A3(new_n580), .A4(new_n568), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n538), .B1(new_n582), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n536), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n436), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT95), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(new_n376), .ZN(G3));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n582), .A2(new_n597), .A3(new_n591), .ZN(new_n598));
  AOI21_X1  g412(.A(G902), .B1(new_n588), .B2(new_n589), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n599), .A2(KEYINPUT96), .A3(new_n580), .A4(new_n568), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n598), .A2(new_n484), .A3(new_n537), .A4(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n502), .A2(KEYINPUT98), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n500), .B1(new_n603), .B2(new_n501), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n511), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT97), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT97), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n511), .A2(new_n609), .A3(new_n605), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n606), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n277), .A2(G478), .ZN(new_n612));
  AOI21_X1  g426(.A(G478), .B1(new_n511), .B2(new_n277), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n613), .A2(KEYINPUT99), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(KEYINPUT99), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n611), .A2(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n534), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n601), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n304), .A2(new_n277), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n620), .A2(G472), .B1(new_n304), .B2(new_n306), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n434), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n357), .A2(new_n360), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  INV_X1    g441(.A(new_n516), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n534), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n601), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n624), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  INV_X1    g447(.A(KEYINPUT36), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n347), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n340), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n359), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n357), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n536), .A2(new_n592), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n622), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT37), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G110), .ZN(G12));
  AND2_X1   g456(.A1(new_n357), .A2(new_n637), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n304), .A2(new_n306), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT32), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n643), .B1(new_n647), .B2(new_n292), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n598), .A2(new_n537), .A3(new_n600), .ZN(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n478), .B1(new_n482), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n629), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n648), .A2(new_n649), .A3(new_n434), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  AND2_X1   g468(.A1(new_n582), .A2(new_n591), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT100), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n476), .A2(new_n528), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n628), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n301), .A2(new_n194), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n277), .B1(new_n287), .B2(new_n193), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n638), .B1(new_n647), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n651), .B(KEYINPUT39), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n435), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT40), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n661), .A2(new_n537), .A3(new_n665), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  INV_X1    g484(.A(new_n651), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n617), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n648), .A2(new_n649), .A3(new_n434), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  OR2_X1    g489(.A1(new_n416), .A2(new_n419), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n277), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(G469), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n678), .A2(new_n431), .A3(new_n420), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n309), .A2(new_n361), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n619), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT41), .B(G113), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT101), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G15));
  NAND2_X1  g498(.A1(new_n680), .A2(new_n630), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NAND4_X1  g500(.A1(new_n598), .A2(new_n537), .A3(new_n600), .A4(new_n679), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n536), .A3(new_n648), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  OAI211_X1 g504(.A(new_n298), .B(new_n303), .C1(new_n193), .C2(new_n288), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n306), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT102), .B1(new_n620), .B2(G472), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n694));
  INV_X1    g508(.A(G472), .ZN(new_n695));
  AOI211_X1 g509(.A(new_n694), .B(new_n695), .C1(new_n304), .C2(new_n277), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n692), .B(new_n361), .C1(new_n693), .C2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n679), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n659), .A2(KEYINPUT103), .A3(new_n628), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n534), .B2(new_n516), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n598), .A3(new_n537), .A4(new_n600), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n483), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  OAI211_X1 g521(.A(new_n692), .B(new_n638), .C1(new_n693), .C2(new_n696), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n708), .A2(new_n687), .A3(new_n672), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n311), .ZN(G27));
  AOI21_X1  g524(.A(new_n623), .B1(new_n647), .B2(new_n292), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n427), .A2(new_n431), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n582), .A2(new_n712), .A3(new_n537), .A4(new_n591), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n711), .B(new_n673), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(KEYINPUT105), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n713), .B(KEYINPUT104), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(KEYINPUT105), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n711), .A3(new_n673), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G131), .ZN(G33));
  OAI211_X1 g537(.A(new_n711), .B(new_n652), .C1(new_n714), .C2(new_n715), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT106), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n719), .A2(new_n726), .A3(new_n711), .A4(new_n652), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G134), .ZN(G36));
  NAND2_X1  g543(.A1(new_n611), .A2(new_n612), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n614), .A2(new_n615), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n534), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n733), .B(KEYINPUT43), .Z(new_n734));
  INV_X1    g548(.A(new_n621), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n638), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT44), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n655), .A2(new_n537), .ZN(new_n738));
  XOR2_X1   g552(.A(new_n738), .B(KEYINPUT107), .Z(new_n739));
  AND2_X1   g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n424), .A2(new_n425), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G469), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n421), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n745), .B(G469), .C1(new_n742), .C2(G902), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n420), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n431), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n666), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n740), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G137), .ZN(G39));
  NOR4_X1   g565(.A1(new_n738), .A2(new_n309), .A3(new_n361), .A4(new_n672), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT108), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n748), .B(KEYINPUT47), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n755), .B(KEYINPUT109), .Z(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n734), .A2(new_n478), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT114), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n738), .A2(new_n698), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n647), .A2(new_n361), .A3(new_n664), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n764), .A3(new_n478), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n765), .A2(new_n659), .ZN(new_n766));
  OAI22_X1  g580(.A1(new_n762), .A2(new_n708), .B1(new_n732), .B2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n760), .A2(new_n658), .A3(new_n538), .A4(new_n699), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n697), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n760), .A2(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n678), .A2(new_n420), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n754), .B1(new_n431), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n776), .A2(new_n739), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n758), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n776), .A2(new_n688), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n773), .A2(KEYINPUT51), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n783), .B(new_n767), .C1(new_n770), .C2(new_n771), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n780), .A2(KEYINPUT51), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n477), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n781), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n762), .A2(new_n362), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT48), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n765), .A2(new_n618), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n787), .A2(new_n788), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n781), .A2(new_n792), .A3(new_n782), .A4(new_n786), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT116), .B1(new_n794), .B2(new_n790), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n718), .A2(new_n721), .B1(new_n725), .B2(new_n727), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n640), .B1(new_n699), .B2(new_n705), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n629), .B1(new_n534), .B2(new_n616), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n434), .A2(new_n621), .A3(new_n361), .A4(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n592), .A2(new_n484), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n680), .A2(new_n630), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n799), .A2(new_n803), .A3(new_n689), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n738), .A2(new_n651), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n659), .A2(new_n628), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n434), .A4(new_n309), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n719), .A2(new_n673), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n692), .B1(new_n693), .B2(new_n696), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n638), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n436), .A2(new_n593), .B1(new_n680), .B2(new_n619), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n798), .A2(new_n804), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n712), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n704), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n671), .A3(new_n665), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n687), .A2(new_n672), .ZN(new_n817));
  INV_X1    g631(.A(new_n708), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n816), .A2(new_n819), .A3(new_n653), .A4(new_n674), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n309), .A2(new_n434), .A3(new_n638), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n598), .A2(new_n537), .A3(new_n600), .ZN(new_n824));
  INV_X1    g638(.A(new_n652), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n709), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(KEYINPUT52), .A3(new_n674), .A4(new_n816), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n797), .B(new_n813), .C1(new_n822), .C2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT111), .B1(new_n826), .B2(new_n709), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n665), .A2(new_n671), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n821), .B1(new_n831), .B2(new_n815), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n819), .A2(new_n833), .A3(new_n653), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n830), .A2(new_n674), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n835), .A2(new_n822), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n813), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(KEYINPUT53), .ZN(new_n838));
  OR3_X1    g652(.A1(new_n829), .A2(new_n838), .A3(KEYINPUT112), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n829), .A2(KEYINPUT112), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(KEYINPUT54), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT113), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT53), .B1(new_n836), .B2(new_n813), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n722), .A2(new_n728), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n812), .A2(new_n799), .A3(new_n689), .A4(new_n803), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n822), .A2(new_n828), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n797), .A3(new_n847), .A4(new_n811), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n839), .A2(new_n852), .A3(KEYINPUT54), .A4(new_n840), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n842), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n796), .A2(new_n854), .B1(G952), .B2(G953), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n778), .A2(KEYINPUT49), .ZN(new_n856));
  INV_X1    g670(.A(new_n733), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n537), .A2(new_n856), .A3(new_n431), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n778), .A2(KEYINPUT49), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n658), .A2(new_n858), .A3(new_n764), .A4(new_n859), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT110), .Z(new_n861));
  NAND2_X1  g675(.A1(new_n855), .A2(new_n861), .ZN(G75));
  NOR2_X1   g676(.A1(new_n849), .A2(new_n277), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT56), .B1(new_n863), .B2(G210), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n575), .A2(new_n578), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n590), .ZN(new_n866));
  XOR2_X1   g680(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n867));
  XNOR2_X1  g681(.A(new_n866), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n864), .B(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n341), .A2(G952), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT118), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n869), .A2(new_n872), .ZN(G51));
  NAND3_X1  g687(.A1(new_n843), .A2(KEYINPUT54), .A3(new_n848), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n851), .A2(KEYINPUT119), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n849), .A2(new_n876), .A3(new_n850), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n421), .B(KEYINPUT57), .Z(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n676), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT120), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n863), .A2(G469), .A3(new_n742), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n872), .B1(new_n881), .B2(new_n882), .ZN(G54));
  NAND3_X1  g697(.A1(new_n863), .A2(KEYINPUT58), .A3(G475), .ZN(new_n884));
  INV_X1    g698(.A(new_n524), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT121), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n884), .A2(new_n885), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n887), .A2(new_n872), .A3(new_n888), .ZN(G60));
  NAND2_X1  g703(.A1(G478), .A2(G902), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT59), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n611), .B1(new_n854), .B2(new_n891), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n611), .A2(new_n875), .A3(new_n877), .A4(new_n891), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n872), .A3(new_n893), .ZN(G63));
  NAND2_X1  g708(.A1(G217), .A2(G902), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT60), .Z(new_n896));
  NAND3_X1  g710(.A1(new_n843), .A2(new_n848), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n350), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n871), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n900));
  AND4_X1   g714(.A1(new_n636), .A2(new_n843), .A3(new_n848), .A4(new_n896), .ZN(new_n901));
  OR3_X1    g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n872), .B1(new_n897), .B2(new_n350), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n901), .B1(new_n906), .B2(KEYINPUT122), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n903), .B1(new_n908), .B2(new_n900), .ZN(new_n909));
  AOI211_X1 g723(.A(KEYINPUT123), .B(KEYINPUT61), .C1(new_n905), .C2(new_n907), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n902), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n913), .B(new_n902), .C1(new_n909), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(G66));
  NAND2_X1  g729(.A1(new_n845), .A2(new_n341), .ZN(new_n916));
  OAI21_X1  g730(.A(G953), .B1(new_n481), .B2(new_n540), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT125), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n917), .A2(KEYINPUT125), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n575), .B1(G898), .B2(new_n341), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(G69));
  AND3_X1   g736(.A1(new_n830), .A2(new_n674), .A3(new_n834), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n669), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT62), .Z(new_n925));
  NAND3_X1  g739(.A1(new_n667), .A2(new_n711), .A3(new_n800), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n738), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n740), .B2(new_n749), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n925), .A2(new_n756), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n274), .B(new_n519), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n341), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n650), .B2(G953), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n362), .A2(new_n704), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n749), .B1(new_n740), .B2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n756), .A2(new_n923), .A3(new_n798), .A4(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n932), .B1(new_n936), .B2(G953), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n412), .B2(new_n650), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G72));
  NAND2_X1  g754(.A1(G472), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT63), .Z(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n929), .B2(new_n845), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n872), .B1(new_n943), .B2(new_n662), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n935), .B2(new_n845), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n275), .B(KEYINPUT126), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n942), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n662), .A2(new_n275), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n839), .A2(new_n840), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n944), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT127), .ZN(G57));
endmodule


