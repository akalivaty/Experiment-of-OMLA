//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1316, new_n1317, new_n1318, new_n1319, new_n1321,
    new_n1322, new_n1323, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n208), .B1(new_n203), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G107), .ZN(new_n216));
  INV_X1    g0016(.A(G264), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n207), .B1(new_n212), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n207), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT0), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n220), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n202), .A2(new_n203), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT64), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT65), .Z(new_n232));
  AOI21_X1  g0032(.A(new_n225), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G58), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT82), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  AND3_X1   g0053(.A1(new_n253), .A2(KEYINPUT72), .A3(new_n226), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT72), .B1(new_n253), .B2(new_n226), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT8), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G58), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n261), .A2(new_n263), .B1(G150), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT73), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n265), .A2(new_n266), .B1(G20), .B2(new_n204), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  INV_X1    g0068(.A(new_n263), .ZN(new_n269));
  INV_X1    g0069(.A(G150), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n227), .A2(new_n262), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n268), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT73), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n257), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G13), .A3(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n253), .A2(new_n226), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT72), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n253), .A2(KEYINPUT72), .A3(new_n226), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n201), .B1(new_n275), .B2(G20), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n282), .A2(new_n283), .B1(new_n201), .B2(new_n277), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT9), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n274), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n204), .A2(G20), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n272), .B2(KEYINPUT73), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n265), .A2(new_n266), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n256), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(KEYINPUT9), .B1(new_n291), .B2(new_n284), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  AND2_X1   g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(KEYINPUT3), .A2(G33), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT70), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n262), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  NAND2_X1  g0100(.A1(KEYINPUT3), .A2(G33), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n294), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  XOR2_X1   g0103(.A(KEYINPUT71), .B(G223), .Z(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n297), .A2(new_n302), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G222), .A3(new_n294), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n297), .A2(new_n302), .A3(G77), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(G33), .A2(G41), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n226), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT68), .ZN(new_n313));
  OAI21_X1  g0113(.A(G274), .B1(new_n310), .B2(new_n226), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G274), .ZN(new_n317));
  AND2_X1   g0117(.A1(G1), .A2(G13), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G41), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n315), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(KEYINPUT68), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G226), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n315), .A2(KEYINPUT69), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n318), .A2(new_n319), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT69), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(new_n275), .C1(G41), .C2(G45), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n323), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n312), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT75), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(G200), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n330), .B1(new_n309), .B2(new_n311), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT75), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n312), .A2(G190), .A3(new_n331), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n293), .A2(new_n334), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n286), .B1(new_n274), .B2(new_n285), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n291), .A2(KEYINPUT9), .A3(new_n284), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT76), .A4(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT10), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n339), .B(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n275), .A2(G20), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n261), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n282), .A2(new_n347), .B1(new_n277), .B2(new_n268), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  INV_X1    g0149(.A(G159), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n271), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT79), .B1(new_n202), .B2(new_n203), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT79), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(G58), .A3(G68), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n354), .A3(new_n229), .ZN(new_n355));
  AOI211_X1 g0155(.A(new_n349), .B(new_n351), .C1(new_n355), .C2(G20), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT78), .B(G33), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n227), .B(new_n299), .C1(new_n357), .C2(new_n298), .ZN(new_n358));
  OAI21_X1  g0158(.A(G68), .B1(new_n358), .B2(KEYINPUT7), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n262), .A2(KEYINPUT78), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT78), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G33), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n296), .B1(new_n364), .B2(KEYINPUT3), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n360), .B1(new_n365), .B2(new_n227), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n356), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n256), .ZN(new_n368));
  NOR2_X1   g0168(.A1(KEYINPUT7), .A2(G20), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n297), .A2(new_n302), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n301), .A2(new_n227), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n357), .B2(new_n298), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n370), .B(G68), .C1(new_n372), .C2(new_n360), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n351), .B1(new_n355), .B2(G20), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT16), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n348), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT17), .ZN(new_n377));
  NOR2_X1   g0177(.A1(G223), .A2(G1698), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n324), .B2(G1698), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n298), .B1(new_n361), .B2(new_n363), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(new_n296), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G87), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n311), .ZN(new_n384));
  INV_X1    g0184(.A(new_n329), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(G232), .B1(new_n316), .B2(new_n322), .ZN(new_n386));
  INV_X1    g0186(.A(G190), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n387), .A2(KEYINPUT80), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(KEYINPUT80), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n384), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n314), .A2(new_n313), .A3(new_n315), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT68), .B1(new_n320), .B2(new_n321), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n393), .A2(new_n394), .B1(new_n329), .B2(new_n236), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n326), .B1(new_n381), .B2(new_n382), .ZN(new_n396));
  OAI21_X1  g0196(.A(G200), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n376), .A2(new_n377), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n348), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n365), .A2(new_n360), .A3(new_n227), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n358), .A2(KEYINPUT7), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n402), .A3(G68), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n257), .B1(new_n403), .B2(new_n356), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n373), .A2(new_n374), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n349), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n400), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n392), .A2(new_n397), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT17), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n399), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n384), .A2(new_n386), .A3(G179), .ZN(new_n411));
  OAI21_X1  g0211(.A(G169), .B1(new_n395), .B2(new_n396), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT18), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n412), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n376), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n410), .A2(KEYINPUT81), .A3(new_n414), .A4(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(G179), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n335), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n274), .A2(new_n285), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n420), .B(new_n422), .C1(G169), .C2(new_n335), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n377), .B1(new_n376), .B2(new_n398), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT17), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n424), .A2(new_n414), .A3(new_n417), .A4(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT81), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n345), .A2(new_n418), .A3(new_n423), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n236), .A2(G1698), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(G226), .B2(G1698), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n306), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G97), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n326), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n393), .A2(new_n394), .B1(new_n329), .B2(new_n209), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT13), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n385), .A2(G238), .B1(new_n316), .B2(new_n322), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT13), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n431), .B1(new_n302), .B2(new_n297), .ZN(new_n440));
  INV_X1    g0240(.A(new_n434), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n311), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G169), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT77), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT14), .ZN(new_n447));
  INV_X1    g0247(.A(G169), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n437), .B2(new_n443), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT14), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT77), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n450), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n437), .A2(G179), .A3(new_n443), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n447), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n264), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n269), .B2(new_n214), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n256), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n457), .A2(KEYINPUT11), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n277), .A2(new_n203), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT12), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n282), .A2(G68), .A3(new_n346), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(KEYINPUT11), .ZN(new_n462));
  AND4_X1   g0262(.A1(new_n458), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n454), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n387), .B2(new_n444), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n336), .B1(new_n437), .B2(new_n443), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n282), .A2(G77), .A3(new_n346), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n268), .A2(new_n271), .B1(new_n227), .B2(new_n214), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT15), .B(G87), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(new_n269), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n256), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n277), .A2(new_n214), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n470), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n323), .B1(new_n215), .B2(new_n329), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n303), .A2(G238), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n216), .B2(new_n306), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n306), .A2(G232), .A3(new_n294), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT74), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n306), .A2(KEYINPUT74), .A3(G232), .A4(new_n294), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n479), .B1(new_n486), .B2(new_n326), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n477), .B1(new_n487), .B2(new_n448), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n484), .A2(new_n485), .ZN(new_n489));
  INV_X1    g0289(.A(new_n306), .ZN(new_n490));
  AOI22_X1  g0290(.A1(G107), .A2(new_n490), .B1(new_n303), .B2(G238), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n478), .B1(new_n492), .B2(new_n311), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n419), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n476), .B1(new_n493), .B2(G190), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n487), .A2(G200), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n488), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n465), .A2(new_n469), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n252), .B1(new_n429), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n465), .A2(new_n469), .A3(new_n497), .ZN(new_n500));
  XNOR2_X1  g0300(.A(new_n426), .B(KEYINPUT81), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n293), .A2(new_n338), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(new_n344), .A3(new_n334), .A4(new_n337), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n339), .A2(new_n343), .A3(new_n342), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n503), .A2(new_n504), .A3(new_n423), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT82), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G250), .A2(G1698), .ZN(new_n508));
  INV_X1    g0308(.A(G257), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(G1698), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G294), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n365), .A2(new_n511), .B1(new_n512), .B2(new_n357), .ZN(new_n513));
  INV_X1    g0313(.A(G45), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G1), .ZN(new_n515));
  XNOR2_X1  g0315(.A(KEYINPUT5), .B(G41), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n311), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n513), .A2(new_n311), .B1(G264), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n320), .A2(new_n515), .A3(new_n516), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(G179), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n517), .A2(G264), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n299), .B1(new_n357), .B2(new_n298), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(new_n510), .B1(G294), .B2(new_n364), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n519), .C1(new_n523), .C2(new_n326), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G169), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT89), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n526), .B1(new_n520), .B2(new_n525), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT88), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n227), .B(G87), .C1(new_n380), .C2(new_n296), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n210), .A2(KEYINPUT22), .A3(G20), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(KEYINPUT22), .B1(new_n306), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G116), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n357), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n227), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n216), .A2(G20), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n531), .B(new_n532), .C1(new_n535), .C2(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n543), .A2(new_n256), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n533), .A2(KEYINPUT22), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n306), .A2(new_n534), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n547), .A2(KEYINPUT88), .A3(new_n538), .A4(new_n541), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n531), .B1(new_n535), .B2(new_n542), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT24), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n277), .A2(new_n216), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT25), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n275), .A2(G33), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n276), .B(new_n554), .C1(new_n254), .C2(new_n255), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n216), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n524), .B2(new_n387), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n336), .B1(new_n518), .B2(new_n519), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n530), .A2(new_n558), .B1(new_n551), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n253), .A2(new_n226), .B1(G20), .B2(new_n536), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G283), .ZN(new_n564));
  INV_X1    g0364(.A(G97), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n227), .C1(G33), .C2(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n563), .A2(KEYINPUT20), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT20), .B1(new_n563), .B2(new_n566), .ZN(new_n568));
  OAI22_X1  g0368(.A1(new_n567), .A2(new_n568), .B1(G116), .B2(new_n276), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n555), .A2(new_n536), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n448), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G257), .A2(G1698), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n217), .B2(G1698), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n380), .B2(new_n296), .ZN(new_n577));
  XNOR2_X1  g0377(.A(KEYINPUT86), .B(G303), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n297), .A2(new_n302), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n311), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n516), .A2(new_n515), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(G270), .A3(new_n326), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n583), .A2(new_n519), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n574), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n326), .B1(new_n577), .B2(new_n579), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n519), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n586), .A2(new_n587), .A3(new_n419), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n571), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n569), .A2(new_n570), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n581), .A2(G179), .A3(new_n584), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n573), .B1(new_n586), .B2(new_n587), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT87), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(G169), .B1(new_n586), .B2(new_n587), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n572), .B1(new_n598), .B2(new_n592), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n586), .A2(new_n587), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n571), .B1(new_n600), .B2(new_n391), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n336), .B2(new_n600), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n597), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n294), .A2(KEYINPUT4), .A3(G244), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n211), .B2(new_n294), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT70), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n564), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n215), .A2(G1698), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT4), .B1(new_n522), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n311), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n517), .A2(G257), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n519), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(G190), .A3(new_n615), .ZN(new_n616));
  OR3_X1    g0416(.A1(new_n276), .A2(KEYINPUT83), .A3(G97), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT83), .B1(new_n276), .B2(G97), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n555), .B2(new_n565), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n370), .B(G107), .C1(new_n372), .C2(new_n360), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n216), .A2(KEYINPUT6), .A3(G97), .ZN(new_n622));
  AND2_X1   g0422(.A1(G97), .A2(G107), .ZN(new_n623));
  NOR2_X1   g0423(.A1(G97), .A2(G107), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n622), .B1(new_n625), .B2(KEYINPUT6), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(G20), .B1(G77), .B2(new_n264), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n620), .B1(new_n628), .B2(new_n256), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n616), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT84), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n306), .A2(new_n605), .B1(G33), .B2(G283), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT4), .ZN(new_n633));
  INV_X1    g0433(.A(new_n610), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n633), .B1(new_n365), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n326), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n631), .B1(new_n636), .B2(new_n614), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n612), .A2(KEYINPUT84), .A3(new_n615), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(G200), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n630), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n612), .A2(new_n615), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n628), .A2(new_n256), .ZN(new_n642));
  INV_X1    g0442(.A(new_n620), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n641), .A2(new_n448), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n612), .A2(new_n419), .A3(new_n615), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n227), .B(G68), .C1(new_n380), .C2(new_n296), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT19), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n263), .A2(new_n649), .A3(G97), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n624), .A2(new_n210), .B1(new_n434), .B2(new_n227), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(new_n649), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n256), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n472), .A2(new_n277), .ZN(new_n655));
  INV_X1    g0455(.A(new_n555), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G87), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(G238), .A2(G1698), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n215), .B2(G1698), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n380), .B2(new_n296), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n364), .A2(G116), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n326), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n326), .B(G250), .C1(G1), .C2(new_n514), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n320), .A2(new_n515), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT85), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n666), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT85), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n537), .B1(new_n522), .B2(new_n660), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n668), .B(new_n669), .C1(new_n670), .C2(new_n326), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n658), .B1(new_n672), .B2(G190), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n667), .A2(new_n671), .A3(G200), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n419), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n654), .A2(new_n655), .ZN(new_n677));
  INV_X1    g0477(.A(new_n472), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n656), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n667), .A2(new_n671), .A3(new_n448), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n676), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n675), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n647), .A2(new_n683), .ZN(new_n684));
  AND4_X1   g0484(.A1(new_n507), .A2(new_n562), .A3(new_n603), .A4(new_n684), .ZN(G372));
  INV_X1    g0485(.A(new_n423), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n488), .A2(new_n494), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n687), .A2(new_n469), .B1(new_n454), .B2(new_n464), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n424), .A2(new_n425), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n414), .A2(new_n417), .A3(KEYINPUT93), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT93), .B1(new_n414), .B2(new_n417), .ZN(new_n691));
  OAI22_X1  g0491(.A1(new_n688), .A2(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n686), .B1(new_n692), .B2(new_n345), .ZN(new_n693));
  INV_X1    g0493(.A(new_n507), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n419), .A2(new_n672), .B1(new_n677), .B2(new_n679), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n663), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n670), .A2(KEYINPUT90), .A3(new_n326), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n668), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n448), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(G200), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n695), .A2(new_n700), .B1(new_n673), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT26), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n642), .A2(new_n643), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n448), .B1(new_n636), .B2(new_n614), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n704), .A2(new_n645), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n675), .A2(new_n682), .A3(new_n706), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT26), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n695), .A2(new_n700), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n520), .A2(new_n525), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n551), .B2(new_n557), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n448), .B1(new_n581), .B2(new_n584), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT21), .B1(new_n715), .B2(new_n571), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT91), .B1(new_n716), .B2(new_n595), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT91), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n589), .A2(new_n718), .A3(new_n599), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n639), .A2(new_n630), .B1(new_n644), .B2(new_n645), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT24), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n543), .A2(new_n256), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n561), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n702), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT92), .B1(new_n721), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n673), .A2(new_n701), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n725), .A2(new_n710), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT92), .ZN(new_n730));
  INV_X1    g0530(.A(new_n557), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n544), .B2(new_n550), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n719), .B(new_n717), .C1(new_n732), .C2(new_n713), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n729), .A2(new_n730), .A3(new_n733), .A4(new_n722), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n711), .B1(new_n727), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n693), .B1(new_n694), .B2(new_n735), .ZN(G369));
  INV_X1    g0536(.A(G13), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G1), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n227), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT27), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT27), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(new_n741), .A3(new_n227), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n740), .A2(G213), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G343), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT94), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n592), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT95), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n717), .A2(new_n719), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n603), .A2(new_n747), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT96), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n745), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n558), .A2(new_n530), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n712), .A2(KEYINPUT89), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n527), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n725), .B1(new_n757), .B2(new_n732), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n732), .A2(new_n745), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n753), .A2(G330), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n716), .B1(new_n591), .B2(new_n596), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n758), .A2(new_n762), .A3(new_n754), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n732), .A2(new_n713), .A3(new_n754), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n761), .A2(new_n765), .ZN(G399));
  INV_X1    g0566(.A(new_n222), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G41), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n624), .A2(new_n210), .A3(new_n536), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n769), .A2(G1), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n231), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n773), .B2(new_n769), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT97), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT28), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n562), .A2(new_n684), .A3(new_n603), .A4(new_n745), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT99), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n636), .A2(new_n614), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n672), .A2(new_n779), .A3(new_n518), .A4(new_n588), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT30), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND4_X1   g0582(.A1(new_n518), .A2(new_n588), .A3(new_n612), .A4(new_n615), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n783), .A2(KEYINPUT99), .A3(KEYINPUT30), .A4(new_n672), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n780), .A2(new_n781), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n600), .A2(G179), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n699), .A2(new_n524), .A3(new_n786), .A4(new_n641), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n782), .A2(new_n784), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n754), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT31), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT98), .B(KEYINPUT31), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n788), .A2(new_n754), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n777), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n795), .A2(G330), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT29), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n735), .B2(new_n754), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n762), .B1(new_n732), .B2(new_n757), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n647), .A2(KEYINPUT100), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT100), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n722), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n729), .A2(new_n799), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n710), .B1(new_n708), .B2(KEYINPUT26), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n703), .B1(new_n702), .B2(new_n706), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n754), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(KEYINPUT29), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n796), .B1(new_n798), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n776), .B1(new_n809), .B2(G1), .ZN(G364));
  NOR2_X1   g0610(.A1(new_n737), .A2(G20), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n275), .B1(new_n811), .B2(G45), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n768), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n753), .B2(G330), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(G330), .B2(new_n753), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n306), .A2(new_n222), .ZN(new_n817));
  INV_X1    g0617(.A(G355), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n817), .A2(new_n818), .B1(G116), .B2(new_n222), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n250), .A2(new_n514), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n232), .B2(new_n514), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n365), .A2(new_n222), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT101), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n819), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G13), .A2(G33), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(G20), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n226), .B1(G20), .B2(new_n448), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n814), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n227), .A2(new_n419), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(G200), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n390), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n336), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(G190), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n834), .A2(G50), .B1(new_n836), .B2(G77), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n390), .A2(new_n835), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n837), .B1(new_n202), .B2(new_n839), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT102), .Z(new_n841));
  NOR2_X1   g0641(.A1(new_n227), .A2(G179), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(G190), .A3(G200), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G87), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n842), .A2(new_n387), .A3(new_n336), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(G159), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n833), .A2(G190), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n845), .B1(new_n848), .B2(KEYINPUT32), .C1(new_n203), .C2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n842), .A2(new_n387), .A3(G200), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n848), .A2(KEYINPUT32), .B1(G107), .B2(new_n853), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n387), .A2(G179), .A3(G200), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n227), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n854), .B(new_n306), .C1(new_n565), .C2(new_n856), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n841), .A2(new_n851), .A3(new_n857), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n858), .A2(KEYINPUT103), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(KEYINPUT103), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n838), .A2(G322), .B1(new_n836), .B2(G311), .ZN(new_n861));
  INV_X1    g0661(.A(G283), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(new_n862), .B2(new_n852), .ZN(new_n863));
  INV_X1    g0663(.A(new_n856), .ZN(new_n864));
  XNOR2_X1  g0664(.A(KEYINPUT33), .B(G317), .ZN(new_n865));
  AOI22_X1  g0665(.A1(G294), .A2(new_n864), .B1(new_n849), .B2(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n834), .A2(G326), .B1(G303), .B2(new_n844), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n306), .B1(G329), .B2(new_n847), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n859), .B(new_n860), .C1(new_n863), .C2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n831), .B1(new_n870), .B2(new_n828), .ZN(new_n871));
  INV_X1    g0671(.A(new_n827), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n751), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n816), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(G396));
  NAND2_X1  g0675(.A1(new_n497), .A2(new_n745), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n735), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n488), .A2(new_n494), .A3(new_n745), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n495), .A2(new_n496), .B1(new_n476), .B2(new_n754), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(new_n687), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n735), .B2(new_n754), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n796), .ZN(new_n883));
  INV_X1    g0683(.A(new_n814), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n795), .A2(G330), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n877), .A2(new_n885), .A3(new_n881), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT105), .ZN(new_n888));
  INV_X1    g0688(.A(new_n880), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(new_n826), .ZN(new_n890));
  INV_X1    g0690(.A(new_n836), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n891), .A2(new_n536), .B1(new_n852), .B2(new_n210), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(G303), .B2(new_n834), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n306), .B1(G311), .B2(new_n847), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n864), .A2(G97), .B1(new_n844), .B2(G107), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n838), .A2(G294), .B1(new_n849), .B2(G283), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n365), .B1(G132), .B2(new_n847), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n852), .A2(new_n203), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n202), .B2(new_n856), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(G50), .B2(new_n844), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n834), .A2(G137), .B1(new_n836), .B2(G159), .ZN(new_n903));
  INV_X1    g0703(.A(G143), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n903), .B1(new_n904), .B2(new_n839), .C1(new_n270), .C2(new_n850), .ZN(new_n905));
  XNOR2_X1  g0705(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n898), .B(new_n902), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n897), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n828), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n828), .A2(new_n825), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n910), .B1(G77), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n814), .B1(new_n890), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n887), .A2(new_n888), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n888), .B1(new_n887), .B2(new_n914), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(G384));
  OR2_X1    g0718(.A1(new_n626), .A2(KEYINPUT35), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n626), .A2(KEYINPUT35), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n919), .A2(G116), .A3(new_n228), .A4(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(KEYINPUT106), .B(KEYINPUT36), .Z(new_n922));
  XNOR2_X1  g0722(.A(new_n921), .B(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n231), .A2(G77), .A3(new_n354), .A4(new_n352), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n201), .A2(G68), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n275), .B(G13), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT107), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n410), .B1(new_n690), .B2(new_n691), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n376), .A2(new_n743), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n376), .A2(new_n416), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n407), .A2(new_n408), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n930), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT37), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT37), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n933), .A2(new_n930), .A3(new_n934), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT38), .B1(new_n932), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n743), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n403), .A2(new_n374), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n349), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n400), .B1(new_n943), .B2(new_n404), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n934), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n413), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT37), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n938), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n944), .A2(new_n941), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n426), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(KEYINPUT38), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n928), .B1(new_n940), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n789), .A2(new_n792), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n788), .A2(KEYINPUT31), .A3(new_n754), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n777), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n463), .A2(new_n745), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n465), .A2(new_n469), .A3(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n464), .B(new_n754), .C1(new_n454), .C2(new_n468), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n880), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n956), .A2(new_n961), .A3(KEYINPUT40), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT93), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n407), .A2(new_n413), .A3(KEYINPUT18), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n415), .B1(new_n376), .B2(new_n416), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n414), .A2(new_n417), .A3(KEYINPUT93), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n689), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n939), .B1(new_n968), .B2(new_n930), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT38), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(KEYINPUT107), .A3(new_n951), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n953), .A2(new_n962), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(KEYINPUT38), .B1(new_n948), .B2(new_n950), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n956), .B(new_n961), .C1(new_n952), .C2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n973), .B1(KEYINPUT40), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n507), .A2(new_n956), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n978), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(G330), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT39), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n940), .B2(new_n952), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n465), .A2(new_n754), .ZN(new_n984));
  INV_X1    g0784(.A(new_n974), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n985), .A2(new_n951), .A3(KEYINPUT39), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n878), .B1(new_n735), .B2(new_n876), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n951), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n959), .A2(new_n960), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n966), .A2(new_n967), .A3(new_n941), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n987), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n507), .A2(new_n798), .A3(new_n808), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n693), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n993), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n981), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n275), .B2(new_n811), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n981), .A2(new_n996), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n927), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT108), .ZN(G367));
  AOI22_X1  g0801(.A1(new_n838), .A2(new_n578), .B1(new_n864), .B2(G107), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n847), .A2(G317), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(new_n365), .A3(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n834), .A2(G311), .B1(new_n836), .B2(G283), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n853), .A2(G97), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(new_n512), .C2(new_n850), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT46), .B1(new_n843), .B2(new_n536), .ZN(new_n1008));
  OR3_X1    g0808(.A1(new_n843), .A2(KEYINPUT46), .A3(new_n536), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1004), .B(new_n1007), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n849), .A2(G159), .B1(new_n844), .B2(G58), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n201), .B2(new_n891), .C1(new_n270), .C2(new_n839), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n856), .A2(new_n203), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G77), .B2(new_n853), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n834), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1014), .B1(new_n904), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(G137), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n306), .B1(new_n1017), .B2(new_n846), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1012), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1010), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT47), .Z(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n828), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n823), .A2(new_n242), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n830), .B1(new_n767), .B2(new_n678), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n884), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n754), .A2(new_n658), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n702), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n710), .B2(new_n1026), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1022), .B(new_n1025), .C1(new_n872), .C2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n754), .A2(new_n704), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n800), .A2(new_n802), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n706), .A2(new_n754), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n763), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT42), .Z(new_n1035));
  NOR3_X1   g0835(.A1(new_n1031), .A2(new_n732), .A3(new_n757), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n745), .B1(new_n1036), .B2(new_n706), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1028), .B(KEYINPUT43), .Z(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(KEYINPUT109), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1028), .A2(KEYINPUT43), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1035), .A2(new_n1037), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT109), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1038), .A2(new_n1044), .A3(new_n1039), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1041), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1046), .B1(new_n761), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n761), .A2(new_n1047), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1041), .A2(new_n1049), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n761), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n765), .A2(new_n1033), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT45), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n765), .A2(KEYINPUT45), .A3(new_n1033), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1047), .B(KEYINPUT44), .C1(new_n764), .C2(new_n763), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT44), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n765), .B2(new_n1033), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1057), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT110), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1052), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n753), .A2(G330), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n763), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n755), .B1(new_n762), .B2(new_n754), .C1(new_n758), .C2(new_n759), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n753), .A2(G330), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1055), .A2(new_n1056), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1072));
  OAI21_X1  g0872(.A(KEYINPUT110), .B1(new_n1072), .B2(new_n761), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1064), .A2(new_n1071), .A3(new_n809), .A4(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n761), .A3(KEYINPUT111), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(KEYINPUT111), .B1(new_n1072), .B2(new_n761), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n809), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n768), .B(KEYINPUT41), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n813), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1029), .B1(new_n1051), .B2(new_n1081), .ZN(G387));
  NAND2_X1  g0882(.A1(new_n1071), .A2(new_n813), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(KEYINPUT112), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(KEYINPUT112), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n760), .A2(new_n872), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n823), .B1(new_n239), .B2(new_n514), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n771), .B2(new_n817), .ZN(new_n1088));
  OR3_X1    g0888(.A1(new_n268), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1089));
  OAI21_X1  g0889(.A(KEYINPUT50), .B1(new_n268), .B2(G50), .ZN(new_n1090));
  AOI21_X1  g0890(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1089), .A2(new_n771), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1088), .A2(new_n1092), .B1(new_n216), .B2(new_n767), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n814), .B1(new_n1093), .B2(new_n830), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT113), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n838), .A2(G317), .B1(new_n836), .B2(new_n578), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1097), .A2(KEYINPUT115), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(KEYINPUT115), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n834), .A2(G322), .B1(new_n849), .B2(G311), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT48), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n864), .A2(G283), .B1(new_n844), .B2(G294), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT49), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n852), .A2(new_n536), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n522), .B(new_n1110), .C1(G326), .C2(new_n847), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1108), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n838), .A2(G50), .B1(new_n836), .B2(G68), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n268), .B2(new_n850), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n834), .A2(G159), .B1(G77), .B2(new_n844), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n864), .A2(new_n678), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n1006), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n522), .B1(new_n270), .B2(new_n846), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1114), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT114), .Z(new_n1120));
  NAND2_X1  g0920(.A1(new_n1112), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1095), .B1(new_n1121), .B2(new_n828), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1084), .A2(new_n1085), .B1(new_n1086), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n769), .B1(new_n1071), .B2(new_n809), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n809), .B2(new_n1071), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1125), .ZN(G393));
  INV_X1    g0926(.A(KEYINPUT116), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1052), .A2(new_n1062), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1072), .A2(new_n761), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT111), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(KEYINPUT116), .A3(new_n1075), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1128), .A2(new_n1129), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1071), .A2(new_n809), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n768), .A3(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1128), .A2(new_n1133), .A3(new_n813), .A4(new_n1129), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1047), .A2(new_n827), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT117), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G311), .A2(new_n838), .B1(new_n834), .B2(G317), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT52), .Z(new_n1143));
  OAI22_X1  g0943(.A1(new_n891), .A2(new_n512), .B1(new_n852), .B2(new_n216), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n306), .B(new_n1144), .C1(G322), .C2(new_n847), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n844), .A2(G283), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G116), .A2(new_n864), .B1(new_n849), .B2(new_n578), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G150), .A2(new_n834), .B1(new_n838), .B2(G159), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT51), .Z(new_n1150));
  NOR2_X1   g0950(.A1(new_n843), .A2(new_n203), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n856), .A2(new_n214), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(new_n261), .C2(new_n836), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n850), .A2(new_n201), .B1(new_n210), .B2(new_n852), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n365), .B(new_n1154), .C1(G143), .C2(new_n847), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1150), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1148), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n828), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n823), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n829), .B1(new_n565), .B2(new_n222), .C1(new_n1159), .C2(new_n247), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1141), .A2(new_n814), .A3(new_n1158), .A4(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1139), .A2(KEYINPUT118), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT118), .B1(new_n1139), .B2(new_n1161), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1138), .B1(new_n1163), .B2(new_n1164), .ZN(G390));
  NAND3_X1  g0965(.A1(new_n956), .A2(new_n961), .A3(G330), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n984), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n878), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n687), .A2(new_n879), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1169), .B1(new_n807), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n990), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1168), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n953), .A2(new_n972), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n988), .A2(new_n990), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1177), .A2(new_n1168), .B1(new_n983), .B2(new_n986), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1167), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n754), .B(new_n1170), .C1(new_n803), .C2(new_n806), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n990), .B1(new_n1180), .B2(new_n1169), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1181), .A2(new_n1168), .A3(new_n953), .A4(new_n972), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n796), .A2(new_n889), .A3(new_n990), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n983), .A2(new_n986), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n984), .B1(new_n988), .B2(new_n990), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1182), .B(new_n1183), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n990), .B1(new_n796), .B2(new_n889), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n988), .B1(new_n1188), .B2(new_n1167), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n956), .A2(G330), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1173), .B1(new_n1190), .B2(new_n880), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1183), .A2(new_n1172), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n956), .A2(G330), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n507), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n994), .A2(new_n693), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n769), .B1(new_n1187), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1196), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n1179), .A3(new_n1186), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1179), .A2(new_n1186), .A3(new_n813), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n814), .B1(new_n261), .B2(new_n912), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n490), .B1(G125), .B2(new_n847), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n838), .A2(G132), .B1(new_n849), .B2(G137), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(KEYINPUT54), .B(G143), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G159), .A2(new_n864), .B1(new_n836), .B2(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n834), .A2(G128), .B1(G50), .B2(new_n853), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1205), .A2(new_n1206), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n844), .A2(G150), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT53), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1152), .B1(G97), .B2(new_n836), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n306), .B1(G294), .B2(new_n847), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1214), .A2(new_n1215), .A3(new_n845), .A4(new_n900), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n838), .A2(G116), .B1(new_n849), .B2(G107), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n862), .B2(new_n1015), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1211), .A2(new_n1213), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1204), .B1(new_n1219), .B2(new_n828), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1184), .B2(new_n826), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1203), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1202), .A2(new_n1223), .ZN(G378));
  XNOR2_X1  g1024(.A(new_n1196), .B(KEYINPUT121), .ZN(new_n1225));
  INV_X1    g1025(.A(G330), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT40), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n975), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n973), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n422), .A2(new_n743), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT119), .Z(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  XOR2_X1   g1032(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n505), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n505), .A2(new_n1234), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1232), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1237), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(new_n1235), .A3(new_n1231), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1229), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n973), .A2(new_n1228), .A3(new_n1241), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n987), .A2(new_n991), .A3(new_n992), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n973), .A2(new_n1228), .A3(new_n1241), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1241), .B1(new_n973), .B2(new_n1228), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n993), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1201), .A2(new_n1225), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n768), .B1(new_n1250), .B2(KEYINPUT57), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1201), .A2(new_n1225), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1246), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1252), .A2(KEYINPUT57), .A3(new_n1253), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1251), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n813), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n884), .B1(new_n201), .B2(new_n911), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n828), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n834), .A2(G125), .B1(new_n836), .B2(G137), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n838), .A2(G128), .B1(new_n849), .B2(G132), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n864), .A2(G150), .B1(new_n844), .B2(new_n1208), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n853), .A2(G159), .ZN(new_n1265));
  AOI211_X1 g1065(.A(G33), .B(G41), .C1(new_n847), .C2(G124), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n891), .A2(new_n472), .B1(new_n214), .B2(new_n843), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1013), .B(new_n1268), .C1(G283), .C2(new_n847), .ZN(new_n1269));
  INV_X1    g1069(.A(G41), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n1015), .A2(new_n536), .B1(new_n202), .B2(new_n852), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n839), .A2(new_n216), .B1(new_n850), .B2(new_n565), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1269), .A2(new_n1270), .A3(new_n365), .A4(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1275), .A2(KEYINPUT58), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(KEYINPUT58), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G50), .B1(new_n262), .B2(new_n1270), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n522), .B2(G41), .ZN(new_n1279));
  AND4_X1   g1079(.A1(new_n1267), .A2(new_n1276), .A3(new_n1277), .A4(new_n1279), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1257), .B1(new_n1258), .B2(new_n1280), .C1(new_n1241), .C2(new_n826), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT120), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1256), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1255), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT122), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1255), .A2(KEYINPUT122), .A3(new_n1283), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1287), .A2(new_n1289), .ZN(G375));
  NAND2_X1  g1090(.A1(new_n1193), .A2(new_n813), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1173), .A2(new_n825), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(KEYINPUT123), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n884), .B1(new_n203), .B2(new_n911), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1116), .B1(new_n839), .B2(new_n862), .ZN(new_n1295));
  XOR2_X1   g1095(.A(new_n1295), .B(KEYINPUT124), .Z(new_n1296));
  AOI22_X1  g1096(.A1(new_n834), .A2(G294), .B1(new_n849), .B2(G116), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n844), .A2(G97), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n306), .B1(G303), .B2(new_n847), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n836), .A2(G107), .B1(new_n853), .B2(G77), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(new_n834), .A2(G132), .B1(G159), .B2(new_n844), .ZN(new_n1303));
  OAI221_X1 g1103(.A(new_n1303), .B1(new_n202), .B2(new_n852), .C1(new_n1017), .C2(new_n839), .ZN(new_n1304));
  AOI211_X1 g1104(.A(new_n365), .B(new_n1304), .C1(G128), .C2(new_n847), .ZN(new_n1305));
  OAI22_X1  g1105(.A1(new_n891), .A2(new_n270), .B1(new_n856), .B2(new_n201), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n849), .B2(new_n1208), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1302), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1293), .B(new_n1294), .C1(new_n1258), .C2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1291), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1198), .A2(new_n1080), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1189), .A2(new_n1196), .A3(new_n1192), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1310), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(G381));
  NOR2_X1   g1115(.A1(G393), .A2(G396), .ZN(new_n1316));
  INV_X1    g1116(.A(G384), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(new_n1314), .ZN(new_n1318));
  NOR4_X1   g1118(.A1(new_n1318), .A2(G387), .A3(G390), .A4(G378), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n1287), .B2(new_n1289), .ZN(G407));
  AOI21_X1  g1120(.A(G378), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1321));
  INV_X1    g1121(.A(G343), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(G213), .A3(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1124(.A(new_n1081), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(G390), .A2(new_n1327), .A3(new_n1029), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1164), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1162), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(G387), .A3(new_n1138), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n874), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1316), .A2(new_n1332), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1328), .A2(new_n1331), .A3(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1333), .B1(new_n1328), .B2(new_n1331), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  OAI211_X1 g1136(.A(G378), .B(new_n1283), .C1(new_n1251), .C2(new_n1254), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1247), .A2(new_n1248), .A3(new_n993), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1245), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1339));
  OAI21_X1  g1139(.A(KEYINPUT125), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT125), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1249), .A2(new_n1246), .A3(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1340), .A2(new_n813), .A3(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1252), .A2(new_n1080), .A3(new_n1253), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1344), .A3(new_n1282), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1222), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1337), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1322), .A2(G213), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1310), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1198), .A2(KEYINPUT60), .ZN(new_n1352));
  AND2_X1   g1152(.A1(new_n1352), .A2(new_n1313), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1189), .A2(new_n1196), .A3(KEYINPUT60), .A4(new_n1192), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(new_n768), .ZN(new_n1355));
  OAI211_X1 g1155(.A(G384), .B(new_n1351), .C1(new_n1353), .C2(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1355), .B1(new_n1352), .B2(new_n1313), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1317), .B1(new_n1357), .B2(new_n1310), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1322), .A2(G213), .A3(G2897), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1356), .A2(new_n1358), .A3(new_n1359), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1359), .B1(new_n1356), .B2(new_n1358), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(KEYINPUT61), .B1(new_n1350), .B2(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1356), .A2(new_n1358), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1364), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1348), .A2(new_n1349), .A3(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT63), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1366), .A2(new_n1367), .ZN(new_n1368));
  AOI22_X1  g1168(.A1(new_n1337), .A2(new_n1347), .B1(G213), .B2(new_n1322), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1369), .A2(KEYINPUT63), .A3(new_n1365), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1336), .A2(new_n1363), .A3(new_n1368), .A4(new_n1370), .ZN(new_n1371));
  AND4_X1   g1171(.A1(KEYINPUT62), .A2(new_n1348), .A3(new_n1349), .A4(new_n1365), .ZN(new_n1372));
  AOI21_X1  g1172(.A(KEYINPUT62), .B1(new_n1369), .B2(new_n1365), .ZN(new_n1373));
  OAI211_X1 g1173(.A(new_n1363), .B(KEYINPUT126), .C1(new_n1372), .C2(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1336), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1374), .A2(new_n1375), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT62), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1366), .A2(new_n1377), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1369), .A2(KEYINPUT62), .A3(new_n1365), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1378), .A2(new_n1379), .ZN(new_n1380));
  AOI21_X1  g1180(.A(KEYINPUT126), .B1(new_n1380), .B2(new_n1363), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1371), .B1(new_n1376), .B2(new_n1381), .ZN(G405));
  OAI21_X1  g1182(.A(new_n1364), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1328), .A2(new_n1331), .ZN(new_n1384));
  INV_X1    g1184(.A(new_n1333), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1384), .A2(new_n1385), .ZN(new_n1386));
  NAND3_X1  g1186(.A1(new_n1328), .A2(new_n1331), .A3(new_n1333), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n1386), .A2(new_n1365), .A3(new_n1387), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1383), .A2(new_n1388), .ZN(new_n1389));
  AOI21_X1  g1189(.A(new_n1346), .B1(new_n1255), .B2(new_n1283), .ZN(new_n1390));
  NOR2_X1   g1190(.A1(new_n1321), .A2(new_n1390), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1389), .A2(new_n1391), .ZN(new_n1392));
  OAI211_X1 g1192(.A(new_n1383), .B(new_n1388), .C1(new_n1321), .C2(new_n1390), .ZN(new_n1393));
  AND2_X1   g1193(.A1(new_n1392), .A2(new_n1393), .ZN(G402));
endmodule


