//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1086, new_n1087;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G127gat), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G134gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT68), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G113gat), .ZN(new_n210));
  INV_X1    g009(.A(G113gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G120gat), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT1), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n206), .A2(G134gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n204), .A2(G127gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n208), .A2(new_n213), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT67), .ZN(new_n219));
  OR3_X1    g018(.A1(new_n204), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G113gat), .B(G120gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n219), .B(new_n220), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(KEYINPUT23), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227));
  NOR3_X1   g026(.A1(new_n227), .A2(G169gat), .A3(G176gat), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n226), .A2(KEYINPUT25), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(KEYINPUT64), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT64), .B1(new_n232), .B2(new_n233), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n229), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n228), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n231), .A2(KEYINPUT65), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G183gat), .ZN(new_n243));
  INV_X1    g042(.A(G190gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n231), .B1(KEYINPUT65), .B2(new_n241), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n239), .B(new_n240), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n237), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT26), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n224), .B1(new_n251), .B2(new_n225), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n251), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n231), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT28), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT27), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G183gat), .ZN(new_n258));
  AOI21_X1  g057(.A(G190gat), .B1(new_n258), .B2(KEYINPUT66), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n243), .A2(KEYINPUT27), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT66), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n256), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n261), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n264), .A2(new_n256), .A3(G190gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n255), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n223), .B1(new_n250), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n232), .A2(new_n233), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n234), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n272), .A2(new_n229), .B1(KEYINPUT25), .B2(new_n248), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n218), .A2(new_n222), .ZN(new_n274));
  INV_X1    g073(.A(new_n252), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n275), .A2(new_n253), .B1(G183gat), .B2(G190gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n264), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT28), .B1(new_n278), .B2(new_n259), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n276), .B1(new_n279), .B2(new_n265), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n273), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n268), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT32), .ZN(new_n286));
  XOR2_X1   g085(.A(G15gat), .B(G43gat), .Z(new_n287));
  XNOR2_X1  g086(.A(G71gat), .B(G99gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n290));
  AOI21_X1  g089(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n284), .A2(new_n285), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n285), .B1(new_n284), .B2(new_n291), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n286), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n284), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n289), .ZN(new_n297));
  OAI22_X1  g096(.A1(new_n293), .A2(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n250), .A2(new_n267), .A3(new_n223), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n274), .B1(new_n273), .B2(new_n280), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n282), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n283), .B1(new_n268), .B2(new_n281), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT34), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n203), .B1(new_n298), .B2(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n302), .A2(new_n306), .A3(new_n307), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n297), .B1(new_n284), .B2(new_n295), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n284), .A2(new_n291), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT70), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n313), .B2(new_n292), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n314), .A3(KEYINPUT72), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n309), .A2(new_n315), .B1(new_n298), .B2(new_n308), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n202), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n298), .A2(new_n308), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n298), .A2(new_n308), .A3(new_n203), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT72), .B1(new_n310), .B2(new_n314), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(KEYINPUT73), .A3(KEYINPUT36), .ZN(new_n323));
  XNOR2_X1  g122(.A(G8gat), .B(G36gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(G64gat), .B(G92gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT22), .ZN(new_n328));
  INV_X1    g127(.A(G211gat), .ZN(new_n329));
  INV_X1    g128(.A(G218gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G211gat), .B(G218gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n332), .B(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n336), .B(KEYINPUT74), .Z(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT75), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n250), .A2(new_n267), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n280), .A2(new_n249), .A3(new_n237), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n337), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n335), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n337), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n335), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n338), .B1(new_n273), .B2(new_n280), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n326), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n347), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n339), .A2(KEYINPUT29), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n335), .B(new_n350), .C1(new_n351), .C2(new_n337), .ZN(new_n352));
  INV_X1    g151(.A(new_n342), .ZN(new_n353));
  INV_X1    g152(.A(new_n338), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(new_n341), .B2(new_n344), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n346), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n326), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n349), .A2(KEYINPUT30), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n348), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT30), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(new_n357), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT2), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT78), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(new_n367), .A3(KEYINPUT2), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n370));
  INV_X1    g169(.A(G141gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n371), .A3(G148gat), .ZN(new_n372));
  INV_X1    g171(.A(G148gat), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT77), .B1(new_n373), .B2(G141gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(G141gat), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G155gat), .ZN(new_n377));
  INV_X1    g176(.A(G162gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n364), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n369), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT76), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(G155gat), .B2(G162gat), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n382), .A2(new_n384), .A3(new_n364), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT2), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n371), .A2(G148gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n386), .B1(new_n375), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n381), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n274), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n218), .A2(new_n222), .A3(KEYINPUT79), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n381), .A2(new_n395), .A3(new_n389), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n391), .A2(new_n393), .A3(new_n394), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n371), .A2(G148gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n398), .B1(new_n387), .B2(KEYINPUT77), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n399), .A2(new_n372), .B1(new_n364), .B2(new_n379), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n400), .A2(new_n369), .B1(new_n388), .B2(new_n385), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(new_n223), .A3(KEYINPUT4), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n390), .B2(new_n274), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT83), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(KEYINPUT5), .ZN(new_n411));
  AND4_X1   g210(.A1(new_n397), .A2(new_n406), .A3(new_n408), .A4(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n397), .A2(new_n404), .A3(new_n402), .A4(new_n409), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT80), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n381), .A2(new_n395), .A3(new_n389), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n395), .B1(new_n381), .B2(new_n389), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n218), .A2(new_n222), .A3(KEYINPUT79), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT79), .B1(new_n218), .B2(new_n222), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n410), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n402), .A2(new_n404), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT80), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n390), .A2(new_n274), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(KEYINPUT81), .A3(new_n390), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n393), .A2(new_n390), .A3(new_n394), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT5), .B1(new_n432), .B2(new_n409), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n413), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  XOR2_X1   g233(.A(G1gat), .B(G29gat), .Z(new_n435));
  XNOR2_X1  g234(.A(G57gat), .B(G85gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  NAND2_X1  g238(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT5), .ZN(new_n442));
  INV_X1    g241(.A(new_n427), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT81), .B1(new_n422), .B2(new_n390), .ZN(new_n444));
  AND4_X1   g243(.A1(KEYINPUT81), .A2(new_n393), .A3(new_n390), .A4(new_n394), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n442), .B1(new_n446), .B2(new_n410), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n414), .A2(new_n415), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n423), .A2(KEYINPUT80), .A3(new_n424), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n412), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n439), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n440), .A2(new_n441), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n434), .A2(KEYINPUT6), .A3(new_n439), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n363), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(KEYINPUT31), .B(G50gat), .Z(new_n457));
  NOR2_X1   g256(.A1(new_n332), .A2(new_n334), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n333), .B1(new_n331), .B2(new_n327), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n344), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n401), .B1(new_n395), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n335), .B1(new_n396), .B2(new_n344), .ZN(new_n462));
  INV_X1    g261(.A(G228gat), .ZN(new_n463));
  INV_X1    g262(.A(G233gat), .ZN(new_n464));
  OAI22_X1  g263(.A1(new_n461), .A2(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n396), .A2(new_n344), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT84), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n396), .A2(KEYINPUT84), .A3(new_n344), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n335), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT3), .B1(new_n335), .B2(new_n344), .ZN(new_n471));
  OAI211_X1 g270(.A(G228gat), .B(G233gat), .C1(new_n471), .C2(new_n401), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n465), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(G22gat), .ZN(new_n474));
  INV_X1    g273(.A(G22gat), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n475), .B(new_n465), .C1(new_n470), .C2(new_n472), .ZN(new_n476));
  XNOR2_X1  g275(.A(G78gat), .B(G106gat), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n474), .B2(new_n476), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n457), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n477), .ZN(new_n481));
  INV_X1    g280(.A(new_n472), .ZN(new_n482));
  INV_X1    g281(.A(new_n469), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT84), .B1(new_n396), .B2(new_n344), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n346), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n475), .B1(new_n486), .B2(new_n465), .ZN(new_n487));
  INV_X1    g286(.A(new_n476), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n481), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n490));
  INV_X1    g289(.A(new_n457), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n480), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n318), .B(new_n323), .C1(new_n456), .C2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT39), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n432), .B2(new_n409), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n406), .A2(new_n397), .A3(new_n408), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n410), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n497), .A3(new_n410), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n452), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT40), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n501), .A2(KEYINPUT40), .A3(new_n452), .A4(new_n502), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n363), .A2(new_n505), .A3(new_n440), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n455), .A2(KEYINPUT86), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n434), .A2(new_n509), .A3(KEYINPUT6), .A4(new_n439), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n454), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n358), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n352), .A2(new_n356), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT85), .B1(new_n513), .B2(KEYINPUT37), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT37), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n360), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n340), .A2(new_n342), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n516), .B1(new_n519), .B2(new_n335), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n346), .B(new_n350), .C1(new_n351), .C2(new_n337), .ZN(new_n521));
  AOI211_X1 g320(.A(KEYINPUT38), .B(new_n357), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n512), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n326), .B1(new_n360), .B2(new_n516), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(new_n514), .B2(new_n517), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n507), .B(new_n494), .C1(new_n511), .C2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n441), .B1(new_n451), .B2(new_n452), .ZN(new_n529));
  AOI211_X1 g328(.A(new_n439), .B(new_n412), .C1(new_n450), .C2(new_n447), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n455), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n363), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n309), .A2(new_n315), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(new_n480), .A3(new_n319), .A4(new_n492), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT35), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT87), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n322), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n316), .A2(KEYINPUT87), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT35), .B1(new_n359), .B2(new_n362), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n480), .A2(new_n540), .A3(new_n492), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n511), .A2(new_n538), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n496), .A2(new_n528), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  INV_X1    g344(.A(G1gat), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(KEYINPUT16), .A3(new_n546), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(G8gat), .ZN(new_n550));
  INV_X1    g349(.A(G8gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(new_n551), .A3(new_n548), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554));
  INV_X1    g353(.A(G43gat), .ZN(new_n555));
  INV_X1    g354(.A(G50gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G43gat), .A2(G50gat), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT14), .ZN(new_n560));
  INV_X1    g359(.A(G29gat), .ZN(new_n561));
  INV_X1    g360(.A(G36gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G29gat), .A2(G36gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n559), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  INV_X1    g370(.A(new_n559), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n563), .A2(new_n565), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n554), .A3(new_n558), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n567), .A4(new_n574), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n571), .B1(new_n570), .B2(new_n575), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n544), .B(new_n553), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n547), .A2(new_n551), .A3(new_n548), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n551), .B1(new_n547), .B2(new_n548), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT91), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT91), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n550), .A2(new_n582), .A3(new_n552), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n570), .A2(new_n575), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(KEYINPUT17), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n544), .B1(new_n589), .B2(new_n553), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n591), .A2(KEYINPUT92), .A3(KEYINPUT18), .A4(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT92), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n553), .B1(new_n576), .B2(new_n577), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT90), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n596), .A2(new_n592), .A3(new_n578), .A4(new_n585), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT18), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n592), .B(KEYINPUT13), .Z(new_n601));
  INV_X1    g400(.A(new_n585), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n584), .B1(new_n581), .B2(new_n583), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(KEYINPUT93), .B(new_n601), .C1(new_n602), .C2(new_n603), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n606), .A2(new_n607), .B1(new_n597), .B2(new_n598), .ZN(new_n608));
  XOR2_X1   g407(.A(G113gat), .B(G141gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT11), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT88), .ZN(new_n611));
  XNOR2_X1  g410(.A(G169gat), .B(G197gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n600), .A2(new_n608), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n614), .B1(new_n600), .B2(new_n608), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G183gat), .B(G211gat), .Z(new_n618));
  INV_X1    g417(.A(G231gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(new_n464), .ZN(new_n620));
  NAND2_X1  g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT9), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(G64gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(G57gat), .ZN(new_n625));
  INV_X1    g424(.A(G57gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(G64gat), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n623), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(G71gat), .A2(G78gat), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n629), .A2(new_n630), .A3(KEYINPUT94), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n632));
  OR2_X1    g431(.A1(G71gat), .A2(G78gat), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n632), .B1(new_n633), .B2(new_n621), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n628), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT95), .B1(new_n626), .B2(G64gat), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT95), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(new_n624), .A3(G57gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n626), .A2(G64gat), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n633), .A2(KEYINPUT96), .A3(new_n621), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT96), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n629), .B2(new_n630), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n640), .A2(new_n623), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n620), .B1(new_n645), .B2(KEYINPUT21), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n635), .A2(new_n644), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT21), .ZN(new_n648));
  INV_X1    g447(.A(new_n620), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G127gat), .B(G155gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n646), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n651), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n649), .B1(new_n647), .B2(new_n648), .ZN(new_n654));
  AOI211_X1 g453(.A(KEYINPUT21), .B(new_n620), .C1(new_n635), .C2(new_n644), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n652), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n652), .B2(new_n656), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n581), .A2(new_n583), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n645), .A2(KEYINPUT21), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n659), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n651), .B1(new_n646), .B2(new_n650), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n654), .A2(new_n655), .A3(new_n653), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n657), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n656), .A3(new_n658), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n663), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n618), .B1(new_n665), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n664), .B1(new_n659), .B2(new_n660), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n668), .A2(new_n663), .A3(new_n669), .ZN(new_n673));
  INV_X1    g472(.A(new_n618), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677));
  INV_X1    g476(.A(G232gat), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n464), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(KEYINPUT41), .ZN(new_n680));
  XNOR2_X1  g479(.A(G134gat), .B(G162gat), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n680), .B(new_n681), .Z(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(G190gat), .B(G218gat), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT98), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT7), .ZN(new_n686));
  AND3_X1   g485(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT99), .B1(G85gat), .B2(G92gat), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(G85gat), .A2(G92gat), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT99), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT7), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(KEYINPUT98), .ZN(new_n694));
  NAND3_X1  g493(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(G99gat), .A2(G106gat), .ZN(new_n697));
  INV_X1    g496(.A(G85gat), .ZN(new_n698));
  INV_X1    g497(.A(G92gat), .ZN(new_n699));
  AOI22_X1  g498(.A1(KEYINPUT8), .A2(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n689), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(G99gat), .A2(G106gat), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT100), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n703), .A3(new_n697), .ZN(new_n704));
  AND2_X1   g503(.A1(G99gat), .A2(G106gat), .ZN(new_n705));
  NOR2_X1   g504(.A1(G99gat), .A2(G106gat), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT100), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n701), .A2(new_n708), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT101), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n704), .A2(new_n707), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n712), .A2(new_n696), .A3(new_n689), .A4(new_n700), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n701), .A2(new_n708), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n587), .A2(new_n588), .B1(new_n711), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n713), .A2(new_n715), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n584), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n679), .A2(KEYINPUT41), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n684), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n716), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n714), .B1(new_n713), .B2(new_n715), .ZN(new_n724));
  OAI22_X1  g523(.A1(new_n723), .A2(new_n724), .B1(new_n576), .B2(new_n577), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n718), .A2(new_n584), .B1(KEYINPUT41), .B2(new_n679), .ZN(new_n726));
  INV_X1    g525(.A(new_n684), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n722), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT97), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n683), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI211_X1 g530(.A(KEYINPUT97), .B(new_n682), .C1(new_n722), .C2(new_n728), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n677), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n717), .A2(new_n721), .A3(new_n684), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n727), .B1(new_n725), .B2(new_n726), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n730), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n682), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n729), .A2(new_n677), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n729), .A2(new_n730), .A3(new_n683), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n676), .A2(new_n733), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(G230gat), .A2(G233gat), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n718), .A2(new_n645), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT10), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n713), .A2(new_n647), .A3(new_n715), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n718), .A2(KEYINPUT10), .A3(new_n645), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n743), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n744), .A2(new_n746), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(new_n743), .ZN(new_n751));
  XNOR2_X1  g550(.A(G120gat), .B(G148gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(G176gat), .B(G204gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  AOI211_X1 g555(.A(new_n754), .B(new_n749), .C1(new_n750), .C2(new_n743), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n543), .A2(new_n617), .A3(new_n741), .A4(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n531), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT103), .B(G1gat), .Z(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1324gat));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n363), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT42), .B1(new_n765), .B2(new_n551), .ZN(new_n766));
  OR2_X1    g565(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  MUX2_X1   g568(.A(KEYINPUT42), .B(new_n766), .S(new_n769), .Z(G1325gat));
  INV_X1    g569(.A(G15gat), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n534), .A2(KEYINPUT87), .A3(new_n319), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT87), .B1(new_n534), .B2(new_n319), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n316), .A2(new_n317), .A3(new_n202), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT36), .B1(new_n322), .B2(KEYINPUT73), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n759), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n780), .B2(new_n771), .ZN(G1326gat));
  NAND2_X1  g580(.A1(new_n759), .A2(new_n493), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT43), .B(G22gat), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1327gat));
  NAND2_X1  g583(.A1(new_n542), .A2(new_n536), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n494), .A2(new_n507), .ZN(new_n786));
  INV_X1    g585(.A(new_n527), .ZN(new_n787));
  INV_X1    g586(.A(new_n511), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n785), .B1(new_n789), .B2(new_n495), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n733), .A2(new_n740), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n617), .A2(new_n676), .A3(new_n758), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n561), .A3(new_n760), .ZN(new_n796));
  XOR2_X1   g595(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n799));
  XOR2_X1   g598(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n800));
  AND4_X1   g599(.A1(KEYINPUT106), .A2(new_n790), .A3(new_n791), .A4(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n733), .A2(new_n740), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n531), .A2(new_n532), .B1(new_n492), .B2(new_n480), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n528), .A2(new_n778), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n802), .B1(new_n805), .B2(new_n785), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n800), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT106), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n801), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n799), .B1(new_n810), .B2(new_n794), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT44), .B1(new_n543), .B2(new_n802), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n812), .A2(KEYINPUT106), .B1(new_n806), .B2(new_n800), .ZN(new_n813));
  OAI211_X1 g612(.A(KEYINPUT107), .B(new_n793), .C1(new_n813), .C2(new_n801), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n811), .A2(new_n760), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n798), .B1(new_n815), .B2(new_n561), .ZN(G1328gat));
  NAND3_X1  g615(.A1(new_n811), .A2(new_n363), .A3(new_n814), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT108), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT108), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n811), .A2(new_n814), .A3(new_n819), .A4(new_n363), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(G36gat), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n795), .A2(new_n562), .A3(new_n363), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT46), .Z(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1329gat));
  INV_X1    g623(.A(new_n774), .ZN(new_n825));
  NOR4_X1   g624(.A1(new_n792), .A2(G43gat), .A3(new_n825), .A4(new_n794), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n810), .A2(new_n778), .A3(new_n794), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(new_n555), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n811), .A2(new_n779), .A3(new_n814), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n826), .B1(new_n831), .B2(G43gat), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n832), .B2(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g632(.A(new_n808), .B1(new_n790), .B2(new_n791), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT106), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n807), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n801), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n794), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n556), .B1(new_n838), .B2(new_n493), .ZN(new_n839));
  NOR4_X1   g638(.A1(new_n792), .A2(G50gat), .A3(new_n494), .A4(new_n794), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT48), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT109), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT109), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n810), .A2(new_n494), .A3(new_n794), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n845), .B(new_n842), .C1(new_n846), .C2(new_n556), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n811), .A2(new_n493), .A3(new_n814), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n840), .B1(new_n849), .B2(G50gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n850), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g650(.A1(new_n741), .A2(new_n616), .A3(new_n615), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n790), .A2(new_n758), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n760), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n363), .ZN(new_n856));
  NOR2_X1   g655(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n857));
  AND2_X1   g656(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n859), .B1(new_n857), .B2(new_n856), .ZN(G1333gat));
  NAND2_X1  g659(.A1(new_n853), .A2(new_n779), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT110), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n772), .B2(new_n773), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT110), .ZN(new_n864));
  AOI21_X1  g663(.A(G71gat), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n861), .A2(G71gat), .B1(new_n853), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g666(.A1(new_n853), .A2(new_n493), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g668(.A1(new_n600), .A2(new_n608), .ZN(new_n870));
  INV_X1    g669(.A(new_n614), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n600), .A2(new_n608), .A3(new_n614), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n676), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n758), .B(new_n875), .C1(new_n813), .C2(new_n801), .ZN(new_n876));
  OAI21_X1  g675(.A(G85gat), .B1(new_n876), .B2(new_n531), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT111), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n792), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n806), .A2(KEYINPUT111), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT51), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT51), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n879), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n760), .A2(new_n698), .A3(new_n758), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n877), .B1(new_n886), .B2(new_n887), .ZN(G1336gat));
  NAND3_X1  g687(.A1(new_n363), .A2(new_n758), .A3(new_n699), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT113), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(new_n883), .B2(new_n885), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n532), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n699), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT112), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  OAI221_X1 g696(.A(new_n891), .B1(new_n895), .B2(new_n894), .C1(new_n892), .C2(new_n699), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1337gat));
  OAI21_X1  g698(.A(G99gat), .B1(new_n876), .B2(new_n778), .ZN(new_n900));
  INV_X1    g699(.A(new_n758), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n825), .A2(G99gat), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n886), .B2(new_n902), .ZN(G1338gat));
  OAI21_X1  g702(.A(G106gat), .B1(new_n876), .B2(new_n494), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n494), .A2(G106gat), .A3(new_n901), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n905), .B1(new_n883), .B2(new_n885), .ZN(new_n906));
  XNOR2_X1  g705(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n904), .B2(new_n906), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(G1339gat));
  INV_X1    g709(.A(KEYINPUT115), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n911), .B1(new_n852), .B2(new_n901), .ZN(new_n912));
  NOR4_X1   g711(.A1(new_n874), .A2(new_n741), .A3(KEYINPUT115), .A4(new_n758), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n747), .A2(new_n748), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n742), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n747), .A2(new_n748), .A3(new_n743), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(KEYINPUT54), .A3(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n755), .B1(new_n749), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT55), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n751), .A2(new_n755), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n918), .A2(KEYINPUT55), .A3(new_n920), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n925), .B1(new_n872), .B2(new_n873), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n591), .A2(new_n592), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n602), .A2(new_n603), .A3(new_n601), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n613), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n758), .A2(new_n873), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n802), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n924), .A2(new_n923), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(new_n921), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n791), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n873), .A2(new_n929), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n676), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT116), .B1(new_n914), .B2(new_n937), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n617), .A2(new_n676), .A3(new_n802), .A4(new_n901), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT115), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n852), .A2(new_n911), .A3(new_n901), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n676), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n933), .B1(new_n615), .B2(new_n616), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n758), .A2(new_n873), .A3(new_n929), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n791), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n934), .A2(new_n935), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT116), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n942), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n938), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n760), .A2(new_n532), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n825), .A2(new_n493), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n955), .A2(new_n211), .A3(new_n617), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n951), .A2(new_n531), .A3(new_n535), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT117), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n532), .A3(new_n874), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n959), .B2(new_n211), .ZN(G1340gat));
  NOR3_X1   g759(.A1(new_n955), .A2(new_n209), .A3(new_n901), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n958), .A2(new_n532), .A3(new_n758), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n209), .ZN(G1341gat));
  NAND3_X1  g762(.A1(new_n958), .A2(new_n532), .A3(new_n676), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT118), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n943), .A2(new_n206), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n965), .B1(new_n955), .B2(new_n967), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n953), .A2(KEYINPUT118), .A3(new_n954), .A4(new_n966), .ZN(new_n969));
  AOI22_X1  g768(.A1(new_n964), .A2(new_n206), .B1(new_n968), .B2(new_n969), .ZN(G1342gat));
  OAI21_X1  g769(.A(G134gat), .B1(new_n955), .B2(new_n802), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n802), .A2(G134gat), .A3(new_n363), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n958), .A2(KEYINPUT56), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT56), .B1(new_n958), .B2(new_n972), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1343gat));
  NAND3_X1  g774(.A1(new_n778), .A2(new_n760), .A3(new_n532), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n918), .A2(new_n920), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT119), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT55), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n932), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(new_n874), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(new_n945), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n947), .B1(new_n982), .B2(new_n802), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n983), .A2(new_n676), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n493), .B1(new_n984), .B2(new_n914), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n976), .B1(new_n985), .B2(KEYINPUT57), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n942), .A2(new_n949), .A3(new_n948), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n949), .B1(new_n942), .B2(new_n948), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT57), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n989), .A2(new_n990), .A3(new_n493), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(G141gat), .B1(new_n992), .B2(new_n617), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT120), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n778), .A2(new_n493), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n951), .A2(new_n952), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n997), .A2(new_n371), .A3(new_n874), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n995), .A2(new_n999), .A3(KEYINPUT58), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT58), .ZN(new_n1001));
  OAI211_X1 g800(.A(new_n993), .B(new_n998), .C1(new_n994), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1000), .A2(new_n1002), .ZN(G1344gat));
  INV_X1    g802(.A(KEYINPUT59), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n1005));
  INV_X1    g804(.A(new_n939), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1005), .B1(new_n984), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g806(.A(KEYINPUT122), .B(new_n939), .C1(new_n983), .C2(new_n676), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n1007), .A2(new_n990), .A3(new_n493), .A4(new_n1008), .ZN(new_n1009));
  OAI21_X1  g808(.A(KEYINPUT57), .B1(new_n951), .B2(new_n494), .ZN(new_n1010));
  AND2_X1   g809(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g810(.A(new_n976), .B(KEYINPUT121), .Z(new_n1012));
  NAND3_X1  g811(.A1(new_n1011), .A2(new_n758), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n1004), .B1(new_n1013), .B2(G148gat), .ZN(new_n1014));
  INV_X1    g813(.A(new_n992), .ZN(new_n1015));
  AOI211_X1 g814(.A(KEYINPUT59), .B(new_n373), .C1(new_n1015), .C2(new_n758), .ZN(new_n1016));
  NAND4_X1  g815(.A1(new_n989), .A2(new_n760), .A3(new_n493), .A4(new_n778), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n532), .A2(new_n373), .A3(new_n758), .ZN(new_n1018));
  OAI22_X1  g817(.A1(new_n1014), .A2(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(G1345gat));
  AOI21_X1  g818(.A(G155gat), .B1(new_n997), .B2(new_n676), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n943), .A2(new_n377), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1020), .B1(new_n1015), .B2(new_n1021), .ZN(G1346gat));
  OAI21_X1  g821(.A(G162gat), .B1(new_n992), .B2(new_n802), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n791), .A2(new_n378), .A3(new_n532), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1023), .B1(new_n1017), .B2(new_n1024), .ZN(G1347gat));
  NAND2_X1  g824(.A1(new_n863), .A2(new_n864), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n531), .A2(new_n363), .ZN(new_n1027));
  INV_X1    g826(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g828(.A(KEYINPUT124), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g830(.A(new_n1027), .B1(new_n863), .B2(new_n864), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n493), .B1(new_n1032), .B2(KEYINPUT124), .ZN(new_n1033));
  NAND4_X1  g832(.A1(new_n938), .A2(new_n950), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  INV_X1    g833(.A(G169gat), .ZN(new_n1035));
  NOR3_X1   g834(.A1(new_n1034), .A2(new_n1035), .A3(new_n617), .ZN(new_n1036));
  NOR2_X1   g835(.A1(new_n951), .A2(new_n760), .ZN(new_n1037));
  NOR2_X1   g836(.A1(new_n535), .A2(new_n532), .ZN(new_n1038));
  XNOR2_X1  g837(.A(new_n1038), .B(KEYINPUT123), .ZN(new_n1039));
  NAND3_X1  g838(.A1(new_n1037), .A2(new_n874), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g839(.A(new_n1036), .B1(new_n1040), .B2(new_n1035), .ZN(G1348gat));
  OAI21_X1  g840(.A(G176gat), .B1(new_n1034), .B2(new_n901), .ZN(new_n1042));
  NAND2_X1  g841(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1043));
  OR2_X1    g842(.A1(new_n901), .A2(G176gat), .ZN(new_n1044));
  OAI21_X1  g843(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(G1349gat));
  OAI21_X1  g844(.A(G183gat), .B1(new_n1034), .B2(new_n943), .ZN(new_n1046));
  NOR2_X1   g845(.A1(new_n943), .A2(new_n264), .ZN(new_n1047));
  NAND4_X1  g846(.A1(new_n989), .A2(new_n531), .A3(new_n1039), .A4(new_n1047), .ZN(new_n1048));
  NAND3_X1  g847(.A1(new_n1046), .A2(KEYINPUT126), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g848(.A(KEYINPUT125), .ZN(new_n1050));
  NAND2_X1  g849(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g850(.A1(new_n1046), .A2(KEYINPUT125), .A3(new_n1048), .ZN(new_n1052));
  INV_X1    g851(.A(KEYINPUT127), .ZN(new_n1053));
  AND3_X1   g852(.A1(new_n1052), .A2(new_n1053), .A3(KEYINPUT60), .ZN(new_n1054));
  AOI21_X1  g853(.A(new_n1053), .B1(new_n1052), .B2(KEYINPUT60), .ZN(new_n1055));
  OAI21_X1  g854(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g855(.A1(new_n1052), .A2(KEYINPUT60), .ZN(new_n1057));
  NAND2_X1  g856(.A1(new_n1057), .A2(KEYINPUT127), .ZN(new_n1058));
  INV_X1    g857(.A(new_n1051), .ZN(new_n1059));
  NAND3_X1  g858(.A1(new_n1052), .A2(new_n1053), .A3(KEYINPUT60), .ZN(new_n1060));
  NAND3_X1  g859(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AND2_X1   g860(.A1(new_n1056), .A2(new_n1061), .ZN(G1350gat));
  OAI21_X1  g861(.A(G190gat), .B1(new_n1034), .B2(new_n802), .ZN(new_n1063));
  XNOR2_X1  g862(.A(new_n1063), .B(KEYINPUT61), .ZN(new_n1064));
  NAND2_X1  g863(.A1(new_n791), .A2(new_n244), .ZN(new_n1065));
  OAI21_X1  g864(.A(new_n1064), .B1(new_n1043), .B2(new_n1065), .ZN(G1351gat));
  NOR2_X1   g865(.A1(new_n779), .A2(new_n1027), .ZN(new_n1067));
  NAND2_X1  g866(.A1(new_n1011), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g867(.A(G197gat), .ZN(new_n1069));
  NOR3_X1   g868(.A1(new_n1068), .A2(new_n1069), .A3(new_n617), .ZN(new_n1070));
  NOR2_X1   g869(.A1(new_n996), .A2(new_n532), .ZN(new_n1071));
  NAND2_X1  g870(.A1(new_n1037), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g871(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g872(.A(G197gat), .B1(new_n1073), .B2(new_n874), .ZN(new_n1074));
  NOR2_X1   g873(.A1(new_n1070), .A2(new_n1074), .ZN(G1352gat));
  NOR3_X1   g874(.A1(new_n1072), .A2(G204gat), .A3(new_n901), .ZN(new_n1076));
  XNOR2_X1  g875(.A(new_n1076), .B(KEYINPUT62), .ZN(new_n1077));
  NAND3_X1  g876(.A1(new_n1011), .A2(new_n758), .A3(new_n1067), .ZN(new_n1078));
  NAND2_X1  g877(.A1(new_n1078), .A2(G204gat), .ZN(new_n1079));
  NAND2_X1  g878(.A1(new_n1077), .A2(new_n1079), .ZN(G1353gat));
  NAND3_X1  g879(.A1(new_n1073), .A2(new_n329), .A3(new_n676), .ZN(new_n1081));
  NAND3_X1  g880(.A1(new_n1011), .A2(new_n676), .A3(new_n1067), .ZN(new_n1082));
  AND3_X1   g881(.A1(new_n1082), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1083));
  AOI21_X1  g882(.A(KEYINPUT63), .B1(new_n1082), .B2(G211gat), .ZN(new_n1084));
  OAI21_X1  g883(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(G1354gat));
  OAI21_X1  g884(.A(G218gat), .B1(new_n1068), .B2(new_n802), .ZN(new_n1086));
  NAND3_X1  g885(.A1(new_n1073), .A2(new_n330), .A3(new_n791), .ZN(new_n1087));
  NAND2_X1  g886(.A1(new_n1086), .A2(new_n1087), .ZN(G1355gat));
endmodule


