

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704;

  XNOR2_X1 U358 ( .A(n503), .B(KEYINPUT32), .ZN(n699) );
  NOR2_X1 U359 ( .A1(n563), .A2(n355), .ZN(n603) );
  XNOR2_X1 U360 ( .A(n540), .B(KEYINPUT1), .ZN(n623) );
  XNOR2_X1 U361 ( .A(n363), .B(n362), .ZN(n484) );
  XNOR2_X1 U362 ( .A(n364), .B(G107), .ZN(n363) );
  XNOR2_X1 U363 ( .A(KEYINPUT92), .B(G110), .ZN(n362) );
  INV_X2 U364 ( .A(G104), .ZN(n364) );
  XNOR2_X1 U365 ( .A(KEYINPUT4), .B(KEYINPUT67), .ZN(n686) );
  INV_X1 U366 ( .A(n541), .ZN(n621) );
  XNOR2_X1 U367 ( .A(n495), .B(G472), .ZN(n541) );
  XNOR2_X1 U368 ( .A(n489), .B(n488), .ZN(n540) );
  INV_X2 U369 ( .A(G953), .ZN(n690) );
  NOR2_X2 U370 ( .A1(n663), .A2(n670), .ZN(n664) );
  NOR2_X2 U371 ( .A1(n531), .A2(n505), .ZN(n507) );
  XNOR2_X2 U372 ( .A(n501), .B(KEYINPUT22), .ZN(n505) );
  XNOR2_X2 U373 ( .A(n375), .B(n385), .ZN(n588) );
  NAND2_X1 U374 ( .A1(n580), .A2(n579), .ZN(n369) );
  INV_X1 U375 ( .A(G125), .ZN(n391) );
  AND2_X2 U376 ( .A1(n368), .A2(n369), .ZN(n668) );
  XNOR2_X1 U377 ( .A(n569), .B(KEYINPUT107), .ZN(n697) );
  NOR2_X1 U378 ( .A1(n374), .A2(n372), .ZN(n569) );
  NOR2_X1 U379 ( .A1(n515), .A2(n496), .ZN(n497) );
  NOR2_X1 U380 ( .A1(n635), .A2(n384), .ZN(n500) );
  NAND2_X1 U381 ( .A1(n398), .A2(n396), .ZN(n537) );
  INV_X1 U382 ( .A(n499), .ZN(n384) );
  AND2_X1 U383 ( .A1(n399), .A2(n401), .ZN(n398) );
  NAND2_X1 U384 ( .A1(n397), .A2(n400), .ZN(n396) );
  XNOR2_X1 U385 ( .A(n391), .B(G146), .ZN(n441) );
  XNOR2_X1 U386 ( .A(n429), .B(G128), .ZN(n440) );
  XOR2_X1 U387 ( .A(KEYINPUT15), .B(G902), .Z(n582) );
  INV_X1 U388 ( .A(G143), .ZN(n429) );
  XNOR2_X1 U389 ( .A(n440), .B(n430), .ZN(n481) );
  INV_X1 U390 ( .A(G134), .ZN(n430) );
  NOR2_X1 U391 ( .A1(G902), .A2(n654), .ZN(n489) );
  NAND2_X1 U392 ( .A1(n668), .A2(G217), .ZN(n395) );
  INV_X1 U393 ( .A(KEYINPUT73), .ZN(n347) );
  XNOR2_X1 U394 ( .A(KEYINPUT70), .B(G119), .ZN(n357) );
  INV_X1 U395 ( .A(KEYINPUT44), .ZN(n353) );
  INV_X1 U396 ( .A(n700), .ZN(n381) );
  XNOR2_X1 U397 ( .A(n479), .B(G146), .ZN(n376) );
  NOR2_X1 U398 ( .A1(n702), .A2(n406), .ZN(n405) );
  INV_X1 U399 ( .A(n613), .ZN(n406) );
  NOR2_X1 U400 ( .A1(n338), .A2(n582), .ZN(n400) );
  XNOR2_X1 U401 ( .A(n434), .B(n431), .ZN(n390) );
  XNOR2_X1 U402 ( .A(G122), .B(KEYINPUT102), .ZN(n427) );
  XNOR2_X1 U403 ( .A(n389), .B(KEYINPUT100), .ZN(n388) );
  INV_X1 U404 ( .A(KEYINPUT9), .ZN(n389) );
  AND2_X1 U405 ( .A1(n606), .A2(n531), .ZN(n532) );
  AND2_X1 U406 ( .A1(n373), .A2(n412), .ZN(n567) );
  INV_X1 U407 ( .A(n552), .ZN(n412) );
  NOR2_X1 U408 ( .A1(n550), .A2(n551), .ZN(n373) );
  INV_X1 U409 ( .A(n568), .ZN(n411) );
  XNOR2_X1 U410 ( .A(n437), .B(G478), .ZN(n513) );
  NOR2_X1 U411 ( .A1(n666), .A2(G902), .ZN(n437) );
  XNOR2_X1 U412 ( .A(KEYINPUT0), .B(KEYINPUT65), .ZN(n460) );
  INV_X1 U413 ( .A(n530), .ZN(n617) );
  XNOR2_X1 U414 ( .A(n470), .B(n349), .ZN(n669) );
  XNOR2_X1 U415 ( .A(n471), .B(n469), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n422), .B(n421), .ZN(n660) );
  XNOR2_X1 U417 ( .A(G113), .B(G104), .ZN(n420) );
  AND2_X1 U418 ( .A1(n614), .A2(n582), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n348), .B(n347), .ZN(n572) );
  NAND2_X1 U420 ( .A1(n338), .A2(n582), .ZN(n401) );
  XNOR2_X1 U421 ( .A(G131), .B(KEYINPUT5), .ZN(n490) );
  XNOR2_X1 U422 ( .A(n481), .B(n480), .ZN(n684) );
  INV_X1 U423 ( .A(G137), .ZN(n480) );
  XNOR2_X1 U424 ( .A(KEYINPUT72), .B(G122), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n356), .B(n439), .ZN(n493) );
  XNOR2_X1 U426 ( .A(n357), .B(n378), .ZN(n356) );
  INV_X1 U427 ( .A(KEYINPUT3), .ZN(n378) );
  XNOR2_X1 U428 ( .A(KEYINPUT83), .B(KEYINPUT8), .ZN(n432) );
  XOR2_X1 U429 ( .A(KEYINPUT7), .B(KEYINPUT99), .Z(n428) );
  XNOR2_X1 U430 ( .A(G140), .B(G131), .ZN(n482) );
  XNOR2_X1 U431 ( .A(n445), .B(KEYINPUT79), .ZN(n446) );
  AND2_X1 U432 ( .A1(G224), .A2(n690), .ZN(n445) );
  XNOR2_X1 U433 ( .A(n686), .B(G101), .ZN(n479) );
  XNOR2_X1 U434 ( .A(n444), .B(n345), .ZN(n448) );
  XNOR2_X1 U435 ( .A(n346), .B(n441), .ZN(n345) );
  XNOR2_X1 U436 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n442) );
  INV_X1 U437 ( .A(KEYINPUT84), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n358), .B(n493), .ZN(n677) );
  XNOR2_X1 U439 ( .A(n484), .B(n359), .ZN(n358) );
  XNOR2_X1 U440 ( .A(n361), .B(n360), .ZN(n359) );
  INV_X1 U441 ( .A(KEYINPUT16), .ZN(n360) );
  XNOR2_X1 U442 ( .A(G140), .B(KEYINPUT95), .ZN(n464) );
  XNOR2_X1 U443 ( .A(G119), .B(G110), .ZN(n462) );
  XNOR2_X1 U444 ( .A(G122), .B(G143), .ZN(n417) );
  XOR2_X1 U445 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n418) );
  XNOR2_X1 U446 ( .A(n377), .B(n375), .ZN(n654) );
  XNOR2_X1 U447 ( .A(n487), .B(KEYINPUT78), .ZN(n377) );
  XNOR2_X1 U448 ( .A(n486), .B(n485), .ZN(n487) );
  NAND2_X1 U449 ( .A1(n578), .A2(n367), .ZN(n614) );
  NOR2_X1 U450 ( .A1(n581), .A2(n579), .ZN(n367) );
  XNOR2_X1 U451 ( .A(n425), .B(n424), .ZN(n511) );
  XNOR2_X1 U452 ( .A(n423), .B(G475), .ZN(n424) );
  INV_X1 U453 ( .A(KEYINPUT13), .ZN(n423) );
  XNOR2_X1 U454 ( .A(n390), .B(n387), .ZN(n435) );
  XNOR2_X1 U455 ( .A(G116), .B(G107), .ZN(n426) );
  XOR2_X1 U456 ( .A(KEYINPUT106), .B(n539), .Z(n702) );
  XNOR2_X1 U457 ( .A(n382), .B(KEYINPUT35), .ZN(n700) );
  NAND2_X1 U458 ( .A1(n567), .A2(n411), .ZN(n372) );
  NOR2_X1 U459 ( .A1(n512), .A2(n511), .ZN(n606) );
  AND2_X1 U460 ( .A1(n351), .A2(n350), .ZN(n591) );
  NAND2_X1 U461 ( .A1(n393), .A2(n350), .ZN(n392) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n393) );
  INV_X1 U463 ( .A(n669), .ZN(n394) );
  NAND2_X1 U464 ( .A1(n366), .A2(n350), .ZN(n365) );
  XNOR2_X1 U465 ( .A(n587), .B(n586), .ZN(n366) );
  INV_X1 U466 ( .A(KEYINPUT53), .ZN(n407) );
  AND2_X1 U467 ( .A1(G210), .A2(n451), .ZN(n338) );
  XNOR2_X1 U468 ( .A(n684), .B(n376), .ZN(n492) );
  INV_X1 U469 ( .A(n492), .ZN(n375) );
  AND2_X1 U470 ( .A1(n494), .A2(G210), .ZN(n339) );
  XOR2_X1 U471 ( .A(KEYINPUT104), .B(n438), .Z(n566) );
  XOR2_X1 U472 ( .A(KEYINPUT71), .B(KEYINPUT34), .Z(n340) );
  XOR2_X1 U473 ( .A(n588), .B(KEYINPUT62), .Z(n341) );
  XOR2_X1 U474 ( .A(n574), .B(KEYINPUT68), .Z(n342) );
  XOR2_X1 U475 ( .A(KEYINPUT45), .B(KEYINPUT85), .Z(n343) );
  NOR2_X1 U476 ( .A1(G952), .A2(n690), .ZN(n670) );
  INV_X1 U477 ( .A(n670), .ZN(n350) );
  XOR2_X1 U478 ( .A(KEYINPUT86), .B(KEYINPUT56), .Z(n344) );
  INV_X1 U479 ( .A(KEYINPUT2), .ZN(n579) );
  INV_X1 U480 ( .A(n578), .ZN(n671) );
  NAND2_X1 U481 ( .A1(n577), .A2(n578), .ZN(n580) );
  XNOR2_X2 U482 ( .A(n403), .B(n343), .ZN(n578) );
  XNOR2_X1 U483 ( .A(n354), .B(n353), .ZN(n404) );
  INV_X1 U484 ( .A(n440), .ZN(n346) );
  XNOR2_X2 U485 ( .A(n461), .B(n460), .ZN(n518) );
  NAND2_X1 U486 ( .A1(n571), .A2(n570), .ZN(n348) );
  XNOR2_X1 U487 ( .A(n589), .B(n341), .ZN(n351) );
  XNOR2_X1 U488 ( .A(n365), .B(n344), .ZN(G51) );
  XNOR2_X2 U489 ( .A(n352), .B(n453), .ZN(n355) );
  NAND2_X1 U490 ( .A1(n537), .A2(n632), .ZN(n352) );
  NAND2_X1 U491 ( .A1(n379), .A2(n381), .ZN(n354) );
  XNOR2_X1 U492 ( .A(n392), .B(KEYINPUT121), .ZN(G66) );
  NOR2_X2 U493 ( .A1(n355), .A2(n459), .ZN(n461) );
  XNOR2_X1 U494 ( .A(n369), .B(KEYINPUT80), .ZN(n615) );
  INV_X1 U495 ( .A(n577), .ZN(n689) );
  XNOR2_X2 U496 ( .A(n581), .B(n370), .ZN(n577) );
  NAND2_X1 U497 ( .A1(n371), .A2(n405), .ZN(n581) );
  XNOR2_X1 U498 ( .A(n575), .B(n342), .ZN(n371) );
  INV_X1 U499 ( .A(n566), .ZN(n374) );
  XNOR2_X1 U500 ( .A(n380), .B(KEYINPUT91), .ZN(n379) );
  NAND2_X1 U501 ( .A1(n699), .A2(n599), .ZN(n380) );
  NAND2_X1 U502 ( .A1(n383), .A2(n566), .ZN(n382) );
  XNOR2_X1 U503 ( .A(n498), .B(n340), .ZN(n383) );
  NAND2_X1 U504 ( .A1(n513), .A2(n511), .ZN(n635) );
  XNOR2_X1 U505 ( .A(n493), .B(n386), .ZN(n385) );
  XNOR2_X1 U506 ( .A(n491), .B(n339), .ZN(n386) );
  XNOR2_X1 U507 ( .A(n481), .B(n388), .ZN(n387) );
  NAND2_X1 U508 ( .A1(n524), .A2(n404), .ZN(n403) );
  NOR2_X2 U509 ( .A1(n588), .A2(G902), .ZN(n495) );
  INV_X1 U510 ( .A(n583), .ZN(n397) );
  NAND2_X1 U511 ( .A1(n583), .A2(n338), .ZN(n399) );
  XNOR2_X2 U512 ( .A(n402), .B(n449), .ZN(n583) );
  INV_X1 U513 ( .A(n677), .ZN(n402) );
  XNOR2_X1 U514 ( .A(n408), .B(n407), .ZN(G75) );
  NAND2_X1 U515 ( .A1(n409), .A2(n690), .ZN(n408) );
  XNOR2_X1 U516 ( .A(n410), .B(KEYINPUT119), .ZN(n409) );
  NAND2_X1 U517 ( .A1(n653), .A2(n652), .ZN(n410) );
  NOR2_X2 U518 ( .A1(n573), .A2(n572), .ZN(n575) );
  BUF_X1 U519 ( .A(n541), .Z(n519) );
  XNOR2_X2 U520 ( .A(n555), .B(KEYINPUT40), .ZN(n703) );
  INV_X1 U521 ( .A(n537), .ZN(n568) );
  XNOR2_X1 U522 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U523 ( .A(n479), .B(n446), .ZN(n447) );
  AND2_X1 U524 ( .A1(n494), .A2(G214), .ZN(n413) );
  XOR2_X1 U525 ( .A(n419), .B(KEYINPUT11), .Z(n414) );
  XOR2_X1 U526 ( .A(n650), .B(KEYINPUT118), .Z(n415) );
  XNOR2_X1 U527 ( .A(n685), .B(n413), .ZN(n422) );
  XNOR2_X1 U528 ( .A(KEYINPUT69), .B(G469), .ZN(n488) );
  XNOR2_X1 U529 ( .A(n452), .B(KEYINPUT64), .ZN(n453) );
  XNOR2_X1 U530 ( .A(KEYINPUT63), .B(KEYINPUT109), .ZN(n590) );
  XNOR2_X1 U531 ( .A(n591), .B(n590), .ZN(G57) );
  INV_X1 U532 ( .A(n441), .ZN(n416) );
  XNOR2_X1 U533 ( .A(KEYINPUT10), .B(n416), .ZN(n471) );
  XNOR2_X1 U534 ( .A(n471), .B(n482), .ZN(n685) );
  NOR2_X1 U535 ( .A1(G953), .A2(G237), .ZN(n494) );
  XNOR2_X1 U536 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U537 ( .A(n414), .B(n420), .ZN(n421) );
  NOR2_X1 U538 ( .A1(G902), .A2(n660), .ZN(n425) );
  INV_X1 U539 ( .A(n511), .ZN(n514) );
  XNOR2_X1 U540 ( .A(n426), .B(KEYINPUT101), .ZN(n436) );
  XNOR2_X1 U541 ( .A(n428), .B(n427), .ZN(n431) );
  NAND2_X1 U542 ( .A1(n690), .A2(G234), .ZN(n433) );
  XNOR2_X1 U543 ( .A(n433), .B(n432), .ZN(n468) );
  NAND2_X1 U544 ( .A1(G217), .A2(n468), .ZN(n434) );
  XNOR2_X1 U545 ( .A(n436), .B(n435), .ZN(n666) );
  INV_X1 U546 ( .A(n513), .ZN(n512) );
  NAND2_X1 U547 ( .A1(n514), .A2(n512), .ZN(n438) );
  XNOR2_X1 U548 ( .A(G116), .B(G113), .ZN(n439) );
  XOR2_X1 U549 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n443) );
  XNOR2_X1 U550 ( .A(n443), .B(n442), .ZN(n444) );
  NOR2_X1 U551 ( .A1(G902), .A2(G237), .ZN(n450) );
  XOR2_X1 U552 ( .A(KEYINPUT76), .B(n450), .Z(n451) );
  NAND2_X1 U553 ( .A1(n451), .A2(G214), .ZN(n632) );
  INV_X1 U554 ( .A(KEYINPUT19), .ZN(n452) );
  NAND2_X1 U555 ( .A1(G234), .A2(G237), .ZN(n454) );
  XNOR2_X1 U556 ( .A(n454), .B(KEYINPUT14), .ZN(n455) );
  XNOR2_X1 U557 ( .A(KEYINPUT74), .B(n455), .ZN(n456) );
  NAND2_X1 U558 ( .A1(G952), .A2(n456), .ZN(n647) );
  NOR2_X1 U559 ( .A1(G953), .A2(n647), .ZN(n527) );
  AND2_X1 U560 ( .A1(n456), .A2(G953), .ZN(n457) );
  NAND2_X1 U561 ( .A1(G902), .A2(n457), .ZN(n525) );
  NOR2_X1 U562 ( .A1(n525), .A2(G898), .ZN(n458) );
  NOR2_X1 U563 ( .A1(n527), .A2(n458), .ZN(n459) );
  XOR2_X1 U564 ( .A(G137), .B(G128), .Z(n463) );
  XNOR2_X1 U565 ( .A(n463), .B(n462), .ZN(n467) );
  XOR2_X1 U566 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n465) );
  XNOR2_X1 U567 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U568 ( .A(n467), .B(n466), .Z(n470) );
  NAND2_X1 U569 ( .A1(G221), .A2(n468), .ZN(n469) );
  NOR2_X1 U570 ( .A1(G902), .A2(n669), .ZN(n476) );
  INV_X1 U571 ( .A(n582), .ZN(n472) );
  NAND2_X1 U572 ( .A1(G234), .A2(n472), .ZN(n473) );
  XNOR2_X1 U573 ( .A(KEYINPUT20), .B(n473), .ZN(n477) );
  NAND2_X1 U574 ( .A1(n477), .A2(G217), .ZN(n474) );
  XOR2_X1 U575 ( .A(KEYINPUT25), .B(n474), .Z(n475) );
  XNOR2_X1 U576 ( .A(n476), .B(n475), .ZN(n530) );
  NAND2_X1 U577 ( .A1(n477), .A2(G221), .ZN(n478) );
  XNOR2_X1 U578 ( .A(n478), .B(KEYINPUT21), .ZN(n528) );
  INV_X1 U579 ( .A(n528), .ZN(n616) );
  XNOR2_X1 U580 ( .A(n616), .B(KEYINPUT96), .ZN(n499) );
  AND2_X1 U581 ( .A1(n617), .A2(n499), .ZN(n624) );
  INV_X1 U582 ( .A(n482), .ZN(n483) );
  XNOR2_X1 U583 ( .A(n484), .B(n483), .ZN(n486) );
  NAND2_X1 U584 ( .A1(G227), .A2(n690), .ZN(n485) );
  NAND2_X1 U585 ( .A1(n624), .A2(n623), .ZN(n515) );
  XNOR2_X1 U586 ( .A(n490), .B(KEYINPUT77), .ZN(n491) );
  XOR2_X1 U587 ( .A(n621), .B(KEYINPUT6), .Z(n531) );
  INV_X1 U588 ( .A(n531), .ZN(n496) );
  XNOR2_X1 U589 ( .A(n497), .B(KEYINPUT33), .ZN(n648) );
  NOR2_X1 U590 ( .A1(n518), .A2(n648), .ZN(n498) );
  INV_X1 U591 ( .A(n518), .ZN(n516) );
  NAND2_X1 U592 ( .A1(n516), .A2(n500), .ZN(n501) );
  INV_X1 U593 ( .A(n623), .ZN(n534) );
  NOR2_X1 U594 ( .A1(n617), .A2(n534), .ZN(n502) );
  NAND2_X1 U595 ( .A1(n507), .A2(n502), .ZN(n503) );
  NAND2_X1 U596 ( .A1(n534), .A2(n519), .ZN(n504) );
  NOR2_X1 U597 ( .A1(n505), .A2(n504), .ZN(n506) );
  NAND2_X1 U598 ( .A1(n530), .A2(n506), .ZN(n599) );
  XOR2_X1 U599 ( .A(n507), .B(KEYINPUT90), .Z(n508) );
  NOR2_X1 U600 ( .A1(n623), .A2(n508), .ZN(n509) );
  NAND2_X1 U601 ( .A1(n509), .A2(n617), .ZN(n510) );
  XNOR2_X1 U602 ( .A(KEYINPUT103), .B(n510), .ZN(n698) );
  NOR2_X1 U603 ( .A1(n514), .A2(n513), .ZN(n608) );
  NOR2_X1 U604 ( .A1(n606), .A2(n608), .ZN(n637) );
  NOR2_X1 U605 ( .A1(n519), .A2(n515), .ZN(n629) );
  NAND2_X1 U606 ( .A1(n629), .A2(n516), .ZN(n517) );
  XNOR2_X1 U607 ( .A(KEYINPUT31), .B(n517), .ZN(n609) );
  NAND2_X1 U608 ( .A1(n540), .A2(n624), .ZN(n552) );
  NOR2_X1 U609 ( .A1(n518), .A2(n552), .ZN(n520) );
  NAND2_X1 U610 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U611 ( .A(KEYINPUT97), .B(n521), .ZN(n594) );
  NOR2_X1 U612 ( .A1(n609), .A2(n594), .ZN(n522) );
  NOR2_X1 U613 ( .A1(n637), .A2(n522), .ZN(n523) );
  NOR2_X1 U614 ( .A1(n698), .A2(n523), .ZN(n524) );
  XOR2_X1 U615 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n536) );
  NOR2_X1 U616 ( .A1(G900), .A2(n525), .ZN(n526) );
  NOR2_X1 U617 ( .A1(n527), .A2(n526), .ZN(n551) );
  NOR2_X1 U618 ( .A1(n551), .A2(n528), .ZN(n529) );
  NAND2_X1 U619 ( .A1(n530), .A2(n529), .ZN(n542) );
  NAND2_X1 U620 ( .A1(n532), .A2(n632), .ZN(n533) );
  NOR2_X1 U621 ( .A1(n542), .A2(n533), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n534), .A2(n558), .ZN(n535) );
  XNOR2_X1 U623 ( .A(n536), .B(n535), .ZN(n538) );
  NAND2_X1 U624 ( .A1(n538), .A2(n568), .ZN(n539) );
  INV_X1 U625 ( .A(n540), .ZN(n545) );
  NOR2_X1 U626 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U627 ( .A(KEYINPUT28), .B(n543), .Z(n544) );
  OR2_X1 U628 ( .A1(n545), .A2(n544), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT75), .B(KEYINPUT38), .Z(n546) );
  XNOR2_X1 U630 ( .A(n568), .B(n546), .ZN(n633) );
  NAND2_X1 U631 ( .A1(n633), .A2(n632), .ZN(n638) );
  NOR2_X1 U632 ( .A1(n635), .A2(n638), .ZN(n547) );
  XNOR2_X1 U633 ( .A(n547), .B(KEYINPUT41), .ZN(n649) );
  OR2_X1 U634 ( .A1(n563), .A2(n649), .ZN(n548) );
  XNOR2_X1 U635 ( .A(n548), .B(KEYINPUT42), .ZN(n704) );
  NAND2_X1 U636 ( .A1(n621), .A2(n632), .ZN(n549) );
  XNOR2_X1 U637 ( .A(KEYINPUT30), .B(n549), .ZN(n550) );
  AND2_X1 U638 ( .A1(n633), .A2(n567), .ZN(n554) );
  XNOR2_X1 U639 ( .A(KEYINPUT89), .B(KEYINPUT39), .ZN(n553) );
  XNOR2_X1 U640 ( .A(n554), .B(n553), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n576), .A2(n606), .ZN(n555) );
  NAND2_X1 U642 ( .A1(n704), .A2(n703), .ZN(n557) );
  XOR2_X1 U643 ( .A(KEYINPUT46), .B(KEYINPUT88), .Z(n556) );
  XNOR2_X1 U644 ( .A(n557), .B(n556), .ZN(n562) );
  AND2_X1 U645 ( .A1(n411), .A2(n558), .ZN(n560) );
  XNOR2_X1 U646 ( .A(KEYINPUT108), .B(KEYINPUT36), .ZN(n559) );
  XNOR2_X1 U647 ( .A(n560), .B(n559), .ZN(n561) );
  NAND2_X1 U648 ( .A1(n623), .A2(n561), .ZN(n612) );
  NAND2_X1 U649 ( .A1(n562), .A2(n612), .ZN(n573) );
  NAND2_X1 U650 ( .A1(n603), .A2(KEYINPUT66), .ZN(n564) );
  NOR2_X1 U651 ( .A1(n637), .A2(n564), .ZN(n565) );
  XNOR2_X1 U652 ( .A(KEYINPUT47), .B(n565), .ZN(n571) );
  XNOR2_X1 U653 ( .A(n697), .B(KEYINPUT82), .ZN(n570) );
  XNOR2_X1 U654 ( .A(KEYINPUT87), .B(KEYINPUT48), .ZN(n574) );
  NAND2_X1 U655 ( .A1(n576), .A2(n608), .ZN(n613) );
  NAND2_X1 U656 ( .A1(n668), .A2(G210), .ZN(n587) );
  XOR2_X1 U657 ( .A(KEYINPUT81), .B(KEYINPUT55), .Z(n585) );
  XNOR2_X1 U658 ( .A(n583), .B(KEYINPUT54), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n585), .B(n584), .ZN(n586) );
  NAND2_X1 U660 ( .A1(G472), .A2(n668), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n594), .A2(n606), .ZN(n592) );
  XNOR2_X1 U662 ( .A(n592), .B(KEYINPUT110), .ZN(n593) );
  XNOR2_X1 U663 ( .A(G104), .B(n593), .ZN(G6) );
  XOR2_X1 U664 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n596) );
  NAND2_X1 U665 ( .A1(n594), .A2(n608), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U667 ( .A(G107), .B(n597), .ZN(G9) );
  XOR2_X1 U668 ( .A(G110), .B(KEYINPUT111), .Z(n598) );
  XNOR2_X1 U669 ( .A(n599), .B(n598), .ZN(G12) );
  XOR2_X1 U670 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n601) );
  NAND2_X1 U671 ( .A1(n608), .A2(n603), .ZN(n600) );
  XNOR2_X1 U672 ( .A(n601), .B(n600), .ZN(n602) );
  XNOR2_X1 U673 ( .A(G128), .B(n602), .ZN(G30) );
  XOR2_X1 U674 ( .A(G146), .B(KEYINPUT113), .Z(n605) );
  NAND2_X1 U675 ( .A1(n603), .A2(n606), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n605), .B(n604), .ZN(G48) );
  NAND2_X1 U677 ( .A1(n609), .A2(n606), .ZN(n607) );
  XNOR2_X1 U678 ( .A(n607), .B(G113), .ZN(G15) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U680 ( .A(n610), .B(G116), .ZN(G18) );
  XOR2_X1 U681 ( .A(G125), .B(KEYINPUT37), .Z(n611) );
  XNOR2_X1 U682 ( .A(n612), .B(n611), .ZN(G27) );
  XNOR2_X1 U683 ( .A(G134), .B(n613), .ZN(G36) );
  NAND2_X1 U684 ( .A1(n615), .A2(n614), .ZN(n653) );
  NOR2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n619) );
  XOR2_X1 U686 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n618) );
  XNOR2_X1 U687 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X1 U688 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U689 ( .A(KEYINPUT115), .B(n622), .ZN(n627) );
  NOR2_X1 U690 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U691 ( .A(KEYINPUT50), .B(n625), .ZN(n626) );
  NOR2_X1 U692 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U693 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U694 ( .A(KEYINPUT51), .B(n630), .Z(n631) );
  NOR2_X1 U695 ( .A1(n649), .A2(n631), .ZN(n644) );
  NOR2_X1 U696 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U697 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U698 ( .A(n636), .B(KEYINPUT116), .ZN(n640) );
  NOR2_X1 U699 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U700 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U701 ( .A1(n641), .A2(n648), .ZN(n642) );
  XOR2_X1 U702 ( .A(KEYINPUT117), .B(n642), .Z(n643) );
  NOR2_X1 U703 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U704 ( .A(n645), .B(KEYINPUT52), .ZN(n646) );
  NOR2_X1 U705 ( .A1(n647), .A2(n646), .ZN(n651) );
  OR2_X1 U706 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U707 ( .A1(n651), .A2(n415), .ZN(n652) );
  XOR2_X1 U708 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n656) );
  XNOR2_X1 U709 ( .A(n654), .B(KEYINPUT120), .ZN(n655) );
  XNOR2_X1 U710 ( .A(n656), .B(n655), .ZN(n658) );
  NAND2_X1 U711 ( .A1(n668), .A2(G469), .ZN(n657) );
  XNOR2_X1 U712 ( .A(n658), .B(n657), .ZN(n659) );
  NOR2_X1 U713 ( .A1(n670), .A2(n659), .ZN(G54) );
  XOR2_X1 U714 ( .A(n660), .B(KEYINPUT59), .Z(n662) );
  NAND2_X1 U715 ( .A1(n668), .A2(G475), .ZN(n661) );
  XNOR2_X1 U716 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U717 ( .A(n664), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U718 ( .A1(G478), .A2(n668), .ZN(n665) );
  XNOR2_X1 U719 ( .A(n666), .B(n665), .ZN(n667) );
  NOR2_X1 U720 ( .A1(n670), .A2(n667), .ZN(G63) );
  OR2_X1 U721 ( .A1(G953), .A2(n671), .ZN(n675) );
  NAND2_X1 U722 ( .A1(G953), .A2(G224), .ZN(n672) );
  XNOR2_X1 U723 ( .A(KEYINPUT61), .B(n672), .ZN(n673) );
  NAND2_X1 U724 ( .A1(n673), .A2(G898), .ZN(n674) );
  NAND2_X1 U725 ( .A1(n675), .A2(n674), .ZN(n682) );
  XNOR2_X1 U726 ( .A(G101), .B(KEYINPUT122), .ZN(n676) );
  XNOR2_X1 U727 ( .A(n676), .B(KEYINPUT123), .ZN(n678) );
  XNOR2_X1 U728 ( .A(n678), .B(n677), .ZN(n680) );
  NOR2_X1 U729 ( .A1(n690), .A2(G898), .ZN(n679) );
  NOR2_X1 U730 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U731 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U732 ( .A(KEYINPUT124), .B(n683), .ZN(G69) );
  XNOR2_X1 U733 ( .A(n684), .B(KEYINPUT125), .ZN(n688) );
  XNOR2_X1 U734 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U735 ( .A(n688), .B(n687), .ZN(n692) );
  XNOR2_X1 U736 ( .A(n692), .B(n689), .ZN(n691) );
  NAND2_X1 U737 ( .A1(n691), .A2(n690), .ZN(n696) );
  XNOR2_X1 U738 ( .A(G227), .B(n692), .ZN(n693) );
  NAND2_X1 U739 ( .A1(n693), .A2(G900), .ZN(n694) );
  NAND2_X1 U740 ( .A1(n694), .A2(G953), .ZN(n695) );
  NAND2_X1 U741 ( .A1(n696), .A2(n695), .ZN(G72) );
  XNOR2_X1 U742 ( .A(n697), .B(G143), .ZN(G45) );
  XOR2_X1 U743 ( .A(G101), .B(n698), .Z(G3) );
  XNOR2_X1 U744 ( .A(n699), .B(G119), .ZN(G21) );
  XOR2_X1 U745 ( .A(G122), .B(n700), .Z(n701) );
  XNOR2_X1 U746 ( .A(KEYINPUT126), .B(n701), .ZN(G24) );
  XOR2_X1 U747 ( .A(G140), .B(n702), .Z(G42) );
  XNOR2_X1 U748 ( .A(G131), .B(n703), .ZN(G33) );
  XNOR2_X1 U749 ( .A(G137), .B(n704), .ZN(G39) );
endmodule

