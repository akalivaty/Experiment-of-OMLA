//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1253, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n204), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(G58), .A2(G68), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n224), .A2(G50), .A3(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n209), .B1(KEYINPUT1), .B2(new_n219), .C1(new_n222), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT65), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n227), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(new_n212), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT10), .ZN(new_n246));
  INV_X1    g0046(.A(G150), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NOR3_X1   g0049(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n250));
  OAI22_X1  g0050(.A1(new_n247), .A2(new_n249), .B1(new_n250), .B2(new_n204), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n204), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n251), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n220), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n261), .B1(new_n203), .B2(G20), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n262), .B(KEYINPUT69), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(new_n259), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G50), .B2(new_n264), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT9), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n273), .A3(G274), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT66), .B(G226), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(G222), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  INV_X1    g0086(.A(G223), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(G1698), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n285), .B1(new_n286), .B2(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n273), .ZN(new_n290));
  AOI211_X1 g0090(.A(new_n275), .B(new_n280), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G190), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n246), .A2(KEYINPUT73), .ZN(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n292), .B(new_n293), .C1(new_n291), .C2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(KEYINPUT73), .B(new_n246), .C1(new_n268), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n267), .B(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n291), .A2(new_n294), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n246), .A2(KEYINPUT73), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n292), .A2(new_n293), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n298), .A2(new_n299), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n291), .A2(G169), .B1(new_n260), .B2(new_n266), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n291), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n296), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT16), .ZN(new_n308));
  INV_X1    g0108(.A(G68), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT7), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n284), .B2(G20), .ZN(new_n311));
  AND2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n309), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n211), .A2(new_n309), .ZN(new_n317));
  OAI21_X1  g0117(.A(G20), .B1(new_n317), .B2(new_n223), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n248), .A2(G159), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n308), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT7), .B1(new_n314), .B2(new_n204), .ZN(new_n322));
  NOR4_X1   g0122(.A1(new_n312), .A2(new_n313), .A3(new_n310), .A4(G20), .ZN(new_n323));
  OAI21_X1  g0123(.A(G68), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n320), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n321), .A2(new_n326), .A3(new_n258), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n258), .B1(new_n203), .B2(G20), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n253), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n264), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n253), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n273), .A2(G232), .A3(new_n276), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n274), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(G226), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G87), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT67), .ZN(new_n338));
  INV_X1    g0138(.A(G1698), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n340), .B(new_n341), .C1(new_n312), .C2(new_n313), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n336), .B(new_n337), .C1(new_n342), .C2(new_n287), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n335), .B1(new_n343), .B2(new_n290), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(G169), .ZN(new_n345));
  AOI211_X1 g0145(.A(G179), .B(new_n335), .C1(new_n343), .C2(new_n290), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n333), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT18), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT75), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n333), .A2(new_n347), .A3(KEYINPUT18), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT76), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n344), .A2(new_n294), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  AOI211_X1 g0156(.A(new_n356), .B(new_n335), .C1(new_n343), .C2(new_n290), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n354), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n344), .A2(G190), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(KEYINPUT76), .C1(new_n294), .C2(new_n344), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n333), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT17), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n333), .B1(new_n358), .B2(new_n360), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT17), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT18), .B1(new_n333), .B2(new_n347), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT75), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n353), .A2(new_n365), .A3(new_n367), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n331), .A2(new_n309), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT12), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT11), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n249), .A2(new_n261), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n254), .A2(new_n286), .B1(new_n204), .B2(G68), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n258), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI221_X1 g0176(.A(new_n372), .B1(new_n309), .B2(new_n329), .C1(new_n373), .C2(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n376), .A2(new_n373), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT14), .ZN(new_n381));
  INV_X1    g0181(.A(G238), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n274), .B1(new_n382), .B2(new_n277), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n283), .A2(new_n284), .A3(G226), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G97), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(new_n385), .C1(new_n212), .C2(new_n288), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n386), .B2(new_n290), .ZN(new_n387));
  XOR2_X1   g0187(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n388));
  AND2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n387), .A2(new_n388), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n381), .B(G169), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n387), .A2(new_n388), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT13), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n392), .B(G179), .C1(new_n393), .C2(new_n387), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n387), .B(new_n388), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n381), .B1(new_n396), .B2(G169), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n380), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(G200), .B1(new_n389), .B2(new_n390), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n392), .B(G190), .C1(new_n393), .C2(new_n387), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n379), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n275), .B1(G244), .B2(new_n278), .ZN(new_n403));
  INV_X1    g0203(.A(G107), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n288), .A2(new_n382), .B1(new_n404), .B2(new_n284), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT70), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n342), .B2(new_n212), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT70), .A4(G232), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n403), .B1(new_n409), .B2(new_n273), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n410), .A2(G179), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n328), .A2(G77), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n413), .A2(new_n254), .B1(new_n204), .B2(new_n286), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT71), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n252), .B(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n416), .B2(new_n248), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n412), .B1(G77), .B2(new_n264), .C1(new_n417), .C2(new_n259), .ZN(new_n418));
  INV_X1    g0218(.A(G169), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n410), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n411), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n410), .A2(new_n356), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n418), .B1(G200), .B2(new_n410), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT72), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI211_X1 g0225(.A(KEYINPUT72), .B(new_n418), .C1(G200), .C2(new_n410), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n421), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n307), .A2(new_n370), .A3(new_n402), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n204), .B(G68), .C1(new_n312), .C2(new_n313), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT19), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n204), .B1(new_n385), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G87), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(new_n213), .A3(new_n404), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n204), .A2(G33), .A3(G97), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n436), .A2(KEYINPUT82), .A3(new_n431), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT82), .B1(new_n436), .B2(new_n431), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n430), .B(new_n435), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n258), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n413), .A2(new_n331), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n203), .A2(G33), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n264), .A2(new_n442), .A3(new_n220), .A4(new_n257), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(new_n413), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT83), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n439), .A2(new_n258), .B1(new_n331), .B2(new_n413), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT83), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n444), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n270), .A2(G1), .ZN(new_n451));
  INV_X1    g0251(.A(G274), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n203), .A2(G45), .ZN(new_n454));
  INV_X1    g0254(.A(G250), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(new_n273), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G116), .ZN(new_n459));
  OAI211_X1 g0259(.A(G244), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n459), .B(new_n460), .C1(new_n342), .C2(new_n382), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n461), .B2(new_n290), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n462), .A2(new_n304), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n462), .A2(G169), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(G190), .ZN(new_n466));
  INV_X1    g0266(.A(new_n443), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G87), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n440), .A2(new_n441), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n461), .A2(new_n290), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n294), .B1(new_n470), .B2(new_n457), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n450), .A2(new_n465), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n313), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT3), .A2(G33), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(G303), .A3(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(G264), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n477));
  OAI21_X1  g0277(.A(G257), .B1(new_n312), .B2(new_n313), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n340), .A2(new_n341), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n290), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT5), .B(G41), .ZN(new_n482));
  INV_X1    g0282(.A(new_n220), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n482), .A2(new_n451), .B1(new_n483), .B2(new_n272), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n452), .B1(new_n483), .B2(new_n272), .ZN(new_n485));
  NOR2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n454), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n484), .A2(G270), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT20), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n204), .B1(new_n213), .B2(G33), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT78), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT78), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(G33), .A3(G283), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n258), .B1(new_n204), .B2(G116), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n492), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n495), .A2(new_n497), .ZN(new_n501));
  INV_X1    g0301(.A(new_n493), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G116), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n257), .A2(new_n220), .B1(G20), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(KEYINPUT20), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n331), .A2(new_n504), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n443), .B2(new_n504), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT84), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n491), .A2(new_n511), .A3(new_n512), .A4(G179), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n481), .A2(new_n490), .A3(G179), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n509), .B1(new_n500), .B2(new_n506), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT84), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n419), .B1(new_n481), .B2(new_n490), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(new_n511), .A3(KEYINPUT21), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT21), .B1(new_n518), .B2(new_n511), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT85), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n481), .A2(new_n490), .A3(G190), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n515), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n294), .B1(new_n481), .B2(new_n490), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n526), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n528), .A2(KEYINPUT85), .A3(new_n515), .A4(new_n524), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n473), .A2(new_n517), .A3(new_n522), .A4(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n331), .A2(KEYINPUT25), .A3(new_n404), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT25), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n264), .B2(G107), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n467), .A2(G107), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n204), .B(G87), .C1(new_n312), .C2(new_n313), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT22), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT22), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n284), .A2(new_n540), .A3(new_n204), .A4(G87), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n459), .A2(G20), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n204), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n404), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT24), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT24), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n542), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n537), .B1(new_n552), .B2(new_n258), .ZN(new_n553));
  OAI211_X1 g0353(.A(G257), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G294), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n554), .B(new_n555), .C1(new_n342), .C2(new_n455), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n290), .B1(G264), .B2(new_n484), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n489), .A2(new_n485), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n304), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n290), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n484), .A2(G264), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n560), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n559), .B1(new_n562), .B2(G169), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n532), .B1(new_n553), .B2(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n542), .A2(new_n550), .A3(new_n547), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n550), .B1(new_n542), .B2(new_n547), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n258), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n536), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n557), .A2(new_n558), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n419), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n568), .A2(KEYINPUT86), .A3(new_n570), .A4(new_n559), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n562), .A2(G190), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(G200), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n553), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n564), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n531), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT81), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT80), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n283), .A2(new_n284), .A3(G244), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(KEYINPUT77), .A3(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G250), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT79), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n284), .A2(KEYINPUT79), .A3(G250), .A4(G1698), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT77), .B1(new_n579), .B2(new_n580), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT4), .A4(G244), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n501), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n273), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n484), .A2(G257), .B1(new_n485), .B2(new_n489), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n578), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n579), .A2(new_n580), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT77), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n589), .A2(new_n501), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(new_n581), .A4(new_n586), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n290), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(KEYINPUT80), .A3(new_n593), .ZN(new_n602));
  AOI21_X1  g0402(.A(G169), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT6), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n604), .A2(new_n213), .A3(G107), .ZN(new_n605));
  XNOR2_X1  g0405(.A(G97), .B(G107), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n607), .A2(new_n204), .B1(new_n286), .B2(new_n249), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n404), .B1(new_n311), .B2(new_n315), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n258), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n331), .A2(new_n213), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n467), .A2(G97), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n601), .A2(new_n593), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(G179), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n577), .B1(new_n603), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT80), .B1(new_n601), .B2(new_n593), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n578), .B(new_n594), .C1(new_n600), .C2(new_n290), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n419), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n613), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n592), .A2(new_n594), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(new_n304), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(KEYINPUT81), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n595), .A2(new_n602), .A3(G190), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n613), .B1(new_n614), .B2(G200), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n576), .A2(new_n616), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n429), .A2(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n306), .ZN(new_n629));
  INV_X1    g0429(.A(new_n352), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(new_n368), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n366), .B(new_n364), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n401), .ZN(new_n634));
  INV_X1    g0434(.A(new_n421), .ZN(new_n635));
  OAI21_X1  g0435(.A(G169), .B1(new_n389), .B2(new_n390), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n394), .A3(new_n391), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n635), .B1(new_n638), .B2(new_n380), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n632), .B1(new_n634), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n296), .A2(new_n302), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n629), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n450), .A2(new_n465), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n616), .A2(new_n623), .A3(new_n626), .ZN(new_n645));
  INV_X1    g0445(.A(new_n466), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n447), .B(new_n468), .C1(new_n294), .C2(new_n462), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT87), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n472), .A2(KEYINPUT87), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n651), .A2(new_n574), .A3(new_n643), .ZN(new_n652));
  INV_X1    g0452(.A(new_n521), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n517), .A2(new_n653), .A3(new_n519), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n553), .A2(new_n563), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n644), .B1(new_n645), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n603), .A2(new_n615), .A3(new_n577), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT81), .B1(new_n619), .B2(new_n622), .ZN(new_n661));
  OAI211_X1 g0461(.A(KEYINPUT26), .B(new_n473), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n603), .A2(new_n615), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n649), .A2(new_n650), .B1(new_n450), .B2(new_n465), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT26), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n642), .B1(new_n669), .B2(new_n429), .ZN(G369));
  INV_X1    g0470(.A(KEYINPUT89), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT27), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT88), .A4(G13), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G213), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n675), .B1(new_n674), .B2(new_n676), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n671), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n674), .A2(new_n676), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n682), .A2(KEYINPUT89), .A3(G213), .A4(new_n677), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n515), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT90), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n527), .A2(new_n529), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n517), .A2(new_n653), .A3(new_n519), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n530), .A2(new_n522), .A3(KEYINPUT90), .A4(new_n517), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n688), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n691), .A2(new_n688), .ZN(new_n695));
  OAI21_X1  g0495(.A(G330), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n553), .A2(new_n687), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n575), .A2(new_n697), .B1(new_n656), .B2(new_n687), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n691), .A2(new_n687), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT91), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n686), .B(new_n702), .ZN(new_n703));
  OAI22_X1  g0503(.A1(new_n575), .A2(new_n701), .B1(new_n656), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n700), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n207), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n434), .A2(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n226), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  INV_X1    g0513(.A(G330), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n557), .A2(new_n462), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n514), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n595), .A2(new_n602), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT30), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n595), .A2(new_n602), .A3(new_n719), .A4(new_n716), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n491), .A2(G179), .A3(new_n462), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n614), .A2(new_n569), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n703), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n723), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n718), .B2(new_n720), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n726), .B1(new_n730), .B2(new_n687), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n645), .A2(new_n576), .A3(new_n725), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n714), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n473), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n616), .B2(new_n623), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n665), .B1(new_n736), .B2(KEYINPUT26), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n616), .A2(new_n623), .A3(new_n626), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n652), .A2(new_n657), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n643), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n725), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT29), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n664), .A2(new_n619), .A3(new_n622), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n644), .B1(new_n744), .B2(KEYINPUT26), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n564), .A2(new_n571), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n652), .B1(new_n746), .B2(new_n691), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n747), .B2(new_n738), .ZN(new_n748));
  AOI211_X1 g0548(.A(KEYINPUT26), .B(new_n735), .C1(new_n616), .C2(new_n623), .ZN(new_n749));
  OAI211_X1 g0549(.A(KEYINPUT29), .B(new_n687), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n734), .B1(new_n743), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n713), .B1(new_n751), .B2(G1), .ZN(G364));
  NOR3_X1   g0552(.A1(new_n694), .A2(G330), .A3(new_n695), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n204), .A2(G13), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n203), .B1(new_n754), .B2(G45), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n708), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n696), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n220), .B1(G20), .B2(new_n419), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT95), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n204), .A2(new_n304), .A3(new_n294), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT93), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT93), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n761), .B1(new_n765), .B2(G190), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n763), .A2(KEYINPUT95), .A3(new_n356), .A4(new_n764), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n304), .A2(G200), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G20), .A3(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n768), .A2(new_n769), .B1(G322), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT98), .Z(new_n774));
  NOR4_X1   g0574(.A1(new_n204), .A2(new_n294), .A3(G179), .A4(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  INV_X1    g0577(.A(G329), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n204), .A2(G190), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT97), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n765), .A2(new_n356), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G326), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n770), .A2(new_n779), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n314), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n204), .B1(new_n780), .B2(G190), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n788), .B1(G294), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G303), .ZN(new_n792));
  NOR4_X1   g0592(.A1(new_n204), .A2(new_n356), .A3(new_n294), .A4(G179), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT96), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n785), .B(new_n791), .C1(new_n792), .C2(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n774), .A2(new_n783), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n781), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G159), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT32), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n776), .A2(new_n404), .B1(new_n213), .B2(new_n789), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n314), .B1(new_n793), .B2(G87), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT94), .Z(new_n804));
  NAND2_X1  g0604(.A1(new_n784), .A2(G50), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n771), .A2(new_n211), .B1(new_n786), .B2(new_n286), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT92), .Z(new_n807));
  NAND4_X1  g0607(.A1(new_n802), .A2(new_n804), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G68), .B2(new_n768), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n760), .B1(new_n797), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n207), .A2(G355), .A3(new_n284), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n707), .A2(new_n284), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(G45), .B2(new_n226), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n241), .A2(new_n270), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n811), .B1(G116), .B2(new_n207), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G13), .A2(G33), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G20), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n760), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n758), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n810), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n818), .B(KEYINPUT99), .Z(new_n822));
  NOR3_X1   g0622(.A1(new_n694), .A2(new_n695), .A3(new_n822), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n753), .A2(new_n759), .B1(new_n821), .B2(new_n823), .ZN(G396));
  NOR2_X1   g0624(.A1(new_n421), .A2(new_n686), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n418), .A2(new_n686), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n425), .B2(new_n426), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n825), .B1(new_n827), .B2(new_n421), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n741), .A2(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n703), .B(new_n825), .C1(new_n827), .C2(new_n421), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n737), .B2(new_n740), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n627), .A2(new_n703), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n728), .A2(new_n731), .ZN(new_n835));
  OAI21_X1  g0635(.A(G330), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n757), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n836), .B2(new_n833), .ZN(new_n838));
  INV_X1    g0638(.A(new_n784), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n839), .A2(new_n792), .B1(new_n504), .B2(new_n786), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n768), .B2(G283), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT102), .ZN(new_n842));
  INV_X1    g0642(.A(G294), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n314), .B1(new_n771), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G311), .B2(new_n798), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n790), .A2(G97), .B1(new_n775), .B2(G87), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(new_n795), .C2(new_n404), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n314), .B1(new_n798), .B2(G132), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n848), .B1(new_n211), .B2(new_n789), .C1(new_n309), .C2(new_n776), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G50), .B2(new_n794), .ZN(new_n850));
  INV_X1    g0650(.A(new_n786), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n772), .A2(G143), .B1(new_n851), .B2(G159), .ZN(new_n852));
  INV_X1    g0652(.A(G137), .ZN(new_n853));
  INV_X1    g0653(.A(new_n768), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n852), .B1(new_n853), .B2(new_n839), .C1(new_n854), .C2(new_n247), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n850), .B1(new_n856), .B2(KEYINPUT34), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT34), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n842), .A2(new_n847), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n760), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n760), .A2(new_n816), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT100), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n757), .B1(new_n863), .B2(G77), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT101), .Z(new_n865));
  OAI211_X1 g0665(.A(new_n861), .B(new_n865), .C1(new_n817), .C2(new_n828), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n838), .A2(new_n866), .ZN(G384));
  NOR2_X1   g0667(.A1(new_n754), .A2(new_n203), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n680), .A2(KEYINPUT107), .A3(new_n683), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT107), .B1(new_n680), .B2(new_n683), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT37), .B1(new_n872), .B2(new_n333), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT106), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n333), .A2(new_n347), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n333), .B2(new_n347), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n363), .B(new_n873), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT108), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n363), .A2(new_n879), .A3(new_n348), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n343), .A2(new_n290), .ZN(new_n881));
  INV_X1    g0681(.A(new_n335), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n304), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(G169), .B2(new_n344), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n327), .B2(new_n332), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT108), .B1(new_n366), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n872), .A2(new_n333), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n880), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n878), .B1(new_n888), .B2(KEYINPUT37), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n633), .B2(new_n632), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n869), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n362), .A2(new_n684), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n370), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n885), .B1(new_n362), .B2(new_n361), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT105), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n892), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT105), .B1(new_n366), .B2(new_n885), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(KEYINPUT38), .B(new_n893), .C1(new_n899), .C2(new_n878), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n891), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n731), .B(new_n902), .C1(new_n627), .C2(new_n703), .ZN(new_n903));
  INV_X1    g0703(.A(new_n401), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n380), .B(new_n686), .C1(new_n638), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n380), .A2(new_n686), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n398), .A2(new_n401), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n908), .A2(new_n828), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n901), .A2(new_n903), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n903), .A2(new_n911), .A3(new_n909), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n370), .A2(new_n892), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n363), .A2(new_n896), .A3(new_n348), .ZN(new_n914));
  INV_X1    g0714(.A(new_n892), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(new_n898), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n878), .B1(new_n916), .B2(KEYINPUT37), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n869), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n900), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n910), .A2(KEYINPUT40), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT109), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n903), .A2(new_n428), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n714), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n922), .B2(new_n921), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n827), .A2(new_n421), .ZN(new_n925));
  INV_X1    g0725(.A(new_n825), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(new_n725), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n659), .B2(new_n667), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT104), .B1(new_n928), .B2(new_n825), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT104), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n832), .A2(new_n930), .A3(new_n926), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n919), .A3(new_n908), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT39), .B1(new_n891), .B2(new_n900), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n918), .A2(new_n900), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n935), .B2(KEYINPUT39), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n638), .A2(new_n380), .A3(new_n687), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n872), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n631), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n933), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n743), .A2(new_n428), .A3(new_n750), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n642), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n868), .B1(new_n924), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n924), .ZN(new_n947));
  INV_X1    g0747(.A(new_n607), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n504), .B(new_n222), .C1(new_n948), .C2(KEYINPUT35), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(KEYINPUT35), .B2(new_n948), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT36), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n226), .A2(new_n286), .A3(new_n317), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n261), .B2(G68), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n953), .A2(new_n203), .A3(G13), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT103), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(new_n951), .A3(new_n955), .ZN(G367));
  NOR2_X1   g0756(.A1(new_n575), .A2(new_n701), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n703), .A2(new_n613), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n616), .A2(new_n623), .A3(new_n626), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n663), .A2(new_n703), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT42), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n960), .A2(new_n961), .B1(new_n564), .B2(new_n571), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n616), .A2(new_n623), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n725), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n686), .A2(new_n469), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n664), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n643), .B2(new_n967), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n963), .A2(new_n966), .B1(KEYINPUT43), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n700), .B1(new_n960), .B2(new_n961), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n972), .B(new_n973), .Z(new_n974));
  XOR2_X1   g0774(.A(new_n708), .B(KEYINPUT41), .Z(new_n975));
  INV_X1    g0775(.A(KEYINPUT111), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT29), .B1(new_n668), .B2(new_n725), .ZN(new_n977));
  INV_X1    g0777(.A(new_n750), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n836), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n701), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n958), .B1(new_n698), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT110), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n981), .B1(new_n696), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n696), .B(KEYINPUT110), .ZN(new_n985));
  INV_X1    g0785(.A(new_n981), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n976), .B1(new_n979), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n704), .B1(new_n960), .B2(new_n961), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT45), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n960), .A2(new_n704), .A3(new_n961), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT44), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n990), .A2(new_n993), .A3(new_n700), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n700), .B1(new_n990), .B2(new_n993), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n696), .B(new_n982), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n983), .B1(new_n997), .B2(new_n981), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n998), .A2(new_n751), .A3(KEYINPUT111), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n988), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(KEYINPUT112), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT112), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n988), .A2(new_n996), .A3(new_n1002), .A4(new_n999), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n975), .B1(new_n1004), .B2(new_n751), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n974), .B1(new_n1005), .B2(new_n756), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n812), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n819), .B1(new_n207), .B2(new_n413), .C1(new_n1007), .C2(new_n237), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n757), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n851), .A2(G283), .B1(new_n798), .B2(G317), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1010), .B(new_n314), .C1(new_n792), .C2(new_n771), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n793), .B2(G116), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n776), .A2(new_n213), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n789), .A2(new_n404), .ZN(new_n1015));
  NOR4_X1   g0815(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(KEYINPUT46), .A2(G116), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n784), .A2(G311), .B1(new_n794), .B2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1016), .B(new_n1018), .C1(new_n843), .C2(new_n854), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n772), .A2(G150), .B1(new_n798), .B2(G137), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n261), .B2(new_n786), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n314), .B1(new_n775), .B2(G77), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT114), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n793), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1025), .A2(new_n211), .B1(new_n309), .B2(new_n789), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1021), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n784), .A2(G143), .B1(new_n1023), .B2(new_n1022), .ZN(new_n1028));
  INV_X1    g0828(.A(G159), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1027), .B(new_n1028), .C1(new_n854), .C2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1019), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT47), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1009), .B1(new_n1032), .B2(new_n760), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n822), .B2(new_n969), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1006), .A2(new_n1034), .ZN(G387));
  NAND2_X1  g0835(.A1(new_n988), .A2(new_n999), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n708), .C1(new_n751), .C2(new_n998), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n710), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1038), .A2(new_n207), .A3(new_n284), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(G107), .B2(new_n207), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n416), .A2(new_n261), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT117), .Z(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT50), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(KEYINPUT50), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n270), .B1(new_n309), .B2(new_n286), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT115), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1045), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1046), .B2(new_n1038), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT116), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1043), .A2(new_n1044), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1007), .B1(new_n234), .B2(G45), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1040), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n819), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n757), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n784), .A2(G159), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT118), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n768), .A2(new_n253), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n314), .B1(new_n798), .B2(G150), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n261), .B2(new_n771), .C1(new_n309), .C2(new_n786), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1025), .A2(new_n286), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n789), .A2(new_n413), .ZN(new_n1061));
  NOR4_X1   g0861(.A1(new_n1059), .A2(new_n1014), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1056), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n284), .B1(new_n798), .B2(G326), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n1025), .A2(new_n843), .B1(new_n777), .B2(new_n789), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n772), .A2(G317), .B1(new_n851), .B2(G303), .ZN(new_n1066));
  INV_X1    g0866(.A(G322), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1066), .B1(new_n1067), .B2(new_n839), .C1(new_n854), .C2(new_n787), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT48), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1065), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT49), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1064), .B1(new_n504), .B2(new_n776), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1063), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1054), .B1(new_n1075), .B2(new_n760), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n698), .B2(new_n822), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1037), .B(new_n1077), .C1(new_n755), .C2(new_n987), .ZN(G393));
  INV_X1    g0878(.A(new_n996), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n709), .B1(new_n1036), .B2(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1004), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n960), .A2(new_n818), .A3(new_n961), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n784), .A2(G317), .B1(G311), .B2(new_n772), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n314), .B1(new_n781), .B2(new_n1067), .C1(new_n843), .C2(new_n786), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1025), .A2(new_n777), .B1(new_n776), .B2(new_n404), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G116), .C2(new_n790), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n854), .B2(new_n792), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n784), .A2(G150), .B1(G159), .B2(new_n772), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT51), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1025), .A2(new_n309), .B1(new_n286), .B2(new_n789), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n314), .B1(new_n798), .B2(G143), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n433), .B2(new_n776), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1091), .B(new_n1093), .C1(new_n416), .C2(new_n851), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n261), .B2(new_n854), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1084), .A2(new_n1088), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n760), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n819), .B1(new_n213), .B2(new_n207), .C1(new_n1007), .C2(new_n244), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1082), .A2(new_n757), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1079), .B2(new_n755), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1081), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G390));
  NAND3_X1  g0902(.A1(new_n903), .A2(G330), .A3(new_n428), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n943), .A2(new_n642), .A3(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(G330), .B(new_n828), .C1(new_n834), .C2(new_n835), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n908), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n903), .A2(G330), .A3(new_n909), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n932), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n734), .A2(new_n828), .A3(new_n908), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n687), .B(new_n925), .C1(new_n748), .C2(new_n749), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n926), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n903), .A2(G330), .A3(new_n828), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1106), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1111), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1104), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n934), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT39), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n919), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1106), .B1(new_n929), .B2(new_n931), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n938), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n937), .B(new_n901), .C1(new_n1114), .C2(new_n1106), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n1111), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1108), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1119), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1108), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n832), .A2(new_n930), .A3(new_n926), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n930), .B1(new_n832), .B2(new_n926), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n908), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n936), .B1(new_n1132), .B2(new_n937), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1125), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1129), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1124), .A2(new_n1125), .A3(new_n1111), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n1136), .A3(new_n1118), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1128), .A2(new_n708), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1135), .A2(new_n756), .A3(new_n1136), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n757), .B1(new_n863), .B2(new_n253), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n776), .A2(new_n309), .B1(new_n286), .B2(new_n789), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n314), .B1(new_n786), .B2(new_n213), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n771), .A2(new_n504), .B1(new_n781), .B2(new_n843), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n795), .B2(new_n433), .C1(new_n839), .C2(new_n777), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n854), .A2(new_n404), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n854), .A2(new_n853), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n784), .A2(G128), .ZN(new_n1148));
  INV_X1    g0948(.A(G132), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n771), .A2(new_n1149), .B1(new_n786), .B2(new_n1150), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n314), .B(new_n1151), .C1(G125), .C2(new_n798), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n793), .A2(G150), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT53), .Z(new_n1154));
  AOI22_X1  g0954(.A1(new_n790), .A2(G159), .B1(new_n775), .B2(G50), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1148), .A2(new_n1152), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1145), .A2(new_n1146), .B1(new_n1147), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1140), .B1(new_n1157), .B2(new_n760), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT119), .Z(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n936), .B2(new_n817), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1139), .A2(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1138), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(G378));
  AOI21_X1  g0963(.A(new_n1060), .B1(G68), .B2(new_n790), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n211), .B2(new_n776), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n314), .A2(new_n269), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n786), .A2(new_n413), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n771), .A2(new_n404), .B1(new_n781), .B2(new_n777), .ZN(new_n1168));
  NOR4_X1   g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n213), .B2(new_n854), .C1(new_n504), .C2(new_n839), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT58), .ZN(new_n1171));
  INV_X1    g0971(.A(G33), .ZN(new_n1172));
  AOI21_X1  g0972(.A(G50), .B1(new_n1172), .B2(new_n269), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1170), .A2(new_n1171), .B1(new_n1166), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1025), .A2(new_n1150), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n772), .A2(G128), .B1(new_n851), .B2(G137), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n247), .B2(new_n789), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(G125), .C2(new_n784), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1149), .B2(new_n854), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n775), .A2(G159), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G33), .B(G41), .C1(new_n798), .C2(G124), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1174), .B1(new_n1171), .B2(new_n1170), .C1(new_n1180), .C2(new_n1184), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1185), .A2(new_n760), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n757), .B1(new_n863), .B2(G50), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n267), .A2(new_n684), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n307), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n307), .A2(new_n1188), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1186), .B(new_n1187), .C1(new_n1194), .C2(new_n816), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT120), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1194), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n891), .A2(new_n900), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n903), .A2(new_n909), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT40), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n919), .A2(new_n911), .A3(new_n903), .A4(new_n909), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1197), .B1(new_n1202), .B2(G330), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n714), .B(new_n1194), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n942), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1194), .B1(new_n920), .B2(new_n714), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1202), .A2(G330), .A3(new_n1197), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n936), .A2(new_n938), .B1(new_n631), .B2(new_n940), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n933), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1205), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1196), .B1(new_n1210), .B2(new_n756), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1104), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1137), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT57), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1205), .B2(new_n1209), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n708), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1210), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1211), .B1(new_n1217), .B2(new_n1218), .ZN(G375));
  NAND2_X1  g1019(.A1(new_n1106), .A2(new_n816), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n757), .B1(new_n863), .B2(G68), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n854), .A2(new_n1150), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n771), .A2(new_n853), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G128), .B2(new_n798), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n314), .B1(new_n851), .B2(G150), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n790), .A2(G50), .B1(new_n775), .B2(G58), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n1029), .B2(new_n795), .C1(new_n1149), .C2(new_n839), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n854), .A2(new_n504), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n776), .A2(new_n286), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n771), .A2(new_n777), .B1(new_n781), .B2(new_n792), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n314), .B1(new_n786), .B2(new_n404), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1061), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n795), .B2(new_n213), .C1(new_n839), .C2(new_n843), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n1222), .A2(new_n1228), .B1(new_n1229), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1221), .B1(new_n1235), .B2(new_n760), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1220), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1117), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1108), .A2(new_n1107), .B1(new_n929), .B2(new_n931), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1237), .B1(new_n1240), .B2(new_n755), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n975), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1110), .A2(new_n1104), .A3(new_n1117), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1119), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(G381));
  NOR2_X1   g1046(.A1(G375), .A2(G378), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1006), .A2(new_n1034), .A3(new_n1101), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(G407));
  AOI22_X1  g1050(.A1(new_n1137), .A2(new_n1212), .B1(new_n1209), .B2(new_n1205), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1216), .B(new_n708), .C1(KEYINPUT57), .C2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(new_n1162), .A3(new_n1211), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G407), .B(G213), .C1(G343), .C2(new_n1253), .ZN(G409));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(G393), .B(G396), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1101), .B1(new_n1006), .B2(new_n1034), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1248), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G387), .A2(G390), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1006), .A2(new_n1101), .A3(new_n1034), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1261), .A3(new_n1256), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1259), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G375), .A2(G378), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n685), .A2(G213), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1195), .B1(new_n1210), .B2(new_n756), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1138), .A2(new_n1267), .A3(new_n1161), .ZN(new_n1268));
  AOI221_X4 g1068(.A(new_n975), .B1(new_n1205), .B2(new_n1209), .C1(new_n1137), .C2(new_n1212), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1266), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(G384), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1244), .A2(KEYINPUT60), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1110), .A2(new_n1274), .A3(new_n1104), .A4(new_n1117), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n709), .B(new_n1118), .C1(new_n1273), .C2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1272), .B1(new_n1276), .B2(new_n1241), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1118), .A2(new_n709), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(G384), .A3(new_n1242), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1265), .A2(new_n1271), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1265), .A2(new_n1271), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1272), .B(new_n1241), .C1(new_n1278), .C2(new_n1279), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1280), .B2(new_n1242), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n685), .A2(G213), .A3(G2897), .ZN(new_n1290));
  XOR2_X1   g1090(.A(new_n1290), .B(KEYINPUT121), .Z(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1288), .A2(new_n1289), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT122), .B1(new_n1287), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1162), .B1(new_n1252), .B2(new_n1211), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1295), .B(KEYINPUT122), .C1(new_n1297), .C2(new_n1270), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1264), .B(new_n1286), .C1(new_n1296), .C2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1265), .A2(new_n1271), .A3(KEYINPUT63), .A4(new_n1283), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(KEYINPUT123), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1255), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT123), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1301), .B(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1259), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1285), .B2(new_n1284), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1295), .B1(new_n1297), .B2(new_n1270), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT122), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1298), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1305), .A2(new_n1307), .A3(new_n1311), .A4(KEYINPUT124), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1303), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT127), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1270), .B1(G378), .B2(G375), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT62), .B1(new_n1315), .B2(new_n1283), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT126), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NOR4_X1   g1118(.A1(new_n1297), .A2(new_n1270), .A3(new_n1318), .A4(new_n1282), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1316), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1284), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1321));
  XOR2_X1   g1121(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(new_n1287), .B2(new_n1295), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1314), .B1(new_n1320), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1284), .A2(new_n1318), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1315), .A2(KEYINPUT62), .A3(new_n1283), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1327), .A2(new_n1328), .A3(KEYINPUT126), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1329), .A2(KEYINPUT127), .A3(new_n1321), .A4(new_n1323), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1325), .A2(new_n1326), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1313), .A2(new_n1331), .ZN(G405));
  NAND2_X1  g1132(.A1(new_n1265), .A2(new_n1253), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1333), .B(new_n1282), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1334), .B(new_n1326), .ZN(G402));
endmodule


