//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n217), .A2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(G58), .A2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n212), .B1(new_n224), .B2(KEYINPUT1), .C1(new_n227), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n252), .A2(new_n254), .A3(G226), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT76), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT76), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n258), .A2(new_n259), .A3(G226), .A4(new_n255), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G97), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n257), .A2(new_n260), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n226), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT68), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(new_n264), .B2(new_n271), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n267), .A2(G1), .A3(G13), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(KEYINPUT68), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n273), .B1(new_n280), .B2(G238), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT13), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n265), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n282), .B1(new_n265), .B2(new_n281), .ZN(new_n285));
  OAI21_X1  g0085(.A(G200), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XOR2_X1   g0086(.A(KEYINPUT77), .B(KEYINPUT11), .Z(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT78), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n225), .ZN(new_n290));
  INV_X1    g0090(.A(G20), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n217), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(G77), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n294), .A2(new_n201), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n290), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT72), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n277), .A2(G13), .A3(G20), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n290), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n277), .A2(G20), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n277), .A2(G13), .A3(G20), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n304), .A2(KEYINPUT72), .A3(new_n225), .A4(new_n289), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n302), .A2(G68), .A3(new_n303), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n288), .A2(new_n298), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT12), .B1(new_n301), .B2(new_n213), .ZN(new_n308));
  INV_X1    g0108(.A(G13), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G1), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n310), .A2(KEYINPUT12), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n308), .B1(new_n292), .B2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n299), .A2(new_n306), .A3(new_n307), .A4(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n265), .A2(new_n281), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(G190), .A3(new_n283), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n286), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(G169), .B1(new_n284), .B2(new_n285), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT14), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n316), .A2(G179), .A3(new_n283), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT14), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n323), .B(G169), .C1(new_n284), .C2(new_n285), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n319), .B1(new_n325), .B2(new_n313), .ZN(new_n326));
  NOR2_X1   g0126(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT8), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G58), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(new_n291), .A3(G33), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT69), .ZN(new_n333));
  NOR3_X1   g0133(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(new_n291), .ZN(new_n335));
  OAI211_X1 g0135(.A(KEYINPUT69), .B(G20), .C1(new_n203), .C2(G68), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n293), .A2(G150), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n332), .A2(new_n335), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n290), .ZN(new_n339));
  INV_X1    g0139(.A(new_n290), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(KEYINPUT70), .A3(new_n304), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT70), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n301), .B2(new_n290), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n341), .A2(new_n343), .A3(G50), .A4(new_n303), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n301), .A2(new_n201), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n339), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT9), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n252), .A2(new_n254), .A3(G222), .A4(new_n255), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n252), .A2(new_n254), .A3(G223), .A4(G1698), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(new_n350), .C1(new_n296), .C2(new_n258), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n264), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n276), .A2(KEYINPUT68), .A3(new_n278), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT68), .B1(new_n276), .B2(new_n278), .ZN(new_n354));
  OAI21_X1  g0154(.A(G226), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n352), .A2(G190), .A3(new_n272), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n272), .A3(new_n355), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n359), .A2(KEYINPUT74), .A3(G200), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT74), .B1(new_n359), .B2(G200), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n348), .B(new_n358), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n339), .A2(KEYINPUT9), .A3(new_n344), .A4(new_n345), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT73), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n327), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT73), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n363), .B(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n361), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n359), .A2(KEYINPUT74), .A3(G200), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n356), .A2(new_n357), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n347), .B2(new_n346), .ZN(new_n372));
  INV_X1    g0172(.A(new_n327), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n367), .A2(new_n370), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n365), .A2(new_n374), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n331), .A2(new_n293), .B1(G20), .B2(G77), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n295), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n290), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n302), .A2(G77), .A3(new_n303), .A4(new_n305), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n301), .A2(new_n296), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n252), .A2(new_n254), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G107), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n252), .A2(new_n254), .A3(G232), .A4(new_n255), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n252), .A2(new_n254), .A3(G238), .A4(G1698), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT71), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT71), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n385), .A2(new_n390), .A3(new_n386), .A4(new_n387), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n264), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n273), .B1(new_n280), .B2(G244), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(G190), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(G244), .B1(new_n353), .B2(new_n354), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n272), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n276), .B1(new_n388), .B2(KEYINPUT71), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n396), .B1(new_n391), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n383), .B(new_n394), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G179), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n392), .A2(new_n401), .A3(new_n393), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(new_n382), .C1(new_n398), .C2(G169), .ZN(new_n403));
  INV_X1    g0203(.A(G169), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n359), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(new_n346), .C1(G179), .C2(new_n359), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n400), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n326), .A2(new_n375), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n331), .A2(new_n301), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n341), .A2(new_n343), .A3(new_n303), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(new_n331), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n228), .B1(new_n217), .B2(G58), .ZN(new_n412));
  INV_X1    g0212(.A(G159), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n412), .A2(new_n291), .B1(new_n413), .B2(new_n294), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n258), .B2(G20), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n384), .A2(KEYINPUT7), .A3(new_n291), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n213), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n340), .B1(new_n419), .B2(KEYINPUT16), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT64), .B(G68), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n416), .B2(new_n417), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n414), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n411), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n252), .A2(new_n254), .A3(G226), .A4(G1698), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n252), .A2(new_n254), .A3(G223), .A4(new_n255), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G87), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n264), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n264), .A2(new_n271), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n431), .A2(G232), .B1(new_n268), .B2(new_n271), .ZN(new_n432));
  INV_X1    g0232(.A(G190), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT80), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n430), .A2(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n399), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT80), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n430), .A2(new_n432), .A3(new_n438), .A4(new_n433), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT17), .B1(new_n425), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n416), .A2(new_n417), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G68), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n229), .B1(new_n422), .B2(new_n202), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n444), .A2(G20), .B1(G159), .B2(new_n293), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n445), .A3(KEYINPUT16), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n424), .A3(new_n290), .ZN(new_n447));
  INV_X1    g0247(.A(new_n411), .ZN(new_n448));
  AND4_X1   g0248(.A1(KEYINPUT17), .A2(new_n440), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n441), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT18), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n436), .A2(G169), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n401), .B2(new_n436), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n451), .B1(new_n425), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n447), .A2(new_n448), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(KEYINPUT18), .A3(new_n453), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(KEYINPUT79), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n459), .B(new_n451), .C1(new_n425), .C2(new_n454), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n450), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT81), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT81), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n450), .A2(new_n458), .A3(new_n463), .A4(new_n460), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n408), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n293), .A2(G77), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT6), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n467), .A2(new_n205), .A3(G107), .ZN(new_n468));
  XNOR2_X1  g0268(.A(G97), .B(G107), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n466), .B1(new_n470), .B2(new_n291), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n206), .B1(new_n416), .B2(new_n417), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n290), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n304), .A2(G97), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT82), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n277), .A2(G33), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n340), .A2(new_n475), .A3(new_n304), .A4(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n304), .A2(new_n476), .A3(new_n225), .A4(new_n289), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT82), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n474), .B1(new_n480), .B2(G97), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n252), .A2(new_n254), .A3(G244), .A4(new_n255), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G250), .A2(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(KEYINPUT4), .A2(G244), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(G1698), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n486), .B1(new_n258), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n264), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n270), .A2(G1), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(G257), .A3(new_n276), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT5), .B(G41), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n268), .A2(new_n499), .A3(new_n493), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n473), .B(new_n481), .C1(new_n502), .C2(new_n433), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n492), .A2(KEYINPUT83), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n276), .B1(new_n484), .B2(new_n490), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT83), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n399), .B1(new_n508), .B2(KEYINPUT84), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n505), .A2(new_n506), .ZN(new_n510));
  AOI211_X1 g0310(.A(KEYINPUT83), .B(new_n276), .C1(new_n484), .C2(new_n490), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n498), .A2(new_n500), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT84), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n503), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n252), .A2(new_n254), .A3(G244), .A4(G1698), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n252), .A2(new_n254), .A3(G238), .A4(new_n255), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G116), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n264), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n276), .A2(G274), .A3(new_n493), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n277), .A2(G45), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n276), .A2(G250), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n522), .A2(G179), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n404), .B1(new_n522), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n517), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n522), .A2(G179), .A3(new_n527), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n526), .B1(new_n521), .B2(new_n264), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(KEYINPUT85), .C1(new_n404), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n258), .A2(new_n291), .A3(G68), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n291), .B1(new_n261), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(G87), .B2(new_n207), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n535), .B1(new_n295), .B2(new_n205), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n539), .A2(new_n290), .B1(new_n301), .B2(new_n377), .ZN(new_n540));
  INV_X1    g0340(.A(new_n377), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n480), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n530), .A2(new_n533), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n399), .B1(new_n522), .B2(new_n527), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(G190), .B2(new_n532), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n480), .A2(G87), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n512), .A2(G179), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n504), .A2(new_n507), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n473), .A2(new_n481), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n502), .A2(new_n404), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n516), .A2(new_n550), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT21), .ZN(new_n557));
  INV_X1    g0357(.A(G116), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n277), .B2(G33), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n302), .A2(new_n305), .A3(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n304), .A2(G116), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n289), .A2(new_n225), .B1(G20), .B2(new_n558), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n485), .B(new_n291), .C1(G33), .C2(new_n205), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT20), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n563), .A2(KEYINPUT20), .A3(new_n564), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n560), .B(new_n562), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(G303), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n384), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n255), .A2(G264), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G257), .A2(G1698), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n252), .B(new_n254), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(new_n573), .A3(new_n264), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n497), .A2(G270), .A3(new_n276), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n500), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G169), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n557), .B1(new_n568), .B2(new_n577), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n574), .A2(new_n500), .A3(new_n575), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n567), .A2(new_n579), .A3(G179), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n567), .A2(KEYINPUT21), .A3(G169), .A4(new_n576), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(G200), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n566), .A2(new_n565), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n561), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n574), .A2(G190), .A3(new_n500), .A4(new_n575), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n582), .A2(new_n584), .A3(new_n560), .A4(new_n585), .ZN(new_n586));
  AND4_X1   g0386(.A1(new_n578), .A2(new_n580), .A3(new_n581), .A4(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n252), .A2(new_n254), .A3(new_n291), .A4(G87), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT22), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT22), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n258), .A2(new_n590), .A3(new_n291), .A4(G87), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n520), .A2(G20), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT23), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n291), .B2(G107), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n592), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n593), .B1(new_n592), .B2(new_n598), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n290), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n206), .B1(new_n477), .B2(new_n479), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n301), .A2(new_n206), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n604), .B(KEYINPUT25), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n497), .A2(G264), .A3(new_n276), .ZN(new_n607));
  INV_X1    g0407(.A(G294), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n251), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(G250), .A2(G1698), .ZN(new_n610));
  INV_X1    g0410(.A(G257), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n610), .B1(new_n611), .B2(G1698), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n609), .B1(new_n612), .B2(new_n258), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n500), .B(new_n607), .C1(new_n613), .C2(new_n276), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT86), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n611), .A2(G1698), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(G250), .B2(G1698), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n618), .A2(new_n384), .B1(new_n251), .B2(new_n608), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n264), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n620), .A2(KEYINPUT86), .A3(new_n500), .A4(new_n607), .ZN(new_n621));
  AOI21_X1  g0421(.A(G190), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n614), .A2(new_n399), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n602), .B(new_n606), .C1(new_n622), .C2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n616), .A2(G169), .A3(new_n621), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n499), .A2(new_n493), .B1(new_n226), .B2(new_n267), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n619), .A2(new_n264), .B1(new_n627), .B2(G264), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(KEYINPUT87), .A3(G179), .A4(new_n500), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT87), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n614), .B2(new_n401), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n592), .A2(new_n598), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT24), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n340), .B1(new_n634), .B2(new_n599), .ZN(new_n635));
  INV_X1    g0435(.A(new_n606), .ZN(new_n636));
  OAI22_X1  g0436(.A1(new_n626), .A2(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n587), .A2(new_n625), .A3(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n465), .A2(new_n556), .A3(new_n638), .ZN(G372));
  INV_X1    g0439(.A(KEYINPUT90), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n403), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n318), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n324), .A2(new_n322), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n316), .A2(new_n283), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n323), .B1(new_n644), .B2(G169), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n313), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n441), .B(new_n449), .C1(new_n642), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n455), .A2(new_n457), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n375), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n406), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n465), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n555), .A2(new_n544), .A3(new_n549), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT26), .ZN(new_n655));
  INV_X1    g0455(.A(new_n553), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n552), .A2(new_n554), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n531), .B1(new_n404), .B2(new_n532), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n546), .A2(new_n548), .B1(new_n661), .B2(new_n543), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n552), .A2(new_n554), .A3(KEYINPUT89), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n659), .A2(new_n660), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n661), .A2(new_n543), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n655), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n581), .A2(new_n580), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n575), .A2(new_n500), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n404), .B1(new_n668), .B2(new_n574), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT21), .B1(new_n669), .B2(new_n567), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n637), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n616), .A2(new_n621), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n433), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n623), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n635), .A2(new_n636), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n510), .A2(new_n511), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n678), .A2(new_n551), .B1(new_n404), .B2(new_n502), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n676), .A2(new_n677), .B1(new_n679), .B2(new_n553), .ZN(new_n680));
  INV_X1    g0480(.A(new_n503), .ZN(new_n681));
  OAI21_X1  g0481(.A(G200), .B1(new_n513), .B2(new_n514), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n508), .A2(KEYINPUT84), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n680), .A2(new_n684), .A3(new_n662), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n673), .B1(new_n685), .B2(KEYINPUT88), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT88), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n680), .A2(new_n684), .A3(new_n687), .A4(new_n662), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n666), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n652), .B1(new_n653), .B2(new_n689), .ZN(G369));
  NAND2_X1  g0490(.A1(new_n310), .A2(new_n291), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(G213), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n567), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n587), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n671), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  INV_X1    g0500(.A(new_n696), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT91), .B1(new_n677), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT91), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n703), .B(new_n696), .C1(new_n635), .C2(new_n636), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n702), .A2(new_n704), .A3(new_n625), .A4(new_n637), .ZN(new_n705));
  INV_X1    g0505(.A(new_n637), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n696), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n700), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n671), .A2(new_n696), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n705), .A2(new_n712), .B1(new_n637), .B2(new_n696), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n210), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(G87), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n205), .A3(new_n206), .A4(new_n558), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n717), .A2(new_n719), .A3(new_n277), .ZN(new_n720));
  INV_X1    g0520(.A(new_n230), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n717), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT28), .Z(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n689), .B2(new_n696), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n654), .A2(new_n660), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n659), .A2(KEYINPUT26), .A3(new_n662), .A4(new_n663), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n680), .A2(new_n672), .A3(new_n684), .A4(new_n662), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n729), .A3(new_n665), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(KEYINPUT29), .A3(new_n701), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n725), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n522), .A2(new_n527), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n614), .A2(new_n576), .A3(new_n401), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n508), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n733), .A2(new_n576), .A3(new_n401), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n628), .A2(new_n492), .A3(new_n501), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT30), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n579), .A2(G179), .A3(new_n532), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n628), .A2(new_n492), .A3(new_n501), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n735), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n696), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n696), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n661), .A2(new_n517), .B1(new_n540), .B2(new_n542), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n748), .A2(new_n533), .B1(new_n548), .B2(new_n546), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n684), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n587), .A2(new_n625), .A3(new_n637), .A4(new_n701), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n746), .B(new_n747), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n732), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n723), .B1(new_n756), .B2(G1), .ZN(G364));
  INV_X1    g0557(.A(new_n700), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n309), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n277), .B1(new_n759), .B2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OR3_X1    g0561(.A1(new_n717), .A2(new_n761), .A3(KEYINPUT92), .ZN(new_n762));
  OAI21_X1  g0562(.A(KEYINPUT92), .B1(new_n717), .B2(new_n761), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n758), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G330), .B2(new_n699), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n225), .B1(G20), .B2(new_n404), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n716), .A2(new_n258), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G45), .B2(new_n230), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT93), .Z(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n246), .B2(new_n270), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n716), .A2(new_n384), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n778), .A2(G355), .B1(new_n558), .B2(new_n716), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n773), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n771), .ZN(new_n781));
  NAND2_X1  g0581(.A1(G20), .A2(G179), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n782), .A2(new_n433), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G322), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n782), .A2(G190), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n384), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n291), .A2(G179), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(new_n433), .A3(new_n399), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n786), .B(new_n790), .C1(G329), .C2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT94), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G303), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n433), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n291), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n782), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n801), .A2(G190), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n800), .A2(G294), .B1(new_n803), .B2(G326), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n791), .A2(new_n433), .A3(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n801), .A2(new_n433), .A3(G200), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G283), .A2(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n794), .A2(new_n797), .A3(new_n804), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n792), .A2(new_n413), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT32), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n718), .A2(new_n795), .B1(new_n805), .B2(new_n206), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G50), .B2(new_n803), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n258), .B1(new_n784), .B2(new_n202), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G77), .B2(new_n787), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n799), .A2(new_n205), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G68), .B2(new_n808), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n813), .A2(new_n815), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n781), .B1(new_n811), .B2(new_n820), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n780), .A2(new_n821), .A3(new_n764), .ZN(new_n822));
  INV_X1    g0622(.A(new_n770), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n699), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n767), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  NAND2_X1  g0626(.A1(new_n382), .A2(new_n696), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n400), .A2(new_n403), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n827), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(new_n641), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n689), .B2(new_n696), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n828), .A2(new_n696), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n832), .B1(new_n689), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n765), .B1(new_n835), .B2(new_n754), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n754), .B2(new_n835), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n771), .A2(new_n768), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n765), .B1(G77), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT95), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G143), .A2(new_n783), .B1(new_n787), .B2(G159), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  INV_X1    g0643(.A(G150), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n842), .B1(new_n843), .B2(new_n802), .C1(new_n844), .C2(new_n807), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT34), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n258), .B1(new_n792), .B2(new_n848), .C1(new_n213), .C2(new_n805), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G58), .B2(new_n800), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n796), .A2(G50), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n845), .A2(new_n846), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n784), .A2(new_n608), .B1(new_n792), .B2(new_n789), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n258), .B(new_n855), .C1(G116), .C2(new_n787), .ZN(new_n856));
  INV_X1    g0656(.A(G283), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n805), .A2(new_n718), .B1(new_n807), .B2(new_n857), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n818), .B(new_n858), .C1(G303), .C2(new_n803), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n796), .A2(G107), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n856), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n854), .B1(KEYINPUT96), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(KEYINPUT96), .B2(new_n861), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n841), .B1(new_n863), .B2(new_n771), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n403), .A2(KEYINPUT90), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n403), .A2(KEYINPUT90), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(new_n866), .A3(new_n830), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n828), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n864), .B1(new_n868), .B2(new_n769), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n837), .A2(new_n869), .ZN(G384));
  NOR2_X1   g0670(.A1(new_n759), .A2(new_n277), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n421), .B1(new_n414), .B2(new_n418), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n446), .A2(new_n872), .A3(new_n290), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n448), .ZN(new_n874));
  INV_X1    g0674(.A(new_n694), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT98), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT98), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n877), .B(new_n694), .C1(new_n873), .C2(new_n448), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n461), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n456), .B1(new_n453), .B2(new_n875), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n440), .A2(new_n447), .A3(new_n448), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n874), .A2(new_n453), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n883), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n886), .A2(new_n876), .A3(new_n878), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n884), .B1(new_n887), .B2(new_n882), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n753), .A2(new_n868), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n313), .A2(new_n696), .ZN(new_n895));
  INV_X1    g0695(.A(new_n643), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n321), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n326), .B2(new_n895), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT40), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n881), .A2(new_n883), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(new_n882), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n456), .A2(new_n875), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n450), .B2(new_n648), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n890), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n892), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT40), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n894), .A2(new_n898), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n900), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n465), .A2(new_n753), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(G330), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n909), .A2(new_n910), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n897), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n646), .A2(new_n318), .A3(new_n895), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n662), .A2(new_n625), .A3(new_n750), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT88), .B1(new_n920), .B2(new_n516), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n688), .A3(new_n672), .ZN(new_n922));
  INV_X1    g0722(.A(new_n666), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n834), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n403), .A2(new_n696), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n927), .A2(new_n893), .B1(new_n649), .B2(new_n694), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n906), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n325), .A2(new_n313), .A3(new_n701), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n725), .A2(KEYINPUT99), .A3(new_n465), .A4(new_n731), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT99), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n462), .A2(new_n464), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n326), .A2(new_n375), .A3(new_n407), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(new_n731), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n922), .A2(new_n923), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT29), .B1(new_n941), .B2(new_n701), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n937), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n651), .B1(new_n936), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n935), .B(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n871), .B1(new_n916), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n916), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n227), .A2(new_n558), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n470), .B(KEYINPUT97), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT35), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n951), .B2(new_n950), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT36), .Z(new_n954));
  OAI211_X1 g0754(.A(new_n721), .B(G77), .C1(new_n202), .C2(new_n422), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(G50), .B2(new_n213), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(G1), .A3(new_n309), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n947), .A2(new_n954), .A3(new_n957), .ZN(G367));
  OAI211_X1 g0758(.A(new_n684), .B(new_n750), .C1(new_n656), .C2(new_n701), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n659), .A2(new_n663), .A3(new_n696), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n705), .A2(new_n712), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n962), .A2(new_n964), .A3(KEYINPUT42), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT42), .B1(new_n962), .B2(new_n964), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n555), .B1(new_n961), .B2(new_n706), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n965), .B(new_n966), .C1(new_n696), .C2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT100), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n548), .A2(new_n701), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n662), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n665), .B2(new_n971), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n968), .A2(new_n969), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n969), .B1(new_n968), .B2(new_n974), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n976), .A2(new_n977), .B1(new_n710), .B2(new_n962), .ZN(new_n978));
  INV_X1    g0778(.A(new_n977), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n710), .A2(new_n962), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(new_n980), .A3(new_n975), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n978), .A2(new_n981), .A3(new_n983), .ZN(new_n986));
  XNOR2_X1  g0786(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n717), .B(new_n987), .Z(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n705), .A2(new_n707), .A3(new_n712), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n964), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(new_n758), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n756), .A2(KEYINPUT104), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT103), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n714), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT45), .B1(new_n714), .B2(new_n961), .ZN(new_n996));
  XNOR2_X1  g0796(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n714), .A2(new_n961), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n997), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n962), .B2(new_n713), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n995), .A2(new_n996), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n994), .B1(new_n1001), .B2(new_n709), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n709), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n732), .A2(new_n992), .A3(new_n754), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT104), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1001), .A2(new_n994), .A3(new_n709), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n993), .A2(new_n1004), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n989), .B1(new_n1009), .B2(new_n756), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n985), .B(new_n986), .C1(new_n1010), .C2(new_n761), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n774), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n772), .B1(new_n210), .B2(new_n377), .C1(new_n240), .C2(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n765), .A2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n558), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n796), .A2(G116), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1015), .B1(new_n1016), .B2(KEYINPUT46), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n800), .A2(G107), .B1(new_n803), .B2(G311), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G97), .A2(new_n806), .B1(new_n808), .B2(G294), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n258), .B1(G303), .B2(new_n783), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n793), .A2(G317), .B1(G283), .B2(new_n787), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n800), .A2(G68), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n202), .B2(new_n795), .C1(new_n413), .C2(new_n807), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G77), .A2(new_n806), .B1(new_n803), .B2(G143), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n384), .B1(new_n793), .B2(G137), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G50), .A2(new_n787), .B1(new_n783), .B2(G150), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1017), .A2(new_n1022), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n1030));
  XOR2_X1   g0830(.A(new_n1029), .B(new_n1030), .Z(new_n1031));
  OAI221_X1 g0831(.A(new_n1014), .B1(new_n973), .B2(new_n823), .C1(new_n781), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1011), .A2(new_n1032), .ZN(G387));
  INV_X1    g0833(.A(new_n992), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n755), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(new_n717), .A3(new_n1005), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n270), .B1(new_n213), .B2(new_n296), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT106), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1037), .B1(new_n719), .B2(new_n1038), .ZN(new_n1039));
  AND3_X1   g0839(.A1(new_n331), .A2(KEYINPUT50), .A3(new_n201), .ZN(new_n1040));
  AOI21_X1  g0840(.A(KEYINPUT50), .B1(new_n331), .B2(new_n201), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1039), .B1(new_n1038), .B2(new_n719), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n774), .B(new_n1042), .C1(new_n237), .C2(new_n270), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n778), .A2(new_n719), .B1(new_n206), .B2(new_n716), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT107), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(KEYINPUT107), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n772), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n765), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G303), .A2(new_n787), .B1(new_n783), .B2(G317), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n789), .B2(new_n807), .C1(new_n785), .C2(new_n802), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT48), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n795), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n800), .A2(G283), .B1(new_n1055), .B2(G294), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT108), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT49), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n805), .A2(new_n558), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n258), .B(new_n1062), .C1(G326), .C2(new_n793), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n788), .A2(new_n213), .B1(new_n792), .B2(new_n844), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n384), .B(new_n1065), .C1(G50), .C2(new_n783), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1055), .A2(G77), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n800), .A2(new_n541), .B1(new_n808), .B2(new_n331), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G97), .A2(new_n806), .B1(new_n803), .B2(G159), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n781), .B1(new_n1064), .B2(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1049), .B(new_n1071), .C1(new_n708), .C2(new_n770), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n761), .B2(new_n992), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1036), .A2(new_n1073), .ZN(G393));
  OR2_X1    g0874(.A1(new_n1001), .A2(new_n709), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n761), .A3(new_n1003), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n784), .A2(new_n413), .B1(new_n802), .B2(new_n844), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT51), .Z(new_n1078));
  INV_X1    g0878(.A(G143), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n795), .A2(new_n422), .B1(new_n792), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT109), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n384), .B1(new_n787), .B2(new_n331), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n718), .B2(new_n805), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n799), .A2(new_n296), .B1(new_n807), .B2(new_n201), .ZN(new_n1084));
  OR4_X1    g0884(.A1(new_n1078), .A2(new_n1081), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT110), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n803), .A2(G317), .B1(G311), .B2(new_n783), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT52), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n384), .B1(new_n792), .B2(new_n785), .C1(new_n788), .C2(new_n608), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n805), .A2(new_n206), .B1(new_n807), .B2(new_n569), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n799), .A2(new_n558), .B1(new_n795), .B2(new_n857), .ZN(new_n1092));
  OR3_X1    g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1087), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n771), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n249), .A2(new_n774), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n773), .B1(G97), .B2(new_n716), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n764), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1096), .B(new_n1099), .C1(new_n961), .C2(new_n823), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1076), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n717), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1075), .A2(new_n1003), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n1005), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1101), .B1(new_n1104), .B2(new_n1009), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(G390));
  NAND3_X1  g0906(.A1(new_n753), .A2(G330), .A3(new_n868), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(new_n898), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n930), .A2(new_n931), .B1(new_n932), .B2(new_n926), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n892), .A2(new_n905), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n730), .A2(new_n701), .A3(new_n868), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n925), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n898), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1110), .A2(new_n1113), .A3(new_n933), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1108), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n926), .A2(new_n932), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT38), .B1(new_n880), .B2(new_n888), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1117), .A2(new_n1118), .A3(new_n929), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT39), .B1(new_n892), .B2(new_n905), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1116), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n556), .A2(new_n638), .A3(new_n701), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n747), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT31), .B1(new_n743), .B2(new_n696), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n831), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1126), .A2(G330), .A3(new_n919), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n932), .B(new_n906), .C1(new_n1128), .C2(new_n898), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1121), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1115), .A2(new_n761), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT111), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT111), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1115), .A2(new_n1130), .A3(new_n1133), .A4(new_n761), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n936), .A2(new_n943), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1112), .B1(new_n689), .B2(new_n834), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n919), .B1(new_n1126), .B2(G330), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n1108), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1107), .A2(new_n898), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1127), .A2(new_n1140), .A3(new_n1112), .A4(new_n1111), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n465), .A2(G330), .A3(new_n753), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1136), .A2(new_n1142), .A3(new_n652), .A4(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(new_n1115), .A3(new_n1130), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1109), .A2(new_n1108), .A3(new_n1114), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1127), .B1(new_n1121), .B2(new_n1129), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1144), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1146), .A2(new_n1149), .A3(new_n717), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n768), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n765), .B1(new_n331), .B2(new_n839), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n258), .B1(new_n796), .B2(G87), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT114), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n799), .A2(new_n296), .B1(new_n805), .B2(new_n213), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n206), .A2(new_n807), .B1(new_n802), .B2(new_n857), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n793), .A2(G294), .B1(G97), .B2(new_n787), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n558), .C2(new_n784), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n788), .A2(new_n1160), .B1(new_n807), .B2(new_n843), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT112), .Z(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n258), .B1(new_n792), .B2(new_n1163), .C1(new_n799), .C2(new_n413), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G50), .B2(new_n806), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n795), .A2(new_n844), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT53), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1162), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n803), .A2(G128), .B1(G132), .B2(new_n783), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT113), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n1154), .A2(new_n1159), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1152), .B1(new_n1171), .B2(new_n771), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1151), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1135), .A2(new_n1150), .A3(new_n1173), .ZN(G378));
  INV_X1    g0974(.A(KEYINPUT119), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n899), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n907), .ZN(new_n1177));
  XOR2_X1   g0977(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n365), .A2(new_n374), .A3(new_n406), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n346), .A2(new_n875), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT118), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n365), .A2(new_n374), .A3(new_n406), .A4(new_n1181), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1184), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1179), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT118), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n1178), .A3(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n913), .B1(new_n908), .B2(new_n906), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1177), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1193), .B1(new_n1177), .B2(new_n1194), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1175), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n935), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1126), .A2(KEYINPUT40), .A3(new_n919), .ZN(new_n1200));
  OAI21_X1  g1000(.A(G330), .B1(new_n1110), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1199), .B1(new_n900), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1177), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n928), .A2(new_n934), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1175), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1198), .A2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n938), .A2(new_n731), .A3(new_n939), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT99), .B1(new_n1208), .B2(new_n725), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n940), .A2(new_n942), .A3(new_n937), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n652), .B(new_n1143), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1115), .A2(new_n1130), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1142), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1211), .B1(new_n1217), .B2(new_n1142), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n935), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1202), .A2(new_n1205), .A3(new_n1203), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(KEYINPUT57), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n717), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1216), .A2(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n784), .A2(new_n206), .B1(new_n792), .B2(new_n857), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1023), .B1(new_n802), .B2(new_n558), .C1(new_n205), .C2(new_n807), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n541), .C2(new_n787), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n384), .A2(new_n269), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1055), .B2(G77), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT116), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n805), .A2(new_n202), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT115), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1226), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1232));
  XOR2_X1   g1032(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1227), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n1163), .A2(new_n802), .B1(new_n807), .B2(new_n848), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G128), .A2(new_n783), .B1(new_n787), .B2(G137), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n795), .B2(new_n1160), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1237), .B(new_n1239), .C1(G150), .C2(new_n800), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n806), .A2(G159), .ZN(new_n1244));
  AOI211_X1 g1044(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  AND4_X1   g1046(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1246), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n765), .B1(G50), .B2(new_n839), .C1(new_n1247), .C2(new_n781), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1199), .B2(new_n768), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1207), .B2(new_n761), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1223), .A2(new_n1250), .ZN(G375));
  XOR2_X1   g1051(.A(new_n760), .B(KEYINPUT120), .Z(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1142), .A2(new_n1253), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n784), .A2(new_n843), .B1(new_n788), .B2(new_n844), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n384), .B(new_n1255), .C1(G128), .C2(new_n793), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n799), .A2(new_n201), .B1(new_n807), .B2(new_n1160), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G132), .B2(new_n803), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n796), .A2(G159), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1256), .A2(new_n1258), .A3(new_n1231), .A4(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n788), .A2(new_n206), .B1(new_n807), .B2(new_n558), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT121), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G303), .A2(new_n793), .B1(new_n803), .B2(G294), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n800), .A2(new_n541), .B1(new_n783), .B2(G283), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1262), .B(new_n1263), .C1(KEYINPUT123), .C2(new_n1265), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1265), .A2(KEYINPUT123), .B1(G97), .B2(new_n796), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n384), .B1(new_n805), .B2(new_n296), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(KEYINPUT122), .Z(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1260), .B1(new_n1266), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n771), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n764), .B1(new_n213), .B2(new_n838), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1272), .B(new_n1273), .C1(new_n919), .C2(new_n769), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1254), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1144), .A2(new_n988), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1142), .B1(new_n944), .B2(new_n1143), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(G381));
  NAND3_X1  g1079(.A1(new_n1036), .A2(new_n825), .A3(new_n1073), .ZN(new_n1280));
  OR4_X1    g1080(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1280), .ZN(new_n1281));
  OR4_X1    g1081(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1281), .ZN(G407));
  NAND2_X1  g1082(.A1(new_n695), .A2(G213), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(G375), .A2(G378), .A3(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(KEYINPUT124), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1280), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1288), .A2(new_n1105), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1105), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(G387), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1289), .A2(new_n1011), .A3(new_n1032), .A4(new_n1290), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(G384), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1211), .A2(KEYINPUT60), .A3(new_n1214), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT60), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1144), .A2(new_n717), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1295), .B1(new_n1299), .B2(new_n1275), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n717), .B(new_n1144), .C1(new_n1278), .C2(KEYINPUT60), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1276), .B(G384), .C1(new_n1301), .C2(new_n1296), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1283), .A2(KEYINPUT125), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1300), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1283), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(G2897), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1300), .A2(new_n1302), .A3(new_n1306), .A4(new_n1303), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(G378), .B(new_n1250), .C1(new_n1216), .C2(new_n1222), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1206), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1205), .B1(new_n1204), .B2(new_n1175), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1215), .B(new_n988), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1202), .A2(new_n1205), .A3(new_n1203), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1205), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1249), .B1(new_n1317), .B2(new_n1253), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1314), .A2(new_n1318), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1135), .A2(new_n1150), .A3(new_n1173), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1311), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1283), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT61), .B1(new_n1310), .B2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1305), .B1(new_n1311), .B2(new_n1321), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(KEYINPUT62), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1324), .A2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1328), .A2(KEYINPUT62), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1294), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1326), .A2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1322), .A2(new_n1334), .A3(new_n1283), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1338), .B1(new_n1325), .B2(new_n1339), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1337), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1328), .A2(new_n1333), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT126), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1294), .B1(new_n1325), .B2(new_n1334), .ZN(new_n1344));
  AND4_X1   g1144(.A1(KEYINPUT126), .A2(new_n1324), .A3(new_n1342), .A4(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1332), .B1(new_n1343), .B2(new_n1345), .ZN(G405));
  AOI21_X1  g1146(.A(G378), .B1(new_n1223), .B2(new_n1250), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1311), .ZN(new_n1348));
  OR3_X1    g1148(.A1(new_n1347), .A2(new_n1348), .A3(new_n1327), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1327), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1350));
  OR2_X1    g1150(.A1(new_n1294), .A2(KEYINPUT127), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1349), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  AND2_X1   g1152(.A1(new_n1294), .A2(KEYINPUT127), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(new_n1352), .B(new_n1353), .ZN(G402));
endmodule


