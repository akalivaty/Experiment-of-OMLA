//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1298, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1355, new_n1356, new_n1357;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AND2_X1   g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n214), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n207), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n210), .B1(new_n212), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G200), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT3), .B(G33), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G223), .A3(G1698), .ZN(new_n247));
  INV_X1    g0047(.A(G77), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G222), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n247), .B1(new_n248), .B2(new_n246), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  AND2_X1   g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  NOR3_X1   g0055(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT68), .B1(new_n211), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G274), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT67), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT67), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n262), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n261), .A2(new_n269), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(G226), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n245), .B1(new_n260), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n260), .A2(new_n274), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n277), .B2(G190), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n255), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n203), .A2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT70), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n282), .A2(new_n283), .B1(G150), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n203), .A2(KEYINPUT70), .A3(G20), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n281), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT71), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n267), .A2(KEYINPUT71), .A3(G13), .A4(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n281), .ZN(new_n300));
  INV_X1    g0100(.A(G20), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(G1), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(new_n202), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n300), .A2(new_n304), .B1(G50), .B2(new_n299), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n294), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT9), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n294), .A2(KEYINPUT9), .A3(new_n305), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n278), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n278), .B(new_n312), .C1(new_n308), .C2(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n276), .A2(new_n315), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n316), .B1(G179), .B2(new_n276), .C1(new_n294), .C2(new_n305), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT17), .ZN(new_n320));
  INV_X1    g0120(.A(G274), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n211), .B2(new_n257), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G41), .A2(G45), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n324), .A2(KEYINPUT67), .A3(G1), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n322), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n261), .A2(G232), .A3(new_n269), .ZN(new_n327));
  NOR2_X1   g0127(.A1(G223), .A2(G1698), .ZN(new_n328));
  INV_X1    g0128(.A(G226), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(G1698), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(new_n246), .B1(G33), .B2(G87), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n254), .B1(new_n253), .B2(new_n255), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n211), .A2(KEYINPUT68), .A3(new_n257), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n326), .B(new_n327), .C1(new_n331), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n245), .ZN(new_n336));
  INV_X1    g0136(.A(G223), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n249), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n329), .A2(G1698), .ZN(new_n339));
  AND2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  NOR2_X1   g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n338), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G87), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n259), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(new_n326), .A4(new_n327), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n336), .A2(KEYINPUT77), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT77), .B1(new_n336), .B2(new_n347), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n288), .B(KEYINPUT69), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n302), .ZN(new_n352));
  INV_X1    g0152(.A(new_n300), .ZN(new_n353));
  INV_X1    g0153(.A(new_n299), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n352), .A2(new_n353), .B1(new_n354), .B2(new_n351), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n340), .A2(new_n341), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT7), .B1(new_n356), .B2(new_n301), .ZN(new_n357));
  OR2_X1    g0157(.A1(KEYINPUT3), .A2(G33), .ZN(new_n358));
  NAND2_X1  g0158(.A1(KEYINPUT3), .A2(G33), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n358), .A2(KEYINPUT7), .A3(new_n301), .A4(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(G68), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT75), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G58), .A2(G68), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n301), .B1(new_n215), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n301), .A2(new_n291), .ZN(new_n366));
  INV_X1    g0166(.A(G159), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n363), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n364), .ZN(new_n370));
  OAI21_X1  g0170(.A(G20), .B1(new_n370), .B2(new_n201), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n284), .A2(G159), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(KEYINPUT75), .A3(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n362), .A2(KEYINPUT16), .A3(new_n369), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n280), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n358), .A2(new_n301), .A3(new_n359), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(KEYINPUT76), .A3(new_n360), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT76), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n380), .A3(new_n377), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(G68), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n369), .A2(new_n373), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT16), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n355), .B1(new_n375), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n320), .B1(new_n350), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n335), .A2(G169), .ZN(new_n388));
  INV_X1    g0188(.A(new_n327), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n259), .B2(new_n344), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(G179), .A3(new_n326), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT18), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT18), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n386), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT77), .ZN(new_n397));
  INV_X1    g0197(.A(new_n347), .ZN(new_n398));
  AOI21_X1  g0198(.A(G200), .B1(new_n390), .B2(new_n326), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n336), .A2(KEYINPUT77), .A3(new_n347), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n302), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n290), .A2(new_n403), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n404), .A2(new_n300), .B1(new_n299), .B2(new_n290), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n382), .A2(new_n384), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n214), .B1(new_n378), .B2(new_n360), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n383), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n281), .B1(new_n410), .B2(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n405), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n402), .A2(new_n412), .A3(KEYINPUT17), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n387), .A2(new_n394), .A3(new_n396), .A4(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n246), .A2(G238), .A3(G1698), .ZN(new_n416));
  INV_X1    g0216(.A(G107), .ZN(new_n417));
  INV_X1    g0217(.A(G232), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n416), .B1(new_n417), .B2(new_n246), .C1(new_n250), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n259), .ZN(new_n420));
  INV_X1    g0220(.A(G244), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n326), .C1(new_n421), .C2(new_n272), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G200), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G20), .A2(G77), .ZN(new_n424));
  INV_X1    g0224(.A(new_n292), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT15), .B(G87), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n424), .B1(new_n288), .B2(new_n366), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n427), .A2(new_n280), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n300), .A2(new_n248), .A3(new_n302), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n299), .A2(G77), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n423), .B(new_n431), .C1(new_n346), .C2(new_n422), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n422), .A2(G179), .ZN(new_n433));
  INV_X1    g0233(.A(new_n431), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n422), .A2(new_n315), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n319), .A2(new_n415), .A3(new_n432), .A4(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n299), .A2(G68), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT12), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n440), .A2(KEYINPUT73), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(KEYINPUT73), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(new_n442), .C1(new_n439), .C2(new_n438), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n425), .A2(new_n248), .B1(new_n301), .B2(G68), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n366), .A2(new_n202), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n280), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT11), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n353), .A2(G68), .A3(new_n403), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n443), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT14), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT72), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n272), .A2(new_n218), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n271), .B2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n326), .B(KEYINPUT72), .C1(new_n218), .C2(new_n272), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT13), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G97), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n418), .A2(G1698), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(G226), .B2(G1698), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n459), .B2(new_n356), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n259), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n455), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n456), .B1(new_n455), .B2(new_n461), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n450), .B(G169), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n455), .A2(new_n461), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT13), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(G179), .A3(new_n462), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n462), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n450), .B1(new_n470), .B2(G169), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n449), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n449), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(G200), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n473), .B(new_n474), .C1(new_n346), .C2(new_n470), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT74), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n472), .A2(KEYINPUT74), .A3(new_n475), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n437), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n354), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n267), .A2(G33), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n299), .A2(G116), .A3(new_n281), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n279), .A2(new_n255), .B1(G20), .B2(new_n479), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n301), .C1(G33), .C2(new_n486), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n484), .A2(KEYINPUT20), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT20), .B1(new_n484), .B2(new_n487), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT84), .ZN(new_n492));
  OR2_X1    g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n264), .A2(G1), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n495), .A2(new_n496), .B1(new_n211), .B2(new_n257), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n267), .A2(G45), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n493), .B2(new_n494), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n497), .A2(G270), .B1(new_n499), .B2(new_n322), .ZN(new_n500));
  OAI211_X1 g0300(.A(G264), .B(G1698), .C1(new_n340), .C2(new_n341), .ZN(new_n501));
  OAI211_X1 g0301(.A(G257), .B(new_n249), .C1(new_n340), .C2(new_n341), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n358), .A2(G303), .A3(new_n359), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n259), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n491), .B(new_n492), .C1(new_n507), .C2(new_n245), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n245), .B1(new_n500), .B2(new_n505), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n480), .B(new_n482), .C1(new_n489), .C2(new_n488), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT84), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(G190), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n506), .A3(G169), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n500), .A2(G179), .A3(new_n505), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n510), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n510), .A2(new_n506), .A3(KEYINPUT21), .A4(G169), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n513), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G244), .B(new_n249), .C1(new_n340), .C2(new_n341), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT4), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n485), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G250), .A2(G1698), .ZN(new_n526));
  NAND2_X1  g0326(.A1(KEYINPUT4), .A2(G244), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(G1698), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n525), .B1(new_n246), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n259), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT81), .ZN(new_n532));
  INV_X1    g0332(.A(new_n494), .ZN(new_n533));
  NOR2_X1   g0333(.A1(KEYINPUT5), .A2(G41), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n496), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(G257), .A3(new_n261), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n499), .A2(new_n322), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n334), .B1(new_n524), .B2(new_n529), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(new_n537), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT81), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(G190), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n531), .A2(new_n538), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G200), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n354), .A2(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n353), .A2(new_n481), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(G97), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT6), .ZN(new_n551));
  AND2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  NOR2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT78), .ZN(new_n555));
  NAND2_X1  g0355(.A1(KEYINPUT6), .A2(G97), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(G107), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n417), .A2(KEYINPUT78), .A3(KEYINPUT6), .A4(G97), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT79), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n554), .A2(new_n557), .A3(KEYINPUT79), .A4(new_n558), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(G20), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n284), .A2(G77), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT80), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT80), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n567), .A3(new_n564), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n379), .A2(G107), .A3(new_n381), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n546), .B(new_n550), .C1(new_n570), .C2(new_n281), .ZN(new_n571));
  AOI21_X1  g0371(.A(G169), .B1(new_n539), .B2(new_n542), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n544), .A2(G179), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n569), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n565), .B2(KEYINPUT80), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n281), .B1(new_n576), .B2(new_n568), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n574), .B1(new_n577), .B2(new_n549), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT83), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n246), .A2(new_n301), .A3(G68), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT19), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n301), .B1(new_n457), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n553), .A2(new_n219), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n301), .A2(G33), .A3(G97), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT82), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n581), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n586), .B1(new_n585), .B2(new_n581), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n580), .B(new_n584), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n280), .ZN(new_n591));
  INV_X1    g0391(.A(new_n426), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n299), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n579), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  AOI211_X1 g0395(.A(KEYINPUT83), .B(new_n593), .C1(new_n590), .C2(new_n280), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n595), .A2(new_n596), .B1(new_n548), .B2(new_n426), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n496), .A2(new_n220), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n261), .A2(new_n598), .B1(new_n322), .B2(new_n496), .ZN(new_n599));
  NOR2_X1   g0399(.A1(G238), .A2(G1698), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n421), .B2(G1698), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n601), .A2(new_n246), .B1(G33), .B2(G116), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n599), .B1(new_n602), .B2(new_n334), .ZN(new_n603));
  MUX2_X1   g0403(.A(G179), .B(G169), .S(new_n603), .Z(new_n604));
  AOI21_X1  g0404(.A(G20), .B1(new_n358), .B2(new_n359), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n605), .A2(G68), .B1(new_n582), .B2(new_n583), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n585), .A2(new_n581), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT82), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n587), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n281), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT83), .B1(new_n610), .B2(new_n593), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n591), .A2(new_n579), .A3(new_n594), .ZN(new_n612));
  INV_X1    g0412(.A(new_n548), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n611), .A2(new_n612), .B1(G87), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n599), .B(G190), .C1(new_n334), .C2(new_n602), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(G200), .B2(new_n603), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n597), .A2(new_n604), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n521), .A2(new_n571), .A3(new_n578), .A4(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(G257), .B(G1698), .C1(new_n340), .C2(new_n341), .ZN(new_n620));
  OAI211_X1 g0420(.A(G250), .B(new_n249), .C1(new_n340), .C2(new_n341), .ZN(new_n621));
  NAND2_X1  g0421(.A1(G33), .A2(G294), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n259), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT85), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n497), .A2(G264), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n624), .B2(new_n626), .ZN(new_n628));
  INV_X1    g0428(.A(new_n537), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT86), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(G179), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n624), .A2(new_n626), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT85), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n634), .A2(G179), .A3(new_n537), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT86), .ZN(new_n637));
  OAI21_X1  g0437(.A(G169), .B1(new_n633), .B2(new_n629), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n632), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n246), .A2(new_n301), .A3(G87), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT22), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT22), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n605), .A2(new_n642), .A3(G87), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT24), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT23), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n301), .B2(G107), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n417), .A2(KEYINPUT23), .A3(G20), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n647), .A2(new_n648), .B1(new_n292), .B2(G116), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n644), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n645), .B1(new_n644), .B2(new_n649), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n280), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT25), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n299), .B2(G107), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n354), .A2(KEYINPUT25), .A3(new_n417), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n613), .A2(G107), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n639), .A2(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n633), .A2(G190), .A3(new_n629), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n634), .A2(new_n537), .A3(new_n635), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n245), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n657), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n619), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n478), .A2(new_n665), .ZN(G372));
  AND2_X1   g0466(.A1(new_n394), .A2(new_n396), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n472), .A2(new_n436), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n475), .A2(new_n387), .A3(new_n413), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n314), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(new_n317), .ZN(new_n672));
  INV_X1    g0472(.A(new_n478), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n597), .A2(new_n604), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n614), .A2(new_n617), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n674), .B(new_n675), .C1(new_n661), .C2(new_n657), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n520), .A2(new_n516), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(new_n658), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n571), .A2(new_n578), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT87), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n532), .B1(new_n531), .B2(new_n538), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT81), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n315), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n544), .ZN(new_n687));
  INV_X1    g0487(.A(G179), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n683), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n572), .A2(KEYINPUT87), .A3(new_n573), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT26), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n550), .B1(new_n570), .B2(new_n281), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n692), .A2(new_n693), .A3(new_n694), .A4(new_n618), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(new_n674), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n674), .A2(new_n675), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT26), .B1(new_n578), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n682), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n672), .B1(new_n673), .B2(new_n700), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT88), .Z(G369));
  INV_X1    g0502(.A(G213), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT90), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n267), .A2(new_n301), .A3(G13), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT89), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT89), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(new_n267), .A3(new_n301), .A4(G13), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n704), .B1(new_n709), .B2(KEYINPUT27), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT27), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n706), .A2(KEYINPUT90), .A3(new_n711), .A4(new_n708), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n703), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT91), .B1(new_n709), .B2(KEYINPUT27), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n709), .A2(KEYINPUT91), .A3(KEYINPUT27), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT92), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(G343), .ZN(new_n719));
  INV_X1    g0519(.A(G343), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT92), .B1(new_n716), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n491), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n677), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n513), .A2(new_n520), .A3(new_n516), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n724), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n658), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n722), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n662), .B1(new_n657), .B2(new_n639), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n722), .A2(new_n657), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n729), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n678), .A2(new_n722), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n730), .A2(new_n723), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(new_n741), .ZN(G399));
  NOR2_X1   g0542(.A1(new_n583), .A2(G116), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n208), .A2(new_n263), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(G1), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n216), .B2(new_n744), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT28), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n699), .A2(new_n723), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT29), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n693), .B1(new_n578), .B2(new_n697), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT96), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n692), .A2(KEYINPUT26), .A3(new_n694), .A4(new_n618), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT95), .ZN(new_n755));
  OAI211_X1 g0555(.A(KEYINPUT96), .B(new_n693), .C1(new_n578), .C2(new_n697), .ZN(new_n756));
  OAI21_X1  g0556(.A(KEYINPUT87), .B1(new_n572), .B2(new_n573), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n686), .A2(new_n683), .A3(new_n689), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n576), .A2(new_n568), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n549), .B1(new_n760), .B2(new_n280), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT95), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT26), .A4(new_n618), .ZN(new_n764));
  AND4_X1   g0564(.A1(new_n753), .A2(new_n755), .A3(new_n756), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n680), .A2(KEYINPUT97), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT97), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n571), .A2(new_n578), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n679), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n674), .ZN(new_n770));
  OAI211_X1 g0570(.A(KEYINPUT29), .B(new_n723), .C1(new_n765), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n750), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n726), .A2(new_n697), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n681), .A2(new_n732), .A3(new_n773), .A4(new_n723), .ZN(new_n774));
  INV_X1    g0574(.A(new_n603), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n507), .A2(new_n775), .A3(G179), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(KEYINPUT93), .B1(new_n630), .B2(new_n687), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT93), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n660), .A2(new_n779), .A3(new_n544), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n777), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT30), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n517), .A2(new_n539), .A3(new_n542), .A4(new_n775), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n634), .A2(new_n635), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n684), .A2(new_n685), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n627), .A2(new_n628), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n506), .A2(new_n688), .A3(new_n603), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(KEYINPUT30), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g0590(.A(KEYINPUT31), .B(new_n722), .C1(new_n781), .C2(new_n790), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n660), .A2(new_n779), .A3(new_n544), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n779), .B1(new_n660), .B2(new_n544), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n776), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n790), .B1(new_n794), .B2(KEYINPUT94), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT94), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n781), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n723), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n774), .B(new_n791), .C1(new_n798), .C2(KEYINPUT31), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G330), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n772), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n747), .B1(new_n801), .B2(G1), .ZN(G364));
  NAND2_X1  g0602(.A1(new_n301), .A2(G13), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n267), .B1(new_n804), .B2(G45), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n744), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n729), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(G330), .B2(new_n727), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n246), .A2(new_n208), .ZN(new_n810));
  INV_X1    g0610(.A(G355), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n811), .B1(G116), .B2(new_n208), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n243), .A2(G45), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n356), .A2(new_n208), .ZN(new_n814));
  INV_X1    g0614(.A(new_n216), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(new_n264), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n812), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(G13), .A2(G33), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(G20), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n255), .B1(G20), .B2(new_n315), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n807), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G179), .A2(G200), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n825), .A2(G20), .A3(new_n346), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G159), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT98), .B(KEYINPUT32), .ZN(new_n829));
  NOR4_X1   g0629(.A1(new_n301), .A2(new_n245), .A3(G179), .A4(G190), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n828), .A2(new_n829), .B1(G107), .B2(new_n830), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n301), .A2(new_n346), .A3(new_n245), .A4(G179), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(G87), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n301), .A2(new_n688), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G190), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n245), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n831), .B(new_n833), .C1(new_n202), .C2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n834), .A2(new_n346), .A3(new_n245), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n301), .A2(new_n688), .A3(new_n245), .A4(G190), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n246), .B1(new_n248), .B2(new_n839), .C1(new_n841), .C2(new_n214), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n835), .A2(G200), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n301), .B1(new_n825), .B2(G190), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n844), .A2(G58), .B1(G97), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n843), .B(new_n847), .C1(new_n828), .C2(new_n829), .ZN(new_n848));
  XNOR2_X1  g0648(.A(KEYINPUT99), .B(G326), .ZN(new_n849));
  INV_X1    g0649(.A(G294), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n837), .A2(new_n849), .B1(new_n850), .B2(new_n845), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT100), .ZN(new_n852));
  INV_X1    g0652(.A(G311), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n356), .B1(new_n839), .B2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(KEYINPUT33), .B(G317), .Z(new_n855));
  NOR2_X1   g0655(.A1(new_n841), .A2(new_n855), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n854), .B(new_n856), .C1(G329), .C2(new_n827), .ZN(new_n857));
  INV_X1    g0657(.A(new_n832), .ZN(new_n858));
  INV_X1    g0658(.A(G303), .ZN(new_n859));
  INV_X1    g0659(.A(new_n830), .ZN(new_n860));
  INV_X1    g0660(.A(G283), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n858), .A2(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n844), .B2(G322), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n852), .A2(new_n857), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n848), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n824), .B1(new_n865), .B2(new_n821), .ZN(new_n866));
  INV_X1    g0666(.A(new_n820), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n866), .B1(new_n727), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n809), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(G396));
  NAND2_X1  g0670(.A1(new_n722), .A2(new_n434), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n432), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n436), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n436), .A2(new_n722), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n748), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n874), .B1(new_n872), .B2(new_n436), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n677), .B1(new_n639), .B2(new_n657), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n879), .A2(new_n680), .A3(new_n676), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n695), .A2(new_n698), .A3(new_n674), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n723), .B(new_n878), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n807), .B1(new_n883), .B2(new_n800), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n800), .B2(new_n883), .ZN(new_n885));
  INV_X1    g0685(.A(new_n839), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n886), .A2(G159), .B1(new_n840), .B2(G150), .ZN(new_n887));
  INV_X1    g0687(.A(G137), .ZN(new_n888));
  INV_X1    g0688(.A(G143), .ZN(new_n889));
  INV_X1    g0689(.A(new_n844), .ZN(new_n890));
  OAI221_X1 g0690(.A(new_n887), .B1(new_n837), .B2(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT34), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n827), .A2(G132), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n830), .A2(G68), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n896), .A3(new_n246), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n858), .A2(new_n202), .B1(new_n213), .B2(new_n845), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n893), .A2(new_n894), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n860), .A2(new_n219), .B1(new_n853), .B2(new_n826), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT101), .Z(new_n901));
  AOI22_X1  g0701(.A1(new_n844), .A2(G294), .B1(G97), .B2(new_n846), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT102), .ZN(new_n903));
  OAI221_X1 g0703(.A(new_n356), .B1(new_n479), .B2(new_n839), .C1(new_n841), .C2(new_n861), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n837), .A2(new_n859), .B1(new_n417), .B2(new_n858), .ZN(new_n905));
  NOR4_X1   g0705(.A1(new_n901), .A2(new_n903), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n821), .B1(new_n899), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n821), .A2(new_n818), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n806), .B1(new_n248), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n907), .B(new_n909), .C1(new_n878), .C2(new_n819), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n885), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(G384));
  NAND3_X1  g0712(.A1(new_n478), .A2(new_n750), .A3(new_n771), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n913), .A2(new_n672), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT105), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n882), .A2(new_n875), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT103), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n407), .B1(new_n383), .B2(new_n409), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n374), .A3(new_n280), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n355), .ZN(new_n920));
  INV_X1    g0720(.A(new_n713), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n715), .A2(new_n714), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n388), .B(new_n391), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n402), .A2(new_n412), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT37), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n920), .A2(new_n923), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n350), .B2(new_n386), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n402), .A2(new_n412), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n386), .A2(new_n717), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n930), .A2(new_n925), .A3(new_n393), .A4(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n926), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n716), .B1(new_n919), .B2(new_n355), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n414), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT38), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n933), .A2(new_n935), .A3(KEYINPUT38), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n472), .A2(new_n475), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n722), .A2(new_n449), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n472), .A2(new_n475), .A3(new_n942), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n916), .A2(new_n940), .A3(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n667), .A2(new_n717), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT104), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n933), .A2(new_n935), .A3(KEYINPUT38), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT38), .B1(new_n933), .B2(new_n935), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n949), .B(KEYINPUT39), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT39), .ZN(new_n953));
  INV_X1    g0753(.A(new_n931), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n930), .A2(new_n393), .A3(new_n931), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT37), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n414), .A2(new_n954), .B1(new_n956), .B2(new_n932), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n939), .B(new_n953), .C1(KEYINPUT38), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n949), .B1(new_n940), .B2(KEYINPUT39), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n472), .A2(new_n722), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n947), .B(new_n948), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n915), .B(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n785), .A2(new_n789), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n781), .B2(new_n796), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n794), .A2(KEYINPUT94), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n722), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT31), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(KEYINPUT31), .B(new_n722), .C1(new_n966), .C2(new_n967), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n774), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n939), .B1(new_n957), .B2(KEYINPUT38), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n876), .B1(new_n944), .B2(new_n945), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT40), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT40), .B1(new_n938), .B2(new_n939), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(new_n972), .A3(new_n974), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n478), .A2(new_n972), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n979), .A2(new_n980), .ZN(new_n983));
  INV_X1    g0783(.A(G330), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n964), .A2(new_n985), .B1(new_n267), .B2(new_n804), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n964), .B2(new_n985), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n212), .A2(new_n479), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n561), .A2(new_n562), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT35), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n990), .B2(new_n989), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT36), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n815), .A2(G77), .A3(new_n364), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n202), .A2(G68), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n267), .B(G13), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n987), .A2(new_n993), .A3(new_n996), .ZN(G367));
  INV_X1    g0797(.A(KEYINPUT43), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n723), .A2(new_n614), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(new_n697), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT106), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n1001), .B2(new_n1000), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(KEYINPUT43), .B2(new_n1000), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n766), .B(new_n768), .C1(new_n761), .C2(new_n723), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n762), .A2(new_n722), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1007), .A2(new_n732), .A3(new_n737), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT42), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n730), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n722), .B1(new_n1010), .B2(new_n578), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1004), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n736), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT42), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1008), .B(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1011), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n1016), .A3(new_n1003), .ZN(new_n1017));
  AND3_X1   g0817(.A1(new_n1012), .A2(new_n1013), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1013), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n744), .B(KEYINPUT41), .ZN(new_n1021));
  AND4_X1   g0821(.A1(KEYINPUT45), .A2(new_n1007), .A3(new_n739), .A4(new_n738), .ZN(new_n1022));
  AOI21_X1  g0822(.A(KEYINPUT45), .B1(new_n1007), .B2(new_n741), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT44), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(KEYINPUT107), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1005), .A2(new_n740), .A3(new_n1006), .A4(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1025), .A2(KEYINPUT107), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1027), .B(new_n1028), .Z(new_n1029));
  NAND3_X1  g0829(.A1(new_n1024), .A2(new_n736), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n738), .B1(new_n735), .B2(new_n737), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n729), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n728), .B(new_n738), .C1(new_n735), .C2(new_n737), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n772), .A2(new_n1034), .A3(new_n800), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(KEYINPUT108), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT108), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n772), .A2(new_n1034), .A3(new_n1037), .A4(new_n800), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n736), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1027), .B(new_n1028), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1030), .A2(new_n1036), .A3(new_n1038), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1021), .B1(new_n1043), .B2(new_n801), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n805), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1020), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n208), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n823), .B1(new_n1047), .B2(new_n592), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n235), .A2(new_n208), .A3(new_n356), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n806), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(KEYINPUT109), .B(G317), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n841), .A2(new_n850), .B1(new_n826), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n246), .B(new_n1052), .C1(G283), .C2(new_n886), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n832), .A2(G116), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT46), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n836), .A2(G311), .B1(G107), .B2(new_n846), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n860), .A2(new_n486), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G303), .B2(new_n844), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT110), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n837), .A2(new_n889), .B1(new_n213), .B2(new_n858), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G150), .B2(new_n844), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n839), .A2(new_n202), .B1(new_n826), .B2(new_n888), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n356), .B(new_n1063), .C1(G159), .C2(new_n840), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n846), .A2(G68), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n830), .A2(G77), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1060), .A2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n821), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1050), .B1(new_n1000), .B2(new_n867), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1046), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT112), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(G387));
  NAND3_X1  g0876(.A1(new_n731), .A2(new_n734), .A3(new_n820), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n810), .A2(new_n743), .B1(G107), .B2(new_n208), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n232), .A2(G45), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n743), .ZN(new_n1080));
  AOI211_X1 g0880(.A(G45), .B(new_n1080), .C1(G68), .C2(G77), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n288), .A2(G50), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT50), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n814), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1078), .B1(new_n1079), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n807), .B1(new_n1085), .B2(new_n823), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n886), .A2(G303), .B1(new_n840), .B2(G311), .ZN(new_n1087));
  INV_X1    g0887(.A(G322), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1087), .B1(new_n837), .B2(new_n1088), .C1(new_n890), .C2(new_n1051), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT48), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n858), .A2(new_n850), .B1(new_n861), .B2(new_n845), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(KEYINPUT49), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n356), .B1(new_n849), .B2(new_n826), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G116), .B2(new_n830), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT49), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n845), .A2(new_n426), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n858), .B2(new_n248), .C1(new_n837), .C2(new_n367), .ZN(new_n1101));
  INV_X1    g0901(.A(G150), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n246), .B1(new_n826), .B2(new_n1102), .C1(new_n839), .C2(new_n214), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1057), .B(new_n1103), .C1(G50), .C2(new_n844), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n351), .B2(new_n841), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1097), .A2(new_n1098), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1086), .B1(new_n1106), .B2(new_n821), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1034), .A2(new_n1045), .B1(new_n1077), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n801), .A2(new_n1034), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n744), .B(KEYINPUT113), .Z(new_n1110));
  NAND2_X1  g0910(.A1(new_n1035), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1108), .B1(new_n1109), .B2(new_n1111), .ZN(G393));
  NAND2_X1  g0912(.A1(new_n1030), .A2(new_n1042), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1035), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n1043), .A3(new_n1110), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT114), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1030), .A2(KEYINPUT114), .A3(new_n1042), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n1045), .A3(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G311), .A2(new_n844), .B1(new_n836), .B2(G317), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT115), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1121), .A2(KEYINPUT52), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(KEYINPUT52), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n858), .A2(new_n861), .B1(new_n860), .B2(new_n417), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n246), .B1(new_n840), .B2(G303), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1125), .B1(new_n850), .B2(new_n839), .C1(new_n1088), .C2(new_n826), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1124), .B(new_n1126), .C1(G116), .C2(new_n846), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1122), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G150), .A2(new_n836), .B1(new_n844), .B2(G159), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT51), .Z(new_n1130));
  OAI22_X1  g0930(.A1(new_n839), .A2(new_n288), .B1(new_n826), .B2(new_n889), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n356), .B(new_n1131), .C1(G50), .C2(new_n840), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n858), .A2(new_n214), .B1(new_n860), .B2(new_n219), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n845), .A2(new_n248), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1130), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1071), .B1(new_n1128), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n240), .A2(new_n208), .A3(new_n356), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n823), .B1(G97), .B2(new_n1047), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n806), .B(new_n1137), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n1007), .B2(new_n867), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1115), .A2(new_n1119), .A3(new_n1141), .ZN(G390));
  AOI22_X1  g0942(.A1(new_n665), .A2(new_n723), .B1(new_n968), .B2(new_n969), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n984), .B1(new_n1143), .B2(new_n971), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n974), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n962), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n916), .B2(new_n946), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1148), .A2(new_n959), .A3(new_n960), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n962), .B(KEYINPUT116), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n973), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n723), .B(new_n873), .C1(new_n765), .C2(new_n770), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n875), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1151), .B1(new_n1153), .B2(new_n946), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1146), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n882), .A2(new_n875), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n946), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n962), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n959), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n940), .A2(KEYINPUT39), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT104), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1151), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n674), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n571), .A2(new_n578), .A3(new_n767), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n767), .B1(new_n571), .B2(new_n578), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1164), .B1(new_n1167), .B2(new_n679), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n755), .A2(new_n753), .A3(new_n764), .A4(new_n756), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n722), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n874), .B1(new_n1170), .B2(new_n873), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1163), .B1(new_n1171), .B2(new_n1157), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n799), .A2(new_n946), .A3(G330), .A4(new_n878), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1162), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1155), .A2(new_n1174), .A3(new_n1045), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n806), .B1(new_n351), .B2(new_n908), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n837), .A2(new_n861), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1134), .B(new_n1177), .C1(G116), .C2(new_n844), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n839), .A2(new_n486), .B1(new_n826), .B2(new_n850), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n246), .B(new_n1179), .C1(G107), .C2(new_n840), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1178), .A2(new_n833), .A3(new_n896), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(G125), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n841), .A2(new_n888), .B1(new_n1182), .B2(new_n826), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT54), .B(G143), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n356), .B(new_n1183), .C1(new_n886), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n832), .A2(G150), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT53), .Z(new_n1188));
  AOI22_X1  g0988(.A1(new_n844), .A2(G132), .B1(G159), .B2(new_n846), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n836), .A2(G128), .B1(G50), .B2(new_n830), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1186), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1181), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1176), .B1(new_n1071), .B2(new_n1192), .C1(new_n1193), .C2(new_n819), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1175), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1155), .A2(new_n1174), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT117), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n799), .A2(G330), .A3(new_n878), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1144), .A2(new_n974), .B1(new_n1198), .B2(new_n1157), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n946), .B1(new_n1144), .B2(new_n878), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1152), .A2(new_n1173), .A3(new_n875), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1199), .A2(new_n1156), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n478), .A2(new_n1144), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n913), .A2(new_n672), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1197), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1110), .B1(new_n1196), .B2(new_n1205), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1196), .A2(new_n1205), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1195), .B1(new_n1206), .B2(new_n1207), .ZN(G378));
  NOR2_X1   g1008(.A1(new_n306), .A2(new_n716), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n318), .A2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n314), .B(new_n317), .C1(new_n306), .C2(new_n716), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n979), .B2(G330), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n984), .B(new_n1215), .C1(new_n976), .C2(new_n978), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n963), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n947), .A2(new_n948), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1193), .B2(new_n1147), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n972), .A2(new_n974), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1222), .A2(new_n977), .B1(new_n975), .B2(KEYINPUT40), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1215), .B1(new_n1223), .B2(new_n984), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n979), .A2(G330), .A3(new_n1216), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1221), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1219), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1215), .A2(new_n818), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n890), .A2(new_n417), .B1(new_n213), .B2(new_n860), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G116), .B2(new_n836), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n840), .A2(G97), .B1(new_n827), .B2(G283), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n356), .A2(new_n263), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n886), .B2(new_n592), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n832), .A2(G77), .B1(new_n846), .B2(G68), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1230), .A2(new_n1231), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT58), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1232), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n886), .A2(G137), .B1(new_n840), .B2(G132), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT118), .Z(new_n1239));
  AOI22_X1  g1039(.A1(new_n844), .A2(G128), .B1(new_n832), .B2(new_n1185), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n836), .A2(G125), .B1(G150), .B2(new_n846), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n830), .A2(G159), .ZN(new_n1245));
  AOI211_X1 g1045(.A(G33), .B(G41), .C1(new_n827), .C2(G124), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1236), .B(new_n1237), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT119), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1071), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n806), .B(new_n1253), .C1(new_n202), .C2(new_n908), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1227), .A2(new_n1045), .B1(new_n1228), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1155), .A2(new_n1174), .A3(new_n1202), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1204), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(KEYINPUT57), .A3(new_n1227), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1110), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT57), .B1(new_n1257), .B2(new_n1227), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1255), .B1(new_n1259), .B2(new_n1260), .ZN(G375));
  AOI21_X1  g1061(.A(new_n806), .B1(new_n214), .B2(new_n908), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n837), .A2(new_n850), .B1(new_n486), .B2(new_n858), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G283), .B2(new_n844), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n839), .A2(new_n417), .B1(new_n826), .B2(new_n859), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n246), .B(new_n1265), .C1(G116), .C2(new_n840), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1264), .A2(new_n1066), .A3(new_n1100), .A4(new_n1266), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n832), .A2(G159), .B1(new_n827), .B2(G128), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(KEYINPUT120), .Z(new_n1269));
  AOI22_X1  g1069(.A1(new_n844), .A2(G137), .B1(G58), .B2(new_n830), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n836), .A2(G132), .B1(G50), .B2(new_n846), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n840), .A2(new_n1185), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n356), .B1(new_n886), .B2(G150), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1267), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT121), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n821), .ZN(new_n1279));
  OAI221_X1 g1079(.A(new_n1262), .B1(new_n1277), .B2(new_n1279), .C1(new_n946), .C2(new_n819), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1202), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1281), .B2(new_n805), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(KEYINPUT122), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1204), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1021), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1283), .A2(new_n1288), .ZN(G381));
  INV_X1    g1089(.A(G375), .ZN(new_n1290));
  OR3_X1    g1090(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(G381), .A2(G390), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G378), .A2(KEYINPUT123), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT123), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1294), .B(new_n1195), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1075), .A2(new_n1290), .A3(new_n1292), .A4(new_n1296), .ZN(G407));
  NAND3_X1  g1097(.A1(new_n1296), .A2(new_n1290), .A3(new_n720), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(G407), .A2(G213), .A3(new_n1298), .ZN(G409));
  XNOR2_X1  g1099(.A(G393), .B(new_n869), .ZN(new_n1300));
  AND3_X1   g1100(.A1(G390), .A2(new_n1046), .A3(new_n1072), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G390), .B1(new_n1046), .B2(new_n1072), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT125), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT125), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1300), .B(new_n1305), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT127), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1301), .A2(new_n1300), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1309), .B1(new_n1075), .B2(G390), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1307), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1308), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n703), .A2(G343), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1257), .A2(new_n1286), .A3(new_n1227), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT124), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT124), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1257), .A2(new_n1227), .A3(new_n1317), .A4(new_n1286), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1316), .A2(new_n1255), .A3(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1319), .A2(new_n1293), .A3(new_n1295), .ZN(new_n1320));
  OAI211_X1 g1120(.A(G378), .B(new_n1255), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1314), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT60), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1285), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1281), .A2(new_n1284), .A3(KEYINPUT60), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1324), .A2(new_n1287), .A3(new_n1110), .A4(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1283), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n911), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1283), .A2(new_n1326), .A3(G384), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT62), .B1(new_n1322), .B2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1314), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT126), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  AOI211_X1 g1136(.A(new_n1336), .B(new_n1314), .C1(new_n1320), .C2(new_n1321), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1335), .A2(new_n1337), .ZN(new_n1338));
  AND2_X1   g1138(.A1(new_n1331), .A2(KEYINPUT62), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1332), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1314), .A2(G2897), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1330), .B(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1342), .B1(new_n1335), .B2(new_n1337), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT61), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1313), .B1(new_n1340), .B2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1338), .A2(KEYINPUT63), .A3(new_n1331), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT63), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1322), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1348), .B1(new_n1349), .B2(new_n1330), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1351));
  AOI21_X1  g1151(.A(KEYINPUT61), .B1(new_n1342), .B2(new_n1349), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1347), .A2(new_n1350), .A3(new_n1351), .A4(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1346), .A2(new_n1353), .ZN(G405));
  NAND2_X1  g1154(.A1(new_n1296), .A2(G375), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n1321), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1356), .B(new_n1330), .ZN(new_n1357));
  XNOR2_X1  g1157(.A(new_n1357), .B(new_n1351), .ZN(G402));
endmodule


