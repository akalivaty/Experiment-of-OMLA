//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G43gat), .ZN(new_n204));
  INV_X1    g003(.A(G43gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G50gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207));
  NOR3_X1   g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT86), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR3_X1   g010(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(KEYINPUT86), .ZN(new_n217));
  NAND2_X1  g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT84), .B1(new_n205), .B2(G50gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT85), .B1(new_n203), .B2(G43gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(new_n203), .A3(G43gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT85), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(new_n205), .A3(G50gat), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n221), .A2(new_n222), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT83), .B(KEYINPUT15), .Z(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n208), .B1(new_n220), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n209), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n231), .A2(KEYINPUT82), .B1(G29gat), .B2(G36gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n209), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n232), .A2(new_n208), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT17), .B1(new_n230), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT17), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n232), .A2(new_n208), .A3(new_n235), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n217), .B(new_n218), .C1(new_n211), .C2(new_n212), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(new_n227), .B2(new_n228), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n238), .B(new_n239), .C1(new_n241), .C2(new_n208), .ZN(new_n242));
  XNOR2_X1  g041(.A(G15gat), .B(G22gat), .ZN(new_n243));
  INV_X1    g042(.A(G1gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT16), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G8gat), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n246), .B(new_n247), .C1(G1gat), .C2(new_n243), .ZN(new_n248));
  INV_X1    g047(.A(G15gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G22gat), .ZN(new_n250));
  INV_X1    g049(.A(G22gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G15gat), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n245), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(G1gat), .B1(new_n250), .B2(new_n252), .ZN(new_n254));
  OAI21_X1  g053(.A(G8gat), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n237), .A2(new_n242), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n220), .A2(new_n229), .ZN(new_n259));
  INV_X1    g058(.A(new_n208), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n236), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n256), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G229gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n202), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G113gat), .B(G141gat), .Z(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(G197gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT11), .B(G169gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n257), .B1(new_n230), .B2(new_n236), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n264), .B(KEYINPUT13), .Z(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n258), .A2(KEYINPUT18), .A3(new_n264), .A4(new_n262), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n266), .A2(new_n272), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT87), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n277), .A2(new_n279), .A3(new_n276), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(new_n277), .B2(new_n276), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n256), .B1(new_n261), .B2(new_n238), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n282), .A2(new_n237), .B1(new_n261), .B2(new_n256), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT18), .B1(new_n283), .B2(new_n264), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n280), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n272), .B(KEYINPUT81), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n278), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT88), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n277), .A2(new_n276), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT87), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n277), .A2(new_n279), .A3(new_n276), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n266), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT81), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n272), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT88), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n278), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n288), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G228gat), .A2(G233gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300));
  XNOR2_X1  g099(.A(G197gat), .B(G204gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT22), .ZN(new_n302));
  NAND2_X1  g101(.A1(G211gat), .A2(G218gat), .ZN(new_n303));
  INV_X1    g102(.A(G211gat), .ZN(new_n304));
  INV_X1    g103(.A(G218gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT67), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT22), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n303), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n310), .A2(new_n301), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n300), .B1(new_n312), .B2(KEYINPUT29), .ZN(new_n313));
  XOR2_X1   g112(.A(G155gat), .B(G162gat), .Z(new_n314));
  XNOR2_X1  g113(.A(G141gat), .B(G148gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(KEYINPUT2), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(KEYINPUT68), .ZN(new_n317));
  OR2_X1    g116(.A1(KEYINPUT69), .A2(G162gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(KEYINPUT69), .A2(G162gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(G155gat), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT2), .ZN(new_n321));
  XNOR2_X1  g120(.A(G155gat), .B(G162gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n316), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n313), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n315), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n322), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT68), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n315), .B(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n314), .B1(KEYINPUT2), .B2(new_n320), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n300), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT74), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n337), .A3(new_n334), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n312), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n299), .B1(new_n325), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n312), .A2(new_n335), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n311), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n347), .A2(new_n307), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n300), .B1(new_n348), .B2(KEYINPUT29), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n349), .A2(new_n324), .B1(G228gat), .B2(G233gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n312), .A2(new_n335), .A3(KEYINPUT73), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n341), .A2(new_n343), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n352), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n342), .B1(new_n354), .B2(new_n340), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(G22gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(G50gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n353), .A2(new_n359), .A3(new_n355), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n365));
  XNOR2_X1  g164(.A(G113gat), .B(G120gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT1), .ZN(new_n367));
  XNOR2_X1  g166(.A(G127gat), .B(G134gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n367), .B(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n332), .A2(KEYINPUT4), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT4), .B1(new_n332), .B2(new_n370), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT70), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n332), .B2(new_n300), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n324), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n376));
  INV_X1    g175(.A(new_n370), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .A4(new_n333), .ZN(new_n378));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n332), .B(new_n370), .ZN(new_n383));
  INV_X1    g182(.A(new_n379), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n381), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G1gat), .B(G29gat), .ZN(new_n388));
  INV_X1    g187(.A(G85gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT0), .B(G57gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT75), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n365), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n393), .ZN(new_n395));
  NOR4_X1   g194(.A1(new_n382), .A2(new_n386), .A3(KEYINPUT76), .A4(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n379), .B1(new_n373), .B2(new_n378), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT39), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n393), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n383), .A2(new_n384), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n402), .B2(new_n399), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT40), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n312), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT66), .B(G190gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT27), .B(G183gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT28), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412));
  INV_X1    g211(.A(G169gat), .ZN(new_n413));
  INV_X1    g212(.A(G176gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n414), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT26), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n411), .B(new_n412), .C1(new_n415), .C2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n412), .B(KEYINPUT24), .ZN(new_n419));
  INV_X1    g218(.A(new_n407), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n419), .B1(new_n420), .B2(G183gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT23), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n415), .B1(new_n422), .B2(new_n416), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n421), .B(new_n423), .C1(new_n422), .C2(new_n416), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT25), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT65), .B(G169gat), .ZN(new_n426));
  OR3_X1    g225(.A1(new_n426), .A2(new_n422), .A3(G176gat), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n427), .A2(new_n423), .ZN(new_n428));
  OR2_X1    g227(.A1(G183gat), .A2(G190gat), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT25), .B1(new_n419), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n418), .A2(new_n425), .A3(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(G226gat), .A2(G233gat), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n432), .B1(KEYINPUT29), .B2(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(KEYINPUT25), .A2(new_n424), .B1(new_n428), .B2(new_n430), .ZN(new_n435));
  INV_X1    g234(.A(new_n433), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n418), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n406), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(new_n406), .A3(new_n437), .ZN(new_n440));
  XNOR2_X1  g239(.A(G8gat), .B(G36gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G64gat), .B(G92gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n440), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n443), .B1(new_n448), .B2(new_n438), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n439), .A2(KEYINPUT30), .A3(new_n440), .A4(new_n444), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n403), .A2(new_n404), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n397), .A2(new_n405), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT71), .B(KEYINPUT6), .Z(new_n454));
  NAND2_X1  g253(.A1(new_n380), .A2(new_n381), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n380), .A2(new_n385), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n381), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n454), .B1(new_n457), .B2(new_n392), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n394), .B2(new_n396), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT77), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n392), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n387), .A2(new_n462), .A3(new_n454), .ZN(new_n463));
  OR3_X1    g262(.A1(new_n448), .A2(KEYINPUT37), .A3(new_n438), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT37), .B1(new_n448), .B2(new_n438), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n464), .A2(new_n443), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT38), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n458), .B(KEYINPUT77), .C1(new_n394), .C2(new_n396), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n461), .A2(new_n463), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n445), .B1(new_n466), .B2(new_n467), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n364), .B(new_n453), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n458), .B1(new_n392), .B2(new_n457), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n463), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n363), .B1(new_n475), .B2(new_n451), .ZN(new_n476));
  NAND2_X1  g275(.A1(G227gat), .A2(G233gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n477), .B(KEYINPUT64), .Z(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n432), .A2(new_n377), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n435), .A2(new_n370), .A3(new_n418), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT32), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT34), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n480), .A2(new_n479), .A3(new_n481), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G43gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n486), .B(new_n487), .Z(new_n488));
  OAI211_X1 g287(.A(new_n485), .B(new_n488), .C1(new_n482), .C2(KEYINPUT33), .ZN(new_n489));
  INV_X1    g288(.A(new_n481), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n370), .B1(new_n435), .B2(new_n418), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT33), .ZN(new_n493));
  INV_X1    g292(.A(new_n488), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n492), .B(new_n479), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n478), .B1(new_n490), .B2(new_n491), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(KEYINPUT32), .A3(new_n497), .ZN(new_n498));
  AND4_X1   g297(.A1(new_n484), .A2(new_n489), .A3(new_n495), .A4(new_n498), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n495), .A2(new_n489), .B1(new_n484), .B2(new_n498), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n501), .B1(new_n499), .B2(new_n500), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n472), .B(new_n476), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n461), .A2(new_n463), .A3(new_n469), .ZN(new_n506));
  INV_X1    g305(.A(new_n451), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n499), .A2(new_n500), .ZN(new_n508));
  AND4_X1   g307(.A1(new_n507), .A2(new_n508), .A3(new_n361), .A4(new_n362), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT78), .B(KEYINPUT35), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n506), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT79), .ZN(new_n512));
  INV_X1    g311(.A(new_n508), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(new_n363), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(new_n474), .A3(new_n507), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT35), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT79), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n506), .A2(new_n509), .A3(new_n517), .A4(new_n510), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n512), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n298), .B1(new_n505), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521));
  INV_X1    g320(.A(G92gat), .ZN(new_n522));
  AOI22_X1  g321(.A1(KEYINPUT8), .A2(new_n521), .B1(new_n389), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT7), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(new_n389), .B2(new_n522), .ZN(new_n525));
  NAND3_X1  g324(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G99gat), .B(G106gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n237), .A2(new_n242), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G232gat), .A2(G233gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT95), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n261), .A2(new_n529), .B1(KEYINPUT41), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G190gat), .B(G218gat), .Z(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT96), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n533), .A2(KEYINPUT41), .ZN(new_n538));
  XNOR2_X1  g337(.A(G134gat), .B(G162gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n531), .A2(new_n534), .ZN(new_n542));
  INV_X1    g341(.A(new_n535), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n536), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n537), .A2(new_n544), .A3(new_n536), .A4(new_n540), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT91), .ZN(new_n550));
  INV_X1    g349(.A(G64gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(G57gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT90), .B(G57gat), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(G64gat), .ZN(new_n555));
  INV_X1    g354(.A(G71gat), .ZN(new_n556));
  INV_X1    g355(.A(G78gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(KEYINPUT9), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n550), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(KEYINPUT90), .A2(G57gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(KEYINPUT90), .A2(G57gat), .ZN(new_n563));
  OAI21_X1  g362(.A(G64gat), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n552), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n556), .B2(new_n557), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(KEYINPUT91), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT9), .ZN(new_n570));
  INV_X1    g369(.A(G57gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G64gat), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n570), .B1(new_n552), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT89), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT89), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(G71gat), .B2(G78gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n573), .A2(new_n577), .A3(new_n558), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT94), .B1(new_n569), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n581));
  AOI211_X1 g380(.A(new_n581), .B(new_n578), .C1(new_n561), .C2(new_n568), .ZN(new_n582));
  OAI211_X1 g381(.A(KEYINPUT10), .B(new_n529), .C1(new_n580), .C2(new_n582), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n555), .A2(new_n560), .A3(new_n550), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT91), .B1(new_n565), .B2(new_n567), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n579), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n530), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT10), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n578), .B1(new_n561), .B2(new_n568), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n529), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n587), .A2(new_n590), .ZN(new_n595));
  INV_X1    g394(.A(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n586), .A2(new_n581), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(G183gat), .B1(new_n610), .B2(new_n256), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT21), .B1(new_n580), .B2(new_n582), .ZN(new_n612));
  INV_X1    g411(.A(G183gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n257), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n611), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n611), .B2(new_n614), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n606), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n611), .A2(new_n614), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n615), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n611), .A2(new_n614), .A3(new_n616), .ZN(new_n622));
  INV_X1    g421(.A(new_n606), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n304), .B1(new_n586), .B2(new_n607), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n589), .A2(KEYINPUT21), .A3(G211gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629));
  NAND3_X1  g428(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n629), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n625), .B2(new_n627), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n630), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n630), .B2(new_n634), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n619), .A2(new_n624), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n619), .B2(new_n624), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n549), .B(new_n605), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n520), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n474), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n244), .ZN(G1324gat));
  INV_X1    g443(.A(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n451), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n247), .A2(KEYINPUT16), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n247), .A2(KEYINPUT16), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(KEYINPUT42), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(G8gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(KEYINPUT42), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(G1325gat));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n504), .B2(new_n502), .ZN(new_n655));
  INV_X1    g454(.A(new_n502), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(KEYINPUT97), .A3(new_n503), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n657), .A3(KEYINPUT98), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n642), .A2(new_n249), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n508), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n249), .B2(new_n664), .ZN(G1326gat));
  NOR2_X1   g464(.A1(new_n642), .A2(new_n364), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT99), .B(KEYINPUT43), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n638), .A2(new_n639), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n604), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n549), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n520), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(new_n215), .A3(new_n475), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n505), .A2(new_n519), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(new_n548), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n548), .A2(KEYINPUT101), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n546), .A2(new_n683), .A3(new_n547), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n472), .A2(new_n476), .A3(new_n658), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n685), .B(new_n686), .C1(new_n519), .C2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n287), .B(new_n672), .C1(new_n681), .C2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G29gat), .B1(new_n689), .B2(new_n474), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n678), .A2(new_n690), .ZN(G1328gat));
  NOR3_X1   g490(.A1(new_n675), .A2(G36gat), .A3(new_n507), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT46), .ZN(new_n693));
  OAI21_X1  g492(.A(G36gat), .B1(new_n689), .B2(new_n507), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1329gat));
  OAI21_X1  g494(.A(G43gat), .B1(new_n689), .B2(new_n658), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n675), .A2(G43gat), .A3(new_n513), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n696), .A2(new_n698), .A3(KEYINPUT47), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n689), .A2(new_n662), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n697), .B1(new_n700), .B2(G43gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n701), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g501(.A(new_n689), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(G50gat), .A3(new_n363), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT102), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n705), .A2(KEYINPUT102), .ZN(new_n707));
  AOI21_X1  g506(.A(G50gat), .B1(new_n676), .B2(new_n363), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n704), .A2(new_n706), .A3(new_n707), .A4(new_n709), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n689), .A2(new_n203), .A3(new_n364), .ZN(new_n711));
  OAI211_X1 g510(.A(KEYINPUT102), .B(new_n705), .C1(new_n711), .C2(new_n708), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n710), .A2(new_n712), .ZN(G1331gat));
  NAND2_X1  g512(.A1(new_n519), .A2(new_n687), .ZN(new_n714));
  INV_X1    g513(.A(new_n287), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n670), .A2(new_n548), .A3(new_n605), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT103), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n287), .B1(new_n519), .B2(new_n687), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(new_n720), .A3(new_n716), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(new_n723), .A3(new_n475), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n723), .B1(new_n722), .B2(new_n475), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n554), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n726), .ZN(new_n728));
  INV_X1    g527(.A(new_n554), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n728), .A2(new_n729), .A3(new_n724), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(G1332gat));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n732));
  NAND2_X1  g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n722), .A2(new_n732), .A3(new_n451), .A4(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n718), .A2(new_n451), .A3(new_n721), .A4(new_n733), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT105), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n735), .B1(new_n734), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(G1333gat));
  INV_X1    g539(.A(new_n662), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n722), .A2(G71gat), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(G71gat), .B1(new_n722), .B2(new_n508), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT50), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n722), .A2(new_n508), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n746), .B(new_n742), .C1(new_n747), .C2(G71gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n722), .A2(new_n363), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT106), .B(G78gat), .Z(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1335gat));
  INV_X1    g551(.A(new_n681), .ZN(new_n753));
  INV_X1    g552(.A(new_n688), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n670), .A2(new_n715), .A3(new_n604), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT107), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(new_n475), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT108), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n755), .A2(new_n760), .A3(new_n475), .A4(new_n757), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(G85gat), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n719), .A2(new_n548), .A3(new_n670), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT51), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n719), .A2(new_n765), .A3(new_n548), .A4(new_n670), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n604), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n475), .A2(new_n389), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n762), .B1(new_n767), .B2(new_n768), .ZN(G1336gat));
  OAI211_X1 g568(.A(new_n451), .B(new_n757), .C1(new_n681), .C2(new_n688), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G92gat), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n507), .A2(G92gat), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n764), .A2(new_n604), .A3(new_n766), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n771), .B(new_n775), .C1(new_n772), .C2(KEYINPUT52), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(G1337gat));
  INV_X1    g578(.A(G99gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n767), .B2(new_n513), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n755), .A2(G99gat), .A3(new_n741), .A4(new_n757), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n781), .A2(KEYINPUT110), .A3(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(G1338gat));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n363), .B(new_n757), .C1(new_n681), .C2(new_n688), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n364), .A2(G106gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n790), .B1(new_n767), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n792), .B(new_n794), .ZN(G1339gat));
  OAI21_X1  g594(.A(KEYINPUT112), .B1(new_n640), .B2(new_n287), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n619), .A2(new_n624), .ZN(new_n797));
  INV_X1    g596(.A(new_n637), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n619), .A2(new_n624), .A3(new_n637), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n548), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n801), .A2(new_n802), .A3(new_n715), .A4(new_n605), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n796), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n583), .A2(new_n596), .A3(new_n591), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n594), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n592), .A2(new_n593), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(new_n601), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n807), .A2(KEYINPUT55), .A3(new_n601), .A4(new_n809), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n812), .A2(new_n602), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n682), .A2(new_n684), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n283), .A2(new_n264), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n274), .A2(new_n275), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n270), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n278), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n812), .A2(new_n820), .A3(new_n602), .A4(new_n813), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT114), .B1(new_n685), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n604), .A2(new_n820), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n812), .A2(new_n602), .A3(new_n813), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n715), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n685), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n805), .B1(new_n829), .B2(new_n671), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(new_n514), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n474), .A2(new_n451), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT115), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n715), .A2(G113gat), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G113gat), .B1(new_n833), .B2(new_n298), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT116), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n836), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(G1340gat));
  INV_X1    g641(.A(G120gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n834), .A2(new_n843), .A3(new_n604), .ZN(new_n844));
  OAI21_X1  g643(.A(G120gat), .B1(new_n833), .B2(new_n605), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1341gat));
  INV_X1    g645(.A(new_n833), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n671), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n548), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(G134gat), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT56), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(G134gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1343gat));
  INV_X1    g653(.A(G141gat), .ZN(new_n855));
  INV_X1    g654(.A(new_n832), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n655), .B2(new_n657), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n830), .A2(new_n858), .A3(new_n363), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n825), .B1(new_n298), .B2(new_n826), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(new_n549), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n824), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n812), .A2(new_n813), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n864), .A2(new_n288), .A3(new_n297), .A4(new_n602), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n548), .B1(new_n865), .B2(new_n825), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n861), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n670), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n364), .B1(new_n868), .B2(new_n805), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n857), .B(new_n859), .C1(new_n869), .C2(new_n858), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n825), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n295), .A2(new_n296), .A3(new_n278), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n296), .B1(new_n295), .B2(new_n278), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n873), .B1(new_n876), .B2(new_n814), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT117), .B1(new_n877), .B2(new_n548), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n824), .A3(new_n862), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n804), .B1(new_n879), .B2(new_n670), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT57), .B1(new_n880), .B2(new_n364), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n881), .A2(KEYINPUT118), .A3(new_n857), .A4(new_n859), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n872), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n855), .B1(new_n883), .B2(new_n287), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n741), .A2(new_n856), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n830), .A2(new_n363), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n885), .A2(new_n886), .A3(new_n855), .A4(new_n876), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT58), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n881), .A2(new_n876), .A3(new_n857), .A4(new_n859), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G141gat), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  AND4_X1   g691(.A1(KEYINPUT119), .A2(new_n891), .A3(new_n892), .A4(new_n887), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT58), .B1(new_n890), .B2(G141gat), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT119), .B1(new_n894), .B2(new_n887), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n889), .A2(new_n896), .ZN(G1344gat));
  NAND2_X1  g696(.A1(new_n885), .A2(new_n886), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(G148gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n604), .ZN(new_n901));
  AOI211_X1 g700(.A(KEYINPUT59), .B(new_n900), .C1(new_n883), .C2(new_n604), .ZN(new_n902));
  XNOR2_X1  g701(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n822), .A2(new_n549), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n670), .B1(new_n866), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n640), .B2(new_n876), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n801), .A2(new_n298), .A3(KEYINPUT121), .A4(new_n605), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n364), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n904), .B1(new_n911), .B2(KEYINPUT57), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n830), .A2(KEYINPUT57), .A3(new_n363), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n909), .ZN(new_n914));
  INV_X1    g713(.A(new_n905), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(new_n877), .B2(new_n548), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n914), .B1(new_n916), .B2(new_n670), .ZN(new_n917));
  OAI211_X1 g716(.A(KEYINPUT122), .B(new_n858), .C1(new_n917), .C2(new_n364), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n912), .A2(new_n913), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n604), .A3(new_n857), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n903), .B1(new_n920), .B2(G148gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n901), .B1(new_n902), .B2(new_n921), .ZN(G1345gat));
  AOI21_X1  g721(.A(G155gat), .B1(new_n899), .B2(new_n671), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n872), .A2(new_n882), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n670), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n923), .B1(new_n925), .B2(G155gat), .ZN(G1346gat));
  NAND2_X1  g725(.A1(new_n318), .A2(new_n319), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n924), .A2(new_n927), .A3(new_n685), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n899), .A2(new_n548), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n927), .B2(new_n929), .ZN(G1347gat));
  NAND2_X1  g729(.A1(new_n474), .A2(new_n451), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n831), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n298), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n715), .A2(new_n426), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(G1348gat));
  NOR2_X1   g735(.A1(new_n933), .A2(new_n605), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(new_n414), .ZN(G1349gat));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n933), .A2(new_n670), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n941), .B2(G183gat), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT123), .B1(new_n940), .B2(new_n408), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n940), .A2(KEYINPUT123), .A3(new_n408), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT60), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT60), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n942), .B(new_n947), .C1(new_n943), .C2(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n933), .B2(new_n549), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n816), .A2(new_n407), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n933), .B2(new_n952), .ZN(G1351gat));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n954), .B1(new_n662), .B2(new_n932), .ZN(new_n955));
  AOI211_X1 g754(.A(KEYINPUT125), .B(new_n931), .C1(new_n660), .C2(new_n661), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n919), .A2(new_n876), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G197gat), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n830), .A2(new_n363), .A3(new_n662), .A4(new_n932), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n715), .A2(G197gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(G1352gat));
  NOR3_X1   g761(.A1(new_n960), .A2(G204gat), .A3(new_n605), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT62), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n919), .A2(new_n604), .A3(new_n957), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n919), .A2(new_n671), .A3(new_n957), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G211gat), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT63), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT63), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n971), .A3(G211gat), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n960), .A2(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT126), .B1(new_n973), .B2(new_n670), .ZN(new_n974));
  OR4_X1    g773(.A1(KEYINPUT126), .A2(new_n960), .A3(G211gat), .A4(new_n670), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n970), .A2(new_n972), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n970), .A2(new_n976), .A3(new_n979), .A4(new_n972), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1354gat));
  NAND4_X1  g780(.A1(new_n919), .A2(new_n957), .A3(G218gat), .A4(new_n548), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n305), .B1(new_n960), .B2(new_n685), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n982), .A2(new_n983), .ZN(G1355gat));
endmodule


