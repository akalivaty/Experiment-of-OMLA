//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1191, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n205), .B(new_n206), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G107), .A2(G264), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n208), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G116), .B2(G270), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G77), .A2(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n203), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n207), .B(new_n222), .C1(new_n225), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n231), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(KEYINPUT72), .ZN(new_n246));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G20), .ZN(new_n248));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  OAI21_X1  g0049(.A(KEYINPUT68), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT68), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n251), .A2(new_n247), .A3(G13), .A4(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G13), .A2(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n223), .B1(new_n254), .B2(new_n203), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G50), .A3(new_n248), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n250), .A2(new_n252), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n215), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G150), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NOR3_X1   g0069(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n267), .A2(new_n269), .B1(new_n270), .B2(new_n224), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n255), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n259), .A2(new_n261), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G222), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G223), .A2(G1698), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n223), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n280), .B(new_n282), .C1(G77), .C2(new_n276), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT67), .B1(new_n281), .B2(new_n223), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT67), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(G1), .A4(G13), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G41), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  AOI21_X1  g0090(.A(G1), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(G274), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n283), .B(new_n292), .C1(new_n216), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n259), .A2(KEYINPUT9), .A3(new_n261), .A4(new_n272), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(G200), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n275), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n246), .B1(new_n300), .B2(KEYINPUT71), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n300), .A2(new_n246), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n246), .B(KEYINPUT10), .C1(new_n300), .C2(KEYINPUT71), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n295), .A2(G179), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n295), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n273), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  AOI211_X1 g0111(.A(KEYINPUT70), .B(new_n255), .C1(new_n252), .C2(new_n250), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT70), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n253), .B2(new_n256), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n248), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n254), .A2(new_n203), .ZN(new_n318));
  OAI21_X1  g0118(.A(G77), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n269), .A2(KEYINPUT69), .ZN(new_n320));
  INV_X1    g0120(.A(new_n262), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n269), .A2(KEYINPUT69), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  XOR2_X1   g0123(.A(KEYINPUT15), .B(G87), .Z(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n264), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n256), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G77), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n260), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  NOR2_X1   g0132(.A1(KEYINPUT3), .A2(G33), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(G238), .B2(G1698), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n219), .B2(G1698), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n336), .B(new_n282), .C1(G107), .C2(new_n276), .ZN(new_n337));
  INV_X1    g0137(.A(G244), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n292), .C1(new_n338), .C2(new_n294), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(G179), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n308), .B2(new_n339), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n311), .B1(new_n331), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n260), .A2(KEYINPUT76), .A3(new_n210), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT12), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT76), .B1(new_n260), .B2(new_n210), .ZN(new_n345));
  XOR2_X1   g0145(.A(new_n344), .B(new_n345), .Z(new_n346));
  NAND2_X1  g0146(.A1(new_n317), .A2(G68), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n268), .A2(G50), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT75), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n264), .A2(G77), .B1(G20), .B2(new_n210), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n256), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  XOR2_X1   g0151(.A(new_n351), .B(KEYINPUT11), .Z(new_n352));
  NAND3_X1  g0152(.A1(new_n346), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n292), .B1(new_n294), .B2(new_n211), .ZN(new_n354));
  INV_X1    g0154(.A(new_n282), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n216), .A2(new_n277), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n276), .B(new_n356), .C1(G232), .C2(new_n277), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G97), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT73), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT73), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(G33), .A3(G97), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n355), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  OR3_X1    g0163(.A1(new_n354), .A2(KEYINPUT13), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT74), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT13), .B1(new_n354), .B2(new_n363), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n366), .A2(new_n365), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n353), .B1(G190), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n364), .A2(new_n366), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G200), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G179), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n367), .B2(new_n368), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT14), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n371), .B2(G169), .ZN(new_n378));
  AOI211_X1 g0178(.A(KEYINPUT14), .B(new_n308), .C1(new_n364), .C2(new_n366), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n353), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n339), .A2(G200), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n339), .A2(new_n296), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n328), .A2(new_n383), .A3(new_n384), .A4(new_n330), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n374), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n276), .B2(G20), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n334), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n210), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n218), .A2(new_n210), .ZN(new_n393));
  NOR2_X1   g0193(.A1(G58), .A2(G68), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n268), .A2(G159), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n388), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT7), .B1(new_n334), .B2(new_n224), .ZN(new_n399));
  NOR4_X1   g0199(.A1(new_n332), .A2(new_n333), .A3(new_n389), .A4(G20), .ZN(new_n400));
  OAI21_X1  g0200(.A(G68), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n397), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(KEYINPUT16), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n398), .A2(new_n403), .A3(new_n255), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n262), .A2(new_n316), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n258), .A2(new_n405), .B1(new_n260), .B2(new_n262), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G274), .ZN(new_n408));
  AOI211_X1 g0208(.A(new_n408), .B(new_n293), .C1(new_n284), .C2(new_n287), .ZN(new_n409));
  AOI211_X1 g0209(.A(new_n219), .B(new_n291), .C1(new_n284), .C2(new_n287), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT78), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(G226), .B(G1698), .C1(new_n332), .C2(new_n333), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT77), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n276), .A2(KEYINPUT77), .A3(G226), .A4(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n276), .A2(G223), .A3(new_n277), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G87), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n282), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n288), .A2(G232), .A3(new_n293), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT78), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n292), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n411), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n308), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n411), .A2(new_n420), .A3(new_n375), .A4(new_n423), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n407), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n427), .B(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n424), .A2(G200), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n411), .A2(new_n420), .A3(G190), .A4(new_n423), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n430), .A2(new_n406), .A3(new_n404), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n407), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n435), .A2(KEYINPUT17), .A3(new_n431), .A4(new_n430), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n434), .A2(KEYINPUT79), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT79), .B1(new_n434), .B2(new_n436), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n429), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n439), .A2(KEYINPUT80), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(KEYINPUT80), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n342), .A2(new_n387), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(G244), .B1(new_n332), .B2(new_n333), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT4), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n443), .A2(new_n444), .B1(G33), .B2(G283), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n276), .A2(KEYINPUT4), .A3(G244), .A4(new_n277), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n276), .B2(G250), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n445), .B(new_n446), .C1(new_n277), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT5), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G41), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n450), .A2(KEYINPUT84), .A3(new_n247), .A4(G45), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n288), .A2(G274), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n247), .A3(G45), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT84), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n454), .A2(new_n455), .B1(KEYINPUT5), .B2(new_n289), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n448), .A2(new_n282), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n289), .A2(KEYINPUT5), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n458), .A2(new_n459), .B1(new_n284), .B2(new_n287), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G257), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n296), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n448), .A2(new_n282), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n456), .A2(new_n288), .A3(G274), .A4(new_n451), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n463), .A2(new_n464), .A3(new_n461), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n462), .B1(new_n465), .B2(G200), .ZN(new_n466));
  OAI21_X1  g0266(.A(G107), .B1(new_n399), .B2(new_n400), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n268), .A2(G77), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(G97), .B(G107), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT82), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OR2_X1    g0275(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(G107), .A3(new_n472), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n470), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT82), .B1(new_n476), .B2(new_n472), .ZN(new_n479));
  XOR2_X1   g0279(.A(G97), .B(G107), .Z(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT83), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G107), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n473), .A2(new_n474), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n480), .B1(new_n484), .B2(new_n479), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT83), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n475), .A2(new_n470), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n469), .B1(new_n489), .B2(G20), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n490), .A2(new_n256), .ZN(new_n491));
  INV_X1    g0291(.A(G97), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n260), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n263), .A2(G1), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n257), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G97), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n466), .A2(new_n491), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n253), .A2(new_n324), .ZN(new_n498));
  INV_X1    g0298(.A(G87), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n257), .A2(new_n499), .A3(new_n494), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT19), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n224), .B1(new_n362), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n492), .A3(new_n483), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n501), .B1(new_n265), .B2(new_n492), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n276), .A2(new_n224), .A3(G68), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT85), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT85), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n276), .A2(new_n508), .A3(new_n224), .A4(G68), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n504), .A2(new_n505), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  AOI211_X1 g0310(.A(new_n498), .B(new_n500), .C1(new_n510), .C2(new_n255), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n247), .A2(new_n408), .A3(G45), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n288), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G250), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n290), .B2(G1), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G116), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n276), .B1(G244), .B2(new_n277), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G238), .A2(G1698), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n513), .A2(new_n515), .B1(new_n519), .B2(new_n282), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G190), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n282), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n288), .A2(new_n515), .A3(new_n512), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G200), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n498), .B1(new_n510), .B2(new_n255), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n495), .A2(new_n324), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n527), .A2(new_n528), .B1(new_n308), .B2(new_n524), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n520), .A2(new_n375), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n511), .A2(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n493), .B(new_n496), .C1(new_n490), .C2(new_n256), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n465), .A2(new_n375), .ZN(new_n533));
  AOI21_X1  g0333(.A(G169), .B1(new_n457), .B2(new_n461), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n224), .A2(G33), .A3(G116), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n224), .A2(G107), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT23), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n224), .B(G87), .C1(new_n332), .C2(new_n333), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n540), .A2(KEYINPUT22), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(KEYINPUT22), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n537), .B(new_n539), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT24), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n540), .B(KEYINPUT22), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(KEYINPUT24), .A3(new_n537), .A4(new_n539), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n255), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n495), .A2(G107), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n253), .A2(G107), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n550), .B(KEYINPUT25), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G250), .B(new_n277), .C1(new_n332), .C2(new_n333), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT86), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT86), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n276), .A2(new_n556), .A3(G250), .A4(new_n277), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G294), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n276), .A2(G257), .A3(G1698), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n555), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n282), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n460), .A2(G264), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n464), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT87), .B1(new_n563), .B2(G190), .ZN(new_n564));
  INV_X1    g0364(.A(G200), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n560), .A2(new_n282), .B1(new_n460), .B2(G264), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT87), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n296), .A4(new_n464), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n564), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n553), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n497), .A2(new_n531), .A3(new_n536), .A4(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n494), .ZN(new_n573));
  OAI211_X1 g0373(.A(G116), .B(new_n573), .C1(new_n312), .C2(new_n314), .ZN(new_n574));
  AOI21_X1  g0374(.A(G20), .B1(G33), .B2(G283), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(G33), .B2(new_n492), .ZN(new_n576));
  INV_X1    g0376(.A(G116), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G20), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n255), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT20), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n576), .A2(new_n255), .A3(KEYINPUT20), .A4(new_n578), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n581), .A2(new_n582), .B1(new_n260), .B2(new_n577), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n574), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n460), .A2(G270), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n277), .A2(G257), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G264), .A2(G1698), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n276), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(new_n282), .C1(G303), .C2(new_n276), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n585), .A2(new_n464), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n584), .A2(G169), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n584), .A2(KEYINPUT21), .A3(G169), .A4(new_n590), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n590), .A2(new_n375), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n584), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n563), .A2(G179), .ZN(new_n598));
  AOI21_X1  g0398(.A(G169), .B1(new_n567), .B2(new_n464), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n552), .ZN(new_n601));
  OR2_X1    g0401(.A1(new_n590), .A2(new_n296), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n590), .A2(G200), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n602), .A2(new_n583), .A3(new_n574), .A4(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n595), .A2(new_n597), .A3(new_n601), .A4(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n442), .A2(new_n572), .A3(new_n605), .ZN(G372));
  XNOR2_X1  g0406(.A(new_n427), .B(KEYINPUT18), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n331), .A2(new_n341), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n374), .A2(new_n608), .B1(new_n381), .B2(new_n380), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n434), .A2(new_n436), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT79), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n434), .A2(new_n436), .A3(KEYINPUT79), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n607), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n306), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n310), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n534), .B1(new_n375), .B2(new_n465), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n531), .A2(KEYINPUT26), .A3(new_n532), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n527), .A2(new_n528), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n524), .A2(new_n308), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n530), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n500), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n525), .A2(new_n521), .A3(new_n527), .A4(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n619), .A2(new_n532), .A3(new_n623), .A4(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT90), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n626), .B2(new_n628), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n620), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n623), .B(KEYINPUT89), .ZN(new_n633));
  INV_X1    g0433(.A(new_n572), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT88), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n600), .B2(new_n552), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n600), .A2(new_n635), .A3(new_n552), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n637), .A2(new_n595), .A3(new_n597), .A4(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n633), .B1(new_n634), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n632), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n618), .B1(new_n442), .B2(new_n642), .ZN(G369));
  NOR2_X1   g0443(.A1(new_n249), .A2(G20), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n247), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(G213), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G343), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n601), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n571), .A2(new_n601), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n552), .A2(new_n650), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n593), .A2(new_n597), .A3(new_n594), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n651), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n584), .A2(new_n650), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n656), .B(new_n659), .Z(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(G330), .A3(new_n604), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n653), .A2(new_n656), .A3(new_n651), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n638), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n651), .B1(new_n665), .B2(new_n636), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(G399));
  INV_X1    g0467(.A(KEYINPUT29), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n641), .A2(new_n668), .A3(new_n651), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n623), .A2(new_n625), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n628), .B1(new_n536), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n620), .A2(new_n671), .A3(KEYINPUT92), .ZN(new_n672));
  INV_X1    g0472(.A(new_n626), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT92), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(KEYINPUT26), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n633), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n656), .B1(new_n552), .B2(new_n600), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(new_n572), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n651), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT29), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n669), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G330), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n520), .A2(new_n567), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n465), .A2(new_n684), .A3(new_n596), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT30), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n465), .A2(new_n684), .A3(KEYINPUT30), .A4(new_n596), .ZN(new_n688));
  AOI21_X1  g0488(.A(G179), .B1(new_n457), .B2(new_n461), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n563), .A3(new_n524), .A4(new_n590), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  AOI211_X1 g0491(.A(KEYINPUT91), .B(KEYINPUT31), .C1(new_n691), .C2(new_n650), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n605), .A2(new_n572), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(new_n651), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n650), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT91), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT31), .B1(new_n691), .B2(new_n650), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n683), .B1(new_n694), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n682), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n247), .ZN(new_n704));
  INV_X1    g0504(.A(new_n204), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n503), .A2(G116), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n226), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n704), .A2(new_n711), .ZN(G364));
  NAND2_X1  g0512(.A1(new_n644), .A2(G45), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n707), .A2(G1), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n660), .A2(new_n604), .ZN(new_n715));
  NOR3_X1   g0515(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n223), .B1(G20), .B2(new_n308), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n375), .A2(G200), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT95), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n224), .A2(G190), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n483), .ZN(new_n723));
  NAND3_X1  g0523(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n296), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n723), .B1(G50), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g0526(.A(KEYINPUT94), .B(G159), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G179), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n721), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT32), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n224), .A2(new_n296), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n720), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G87), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n726), .A2(new_n276), .A3(new_n732), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n375), .A2(G200), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n721), .A2(new_n738), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n739), .A2(new_n218), .B1(new_n740), .B2(new_n329), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT93), .Z(new_n742));
  NAND2_X1  g0542(.A1(new_n729), .A2(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G97), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n724), .A2(G190), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n747), .B2(new_n210), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT96), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n737), .A2(new_n742), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n739), .ZN(new_n751));
  INV_X1    g0551(.A(new_n730), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G322), .A2(new_n751), .B1(new_n752), .B2(G329), .ZN(new_n753));
  INV_X1    g0553(.A(G294), .ZN(new_n754));
  INV_X1    g0554(.A(new_n744), .ZN(new_n755));
  INV_X1    g0555(.A(G326), .ZN(new_n756));
  INV_X1    g0556(.A(new_n725), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n753), .B1(new_n754), .B2(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n740), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n276), .B1(new_n759), .B2(G311), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n747), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G303), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n734), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G283), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n722), .A2(new_n765), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n758), .A2(new_n762), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n718), .B1(new_n750), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n276), .A2(G355), .A3(new_n204), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n241), .A2(new_n290), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n705), .A2(new_n276), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G45), .B2(new_n226), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n769), .B1(G116), .B2(new_n204), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n718), .A2(new_n716), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n717), .A2(new_n768), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n715), .A2(new_n683), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n661), .A3(new_n714), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n778), .ZN(G396));
  AND3_X1   g0579(.A1(new_n331), .A2(new_n341), .A3(new_n651), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n331), .A2(new_n650), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n385), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(new_n782), .B2(new_n608), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n254), .ZN(new_n785));
  INV_X1    g0585(.A(new_n714), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n718), .A2(new_n254), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n329), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n734), .A2(new_n215), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n751), .A2(G143), .B1(G150), .B2(new_n746), .ZN(new_n790));
  INV_X1    g0590(.A(G137), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n790), .B1(new_n791), .B2(new_n757), .C1(new_n740), .C2(new_n728), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT34), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n722), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n792), .A2(new_n793), .B1(G68), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n752), .A2(G132), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n794), .A2(new_n796), .A3(new_n276), .A4(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n789), .B(new_n798), .C1(G58), .C2(new_n744), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n795), .A2(G87), .B1(G311), .B2(new_n752), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n276), .B1(new_n735), .B2(G107), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n800), .A2(new_n801), .A3(new_n745), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n757), .A2(new_n763), .B1(new_n740), .B2(new_n577), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G283), .B2(new_n746), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT97), .Z(new_n805));
  AOI211_X1 g0605(.A(new_n802), .B(new_n805), .C1(G294), .C2(new_n751), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n718), .B1(new_n799), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n785), .A2(new_n786), .A3(new_n788), .A4(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n784), .B1(new_n642), .B2(new_n650), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n626), .A2(new_n628), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n671), .A2(KEYINPUT90), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n629), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n665), .A2(new_n656), .A3(new_n636), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n677), .B1(new_n813), .B2(new_n572), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n651), .B(new_n783), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n809), .A2(new_n701), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT98), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n701), .B1(new_n809), .B2(new_n815), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(new_n786), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n808), .B1(new_n817), .B2(new_n819), .ZN(G384));
  INV_X1    g0620(.A(KEYINPUT101), .ZN(new_n821));
  INV_X1    g0621(.A(new_n648), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n407), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT99), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(KEYINPUT99), .B1(new_n407), .B2(new_n822), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n432), .A2(new_n427), .ZN(new_n828));
  OAI21_X1  g0628(.A(KEYINPUT37), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n828), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n823), .A2(KEYINPUT100), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT100), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n407), .A2(new_n833), .A3(new_n822), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n829), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n607), .B1(new_n612), .B2(new_n613), .ZN(new_n837));
  INV_X1    g0637(.A(new_n827), .ZN(new_n838));
  OAI211_X1 g0638(.A(KEYINPUT38), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n439), .A2(new_n827), .ZN(new_n841));
  AOI21_X1  g0641(.A(KEYINPUT38), .B1(new_n841), .B2(new_n836), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n821), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(KEYINPUT101), .A3(new_n839), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n634), .A2(new_n678), .A3(new_n604), .A4(new_n651), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n695), .B1(new_n698), .B2(KEYINPUT103), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT103), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n691), .A2(new_n850), .A3(KEYINPUT31), .A4(new_n650), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n353), .A2(new_n650), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n373), .B(new_n853), .C1(new_n380), .C2(new_n381), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n382), .A2(new_n650), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n852), .A2(new_n783), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n843), .A2(new_n847), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT40), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT102), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n832), .A2(new_n834), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT37), .B1(new_n861), .B2(new_n828), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n835), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n861), .B1(new_n607), .B2(new_n610), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n839), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n841), .A2(KEYINPUT102), .A3(KEYINPUT38), .A4(new_n836), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n859), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n858), .A2(new_n859), .B1(new_n857), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n852), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n442), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n869), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(G330), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n607), .A2(new_n648), .ZN(new_n874));
  INV_X1    g0674(.A(new_n856), .ZN(new_n875));
  INV_X1    g0675(.A(new_n780), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n815), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n843), .A2(new_n877), .A3(new_n847), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n866), .A2(new_n867), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n846), .A2(KEYINPUT39), .A3(new_n839), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n380), .A2(new_n381), .A3(new_n650), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n874), .B(new_n878), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n682), .A2(new_n442), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(new_n617), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n886), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n873), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n247), .B2(new_n644), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n577), .B1(new_n489), .B2(KEYINPUT35), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n892), .B(new_n225), .C1(KEYINPUT35), .C2(new_n489), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT36), .ZN(new_n894));
  OAI21_X1  g0694(.A(G77), .B1(new_n218), .B2(new_n210), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n895), .A2(new_n226), .B1(G50), .B2(new_n210), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(G1), .A3(new_n249), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n891), .A2(new_n894), .A3(new_n897), .ZN(G367));
  INV_X1    g0698(.A(new_n231), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n771), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n716), .B(new_n718), .C1(new_n324), .C2(new_n705), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n714), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n735), .A2(G58), .B1(G137), .B2(new_n752), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n276), .B1(new_n747), .B2(new_n728), .C1(new_n904), .C2(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(KEYINPUT104), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n795), .A2(G77), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n751), .A2(G150), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n744), .A2(G68), .B1(G143), .B2(new_n725), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n906), .A2(new_n907), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n905), .B(new_n910), .C1(G50), .C2(new_n759), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT105), .Z(new_n912));
  NOR2_X1   g0712(.A1(new_n740), .A2(new_n765), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n744), .A2(G107), .B1(G294), .B2(new_n746), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n752), .A2(G317), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(new_n334), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n722), .A2(new_n492), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n916), .B(new_n917), .C1(G311), .C2(new_n725), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n735), .A2(G116), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT46), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n918), .B(new_n920), .C1(new_n763), .C2(new_n739), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n912), .B1(new_n913), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT47), .Z(new_n923));
  INV_X1    g0723(.A(new_n718), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n902), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT106), .Z(new_n926));
  OR3_X1    g0726(.A1(new_n677), .A2(new_n511), .A3(new_n651), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n531), .B1(new_n511), .B2(new_n651), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n926), .B1(new_n716), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n706), .B(KEYINPUT41), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n658), .A2(new_n661), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n664), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n703), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n663), .A2(new_n666), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n532), .A2(new_n650), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n497), .A2(new_n536), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n619), .A2(new_n532), .A3(new_n650), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT44), .Z(new_n943));
  NAND2_X1  g0743(.A1(new_n937), .A2(new_n941), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT45), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n935), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n932), .B1(new_n947), .B2(new_n703), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(G1), .A3(new_n713), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n663), .A2(new_n939), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT42), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n536), .B1(new_n939), .B2(new_n601), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n651), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n951), .A2(new_n953), .B1(KEYINPUT43), .B2(new_n929), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n941), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n662), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n956), .B(new_n958), .Z(new_n959));
  AOI21_X1  g0759(.A(new_n931), .B1(new_n949), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(G387));
  AOI21_X1  g0761(.A(new_n707), .B1(new_n703), .B2(new_n934), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n935), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n734), .A2(new_n329), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n744), .A2(new_n324), .ZN(new_n965));
  INV_X1    g0765(.A(G159), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n965), .B1(new_n757), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n276), .B1(new_n739), .B2(new_n215), .ZN(new_n968));
  OR4_X1    g0768(.A1(new_n917), .A2(new_n964), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G150), .B2(new_n752), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n210), .B2(new_n740), .C1(new_n262), .C2(new_n747), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n734), .A2(new_n754), .B1(new_n765), .B2(new_n755), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT108), .Z(new_n973));
  AOI22_X1  g0773(.A1(new_n751), .A2(G317), .B1(G311), .B2(new_n746), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n725), .A2(G322), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(new_n763), .C2(new_n740), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT48), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n973), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT49), .Z(new_n981));
  OAI221_X1 g0781(.A(new_n334), .B1(new_n756), .B2(new_n730), .C1(new_n722), .C2(new_n577), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n971), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n718), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n236), .A2(G45), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT107), .Z(new_n986));
  NOR2_X1   g0786(.A1(new_n262), .A2(G50), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT50), .ZN(new_n988));
  AOI21_X1  g0788(.A(G45), .B1(G68), .B2(G77), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n988), .A2(new_n708), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n771), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n276), .A2(new_n204), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n991), .B1(G107), .B2(new_n204), .C1(new_n708), .C2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n774), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n714), .B1(new_n655), .B2(new_n716), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n984), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n713), .A2(G1), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n963), .B(new_n996), .C1(new_n998), .C2(new_n934), .ZN(G393));
  XOR2_X1   g0799(.A(new_n946), .B(new_n662), .Z(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n947), .B1(new_n1001), .B2(new_n935), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n706), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n774), .B1(new_n492), .B2(new_n204), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n244), .B2(new_n771), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n334), .B1(new_n747), .B2(new_n763), .C1(new_n755), .C2(new_n577), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1006), .B(new_n723), .C1(G322), .C2(new_n752), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n735), .A2(G283), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n759), .A2(G294), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n751), .A2(G311), .B1(G317), .B2(new_n725), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n751), .A2(G159), .B1(G150), .B2(new_n725), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT51), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G87), .B2(new_n795), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n735), .A2(G68), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n759), .A2(new_n321), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n276), .B1(new_n747), .B2(new_n215), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G143), .B2(new_n752), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n755), .A2(new_n329), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1013), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n714), .B(new_n1005), .C1(new_n1023), .C2(new_n718), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n957), .A2(new_n716), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT109), .Z(new_n1026));
  AOI22_X1  g0826(.A1(new_n1000), .A2(new_n997), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1003), .A2(new_n1027), .ZN(G390));
  NAND3_X1  g0828(.A1(new_n852), .A2(G330), .A3(new_n783), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1029), .A2(new_n875), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n815), .A2(new_n876), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n884), .B1(new_n1031), .B2(new_n856), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n881), .B2(new_n882), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n782), .A2(new_n608), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n651), .B(new_n1034), .C1(new_n676), .C2(new_n679), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n856), .B1(new_n1036), .B2(new_n780), .ZN(new_n1037));
  AND3_X1   g0837(.A1(new_n1037), .A2(new_n879), .A3(new_n885), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1030), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n694), .A2(new_n700), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1040), .A2(G330), .A3(new_n783), .A4(new_n856), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1037), .A2(new_n879), .A3(new_n885), .ZN(new_n1042));
  AOI21_X1  g0842(.A(KEYINPUT39), .B1(new_n866), .B2(new_n867), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n882), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1041), .B(new_n1042), .C1(new_n1045), .C2(new_n1032), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n442), .A2(new_n683), .A3(new_n870), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n887), .A2(new_n617), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1029), .A2(new_n875), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1035), .A2(new_n876), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n1041), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(KEYINPUT111), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n856), .B1(new_n701), .B2(new_n783), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1031), .B1(new_n1053), .B2(new_n1030), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT111), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1049), .A2(new_n1041), .A3(new_n1050), .A4(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1039), .A2(new_n1046), .A3(new_n1048), .A4(new_n1057), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(new_n706), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1039), .A2(new_n1046), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1048), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n997), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n883), .A2(new_n254), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n787), .A2(new_n262), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1022), .B1(G97), .B2(new_n759), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n334), .C1(new_n577), .C2(new_n739), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n735), .A2(G87), .B1(new_n746), .B2(G107), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n210), .B2(new_n722), .C1(new_n754), .C2(new_n730), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1068), .B(new_n1070), .C1(G283), .C2(new_n725), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n795), .A2(G50), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n734), .A2(new_n267), .ZN(new_n1073));
  XOR2_X1   g0873(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n1074));
  XNOR2_X1  g0874(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n334), .B1(new_n752), .B2(G125), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n755), .A2(new_n966), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT54), .B(G143), .Z(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1079), .A2(new_n740), .B1(new_n791), .B2(new_n747), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1077), .B(new_n1080), .C1(G128), .C2(new_n725), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1075), .A2(new_n1076), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G132), .B2(new_n751), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1071), .B1(new_n1072), .B2(new_n1083), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT113), .Z(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n718), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1065), .A2(new_n786), .A3(new_n1066), .A4(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1063), .A2(new_n1064), .A3(new_n1087), .ZN(G378));
  INV_X1    g0888(.A(KEYINPUT57), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1058), .A2(new_n1048), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n886), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n858), .A2(new_n859), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n868), .A2(new_n857), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT119), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n273), .A2(new_n822), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n306), .A2(new_n310), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n306), .B2(new_n310), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1100), .A2(new_n1096), .A3(new_n1101), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1095), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1104), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(KEYINPUT119), .A3(new_n1102), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  AND4_X1   g0908(.A1(G330), .A2(new_n1093), .A3(new_n1094), .A4(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n869), .B2(G330), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1092), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1093), .A2(G330), .A3(new_n1094), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1110), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n869), .A2(G330), .A3(new_n1108), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n886), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1089), .B1(new_n1091), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1090), .A2(KEYINPUT57), .A3(new_n1112), .A4(new_n1117), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n706), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1112), .A2(new_n997), .A3(new_n1117), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1105), .A2(new_n1107), .A3(new_n254), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n964), .B1(G97), .B2(new_n746), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n759), .A2(new_n324), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(new_n218), .C2(new_n722), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n744), .A2(G68), .B1(G116), .B2(new_n725), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1127), .B(new_n289), .C1(new_n765), .C2(new_n730), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n739), .A2(new_n483), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT114), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1126), .A2(new_n276), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT115), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n1133));
  XNOR2_X1  g0933(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n735), .A2(new_n1078), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n751), .A2(G128), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n759), .A2(G137), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G125), .A2(new_n725), .B1(new_n746), .B2(G132), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G150), .B2(new_n744), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT117), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT59), .ZN(new_n1142));
  INV_X1    g0942(.A(G124), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n730), .B1(KEYINPUT118), .B2(new_n1143), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1143), .A2(KEYINPUT118), .ZN(new_n1145));
  AOI211_X1 g0945(.A(G33), .B(G41), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1142), .B(new_n1146), .C1(new_n722), .C2(new_n728), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n215), .B1(new_n332), .B2(G41), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1134), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n718), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n787), .A2(new_n215), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1123), .A2(new_n786), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT120), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1122), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT121), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1122), .A2(new_n1155), .A3(KEYINPUT121), .A4(new_n1154), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1121), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT122), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1121), .A2(KEYINPUT122), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(G375));
  OR2_X1    g0964(.A1(new_n1057), .A2(new_n1048), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n932), .A3(new_n1061), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n795), .A2(G58), .B1(G150), .B2(new_n759), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1167), .B1(new_n966), .B2(new_n734), .C1(new_n747), .C2(new_n1079), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G137), .B2(new_n751), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n744), .A2(G50), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n334), .B1(new_n725), .B2(G132), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G128), .B2(new_n752), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n907), .B1(new_n765), .B2(new_n739), .C1(new_n763), .C2(new_n730), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n276), .B1(new_n725), .B2(G294), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n965), .C1(new_n483), .C2(new_n740), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n747), .A2(new_n577), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n734), .A2(new_n492), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n718), .B1(new_n1173), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n254), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n786), .B(new_n1180), .C1(new_n856), .C2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n210), .B2(new_n787), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1057), .B2(new_n997), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1166), .A2(new_n1184), .ZN(G381));
  NOR2_X1   g0985(.A1(G375), .A2(G378), .ZN(new_n1186));
  INV_X1    g0986(.A(G390), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(G393), .A2(G396), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(G387), .A2(G384), .A3(G381), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(G407));
  NAND2_X1  g0990(.A1(new_n1186), .A2(new_n649), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(G407), .A2(G213), .A3(new_n1191), .ZN(G409));
  XOR2_X1   g0992(.A(G393), .B(G396), .Z(new_n1193));
  NAND2_X1  g0993(.A1(new_n960), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT126), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n960), .A2(new_n1196), .A3(new_n1193), .ZN(new_n1197));
  OR3_X1    g0997(.A1(new_n1195), .A2(new_n1197), .A3(new_n1187), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1187), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT60), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n707), .B1(new_n1165), .B2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1202), .B(new_n1061), .C1(new_n1201), .C2(new_n1165), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1203), .A2(G384), .A3(new_n1184), .ZN(new_n1204));
  AOI21_X1  g1004(.A(G384), .B1(new_n1203), .B2(new_n1184), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n649), .A2(G213), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1122), .A2(new_n1152), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT124), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT123), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1210), .A2(new_n1211), .A3(new_n932), .A4(new_n1090), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1090), .A2(new_n932), .A3(new_n1112), .A4(new_n1117), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT123), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT124), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1122), .A2(new_n1215), .A3(new_n1152), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1209), .A2(new_n1212), .A3(new_n1214), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT125), .ZN(new_n1218));
  INV_X1    g1018(.A(G378), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1121), .A2(G378), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1218), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1206), .B(new_n1207), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1200), .B1(new_n1225), .B2(KEYINPUT63), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n649), .A2(G213), .A3(G2897), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1206), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1227), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT125), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1231), .B1(new_n1234), .B2(new_n1207), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT63), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1224), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT61), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1226), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1224), .A2(KEYINPUT62), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1207), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1231), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1238), .B1(new_n1224), .B2(KEYINPUT62), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1200), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1239), .A2(new_n1246), .ZN(G405));
  AND2_X1   g1047(.A1(new_n1221), .A2(KEYINPUT127), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G375), .B2(new_n1219), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT127), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1250), .B(G378), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1206), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(G375), .A2(KEYINPUT127), .A3(new_n1219), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1206), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G378), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1253), .B(new_n1254), .C1(new_n1255), .C2(new_n1248), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1200), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1252), .A2(new_n1256), .A3(new_n1199), .A4(new_n1198), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(G402));
endmodule


