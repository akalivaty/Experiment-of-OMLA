//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(KEYINPUT65), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n210), .B1(new_n211), .B2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G13), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n213), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(G50), .B2(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n203), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n233));
  INV_X1    g0033(.A(KEYINPUT66), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G20), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(G1), .A2(G13), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G50), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n206), .A2(new_n239), .ZN(new_n240));
  AOI211_X1 g0040(.A(new_n217), .B(new_n231), .C1(new_n238), .C2(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G250), .B(G257), .Z(new_n246));
  XNOR2_X1  g0046(.A(G264), .B(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G68), .B(G77), .Z(new_n253));
  XNOR2_X1  g0053(.A(G50), .B(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT70), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G223), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G222), .ZN(new_n264));
  OR3_X1    g0064(.A1(new_n263), .A2(KEYINPUT69), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT69), .B1(new_n263), .B2(new_n264), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G77), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n261), .A2(new_n265), .A3(new_n266), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT71), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n274), .A2(KEYINPUT71), .A3(G1), .A4(G13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(G41), .B2(G45), .ZN(new_n282));
  OR2_X1    g0082(.A1(KEYINPUT68), .A2(G226), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT68), .A2(G226), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n275), .A2(new_n282), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT67), .B(G41), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n281), .B(G274), .C1(new_n286), .C2(G45), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n280), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(G20), .B1(new_n207), .B2(G50), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G150), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n236), .A2(G33), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n291), .B(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n237), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n281), .A2(G13), .A3(G20), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n296), .A2(new_n298), .B1(new_n239), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n297), .A2(new_n237), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n281), .A2(G20), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G50), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n290), .B(new_n307), .C1(G179), .C2(new_n288), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n288), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n307), .B(KEYINPUT9), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n288), .A2(G200), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT10), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n311), .A2(new_n316), .A3(new_n312), .A4(new_n313), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n309), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n303), .ZN(new_n319));
  OR3_X1    g0119(.A1(new_n295), .A2(new_n319), .A3(KEYINPUT77), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT77), .B1(new_n295), .B2(new_n319), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n320), .A2(new_n302), .A3(new_n299), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n295), .A2(new_n300), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT76), .B1(new_n269), .B2(G33), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT76), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(new_n267), .A3(KEYINPUT3), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n327), .A3(new_n270), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT7), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n233), .B2(new_n235), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n329), .B1(new_n257), .B2(G20), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n203), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n335), .A2(G20), .B1(G159), .B2(new_n292), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT16), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT7), .B1(new_n257), .B2(G20), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n236), .A2(new_n271), .A3(new_n329), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n339), .A3(G68), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(new_n336), .A3(KEYINPUT16), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n298), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n324), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n268), .A2(new_n270), .A3(G226), .A4(G1698), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT78), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT78), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n257), .A2(new_n346), .A3(G226), .A4(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G87), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n257), .A2(G223), .A3(new_n262), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n345), .A2(new_n347), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n279), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n275), .A2(new_n282), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n287), .B1(new_n224), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(G179), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n353), .B1(new_n350), .B2(new_n279), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n355), .B1(new_n289), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n343), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT18), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT16), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n335), .A2(G20), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n292), .A2(G159), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n360), .B1(new_n333), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(new_n298), .A3(new_n341), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n351), .A2(new_n310), .A3(new_n354), .ZN(new_n366));
  AOI21_X1  g0166(.A(G200), .B1(new_n351), .B2(new_n354), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n365), .B(new_n324), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT17), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n368), .B(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n359), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n295), .B(KEYINPUT72), .ZN(new_n372));
  INV_X1    g0172(.A(new_n292), .ZN(new_n373));
  XOR2_X1   g0173(.A(KEYINPUT15), .B(G87), .Z(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n372), .A2(new_n373), .B1(new_n294), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G77), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n236), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n298), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n304), .A2(new_n377), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n299), .A2(G77), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n379), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n271), .A2(G107), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n257), .A2(G232), .A3(new_n262), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n258), .B(KEYINPUT70), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n385), .B(new_n386), .C1(new_n387), .C2(new_n228), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n279), .ZN(new_n389));
  INV_X1    g0189(.A(G244), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n352), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(new_n287), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n384), .B1(new_n393), .B2(G200), .ZN(new_n394));
  INV_X1    g0194(.A(new_n287), .ZN(new_n395));
  AOI211_X1 g0195(.A(new_n395), .B(new_n391), .C1(new_n388), .C2(new_n279), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G190), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n318), .A2(new_n371), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n292), .A2(G50), .ZN(new_n400));
  OAI221_X1 g0200(.A(new_n400), .B1(new_n232), .B2(G68), .C1(new_n294), .C2(new_n377), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n298), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT11), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n305), .A2(G68), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n299), .A2(G68), .ZN(new_n405));
  XNOR2_X1  g0205(.A(KEYINPUT74), .B(KEYINPUT12), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT12), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n407), .A2(KEYINPUT75), .B1(new_n408), .B2(new_n405), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(KEYINPUT75), .B2(new_n407), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n403), .A2(new_n404), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n352), .A2(new_n228), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n257), .A2(G226), .A3(new_n262), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G97), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n268), .A2(new_n270), .A3(G232), .A4(G1698), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n412), .B1(new_n416), .B2(new_n279), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT13), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n417), .A2(new_n418), .A3(new_n287), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n418), .B1(new_n417), .B2(new_n287), .ZN(new_n420));
  OAI21_X1  g0220(.A(G169), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT14), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT14), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(G169), .C1(new_n419), .C2(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G179), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n417), .A2(new_n287), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT13), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n417), .A2(new_n418), .A3(new_n287), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(KEYINPUT73), .A3(new_n429), .ZN(new_n430));
  OR3_X1    g0230(.A1(new_n427), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n411), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n431), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G190), .ZN(new_n435));
  INV_X1    g0235(.A(new_n411), .ZN(new_n436));
  OAI21_X1  g0236(.A(G200), .B1(new_n419), .B2(new_n420), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n389), .A2(new_n426), .A3(new_n287), .A4(new_n392), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(new_n384), .C1(new_n396), .C2(G169), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n433), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n399), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT85), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT24), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT66), .B(G20), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT23), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n225), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT23), .B1(new_n232), .B2(G107), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n236), .A2(new_n257), .A3(G87), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT22), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT22), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n236), .A2(new_n257), .A3(new_n452), .A4(G87), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n449), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n443), .A2(KEYINPUT24), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n232), .A2(G33), .A3(G116), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n456), .B1(new_n454), .B2(new_n457), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n444), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n281), .A2(G33), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n302), .A2(new_n299), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n461), .A2(new_n298), .B1(G107), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n299), .A2(G107), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n466), .B(KEYINPUT25), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n281), .B(G45), .C1(new_n468), .C2(G41), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n286), .B2(new_n468), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G274), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n257), .A2(G257), .A3(G1698), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n257), .A2(G250), .A3(new_n262), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G294), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n279), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT86), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n237), .B1(G33), .B2(G41), .ZN(new_n478));
  NOR4_X1   g0278(.A1(new_n470), .A2(new_n477), .A3(new_n226), .A4(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n469), .ZN(new_n480));
  INV_X1    g0280(.A(G41), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT67), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT67), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G41), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n484), .A3(new_n468), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n478), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT86), .B1(new_n486), .B2(G264), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n471), .B(new_n476), .C1(new_n479), .C2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(new_n310), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(G200), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n465), .A2(new_n467), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n464), .A2(G107), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n451), .A2(new_n453), .ZN(new_n494));
  INV_X1    g0294(.A(new_n449), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n457), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n455), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(new_n458), .B1(new_n443), .B2(KEYINPUT24), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n493), .B(new_n467), .C1(new_n498), .C2(new_n302), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n488), .A2(G169), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n482), .A2(new_n484), .A3(new_n468), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n275), .B1(new_n501), .B2(new_n469), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n477), .B1(new_n502), .B2(new_n226), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n486), .A2(KEYINPUT86), .A3(G264), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(G179), .A3(new_n471), .A4(new_n476), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT87), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n500), .A2(new_n506), .A3(KEYINPUT87), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n499), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n464), .A2(G116), .ZN(new_n511));
  INV_X1    g0311(.A(G116), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n300), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n302), .B1(G20), .B2(new_n512), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  INV_X1    g0315(.A(G97), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n236), .B(new_n515), .C1(G33), .C2(new_n516), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n514), .A2(KEYINPUT20), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT20), .B1(new_n514), .B2(new_n517), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n511), .B(new_n513), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n257), .A2(G257), .A3(new_n262), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n271), .A2(G303), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n258), .C2(new_n226), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n279), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n486), .A2(G270), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n471), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(G169), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n520), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n526), .A2(G200), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(new_n531), .C1(new_n310), .C2(new_n526), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n526), .A2(new_n426), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n520), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n520), .A2(KEYINPUT21), .A3(G169), .A4(new_n526), .ZN(new_n535));
  AND4_X1   g0335(.A1(new_n529), .A2(new_n532), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n492), .A2(new_n510), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(G257), .B(new_n275), .C1(new_n501), .C2(new_n469), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT82), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n486), .A2(KEYINPUT82), .A3(G257), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n540), .A2(new_n471), .A3(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n268), .A2(new_n270), .A3(G244), .A4(new_n262), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n515), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n279), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT81), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(KEYINPUT81), .A3(new_n279), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n542), .A2(new_n426), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n549), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n540), .A2(new_n471), .A3(new_n541), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n289), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n463), .A2(G97), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n299), .A2(new_n516), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT80), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n557), .A2(KEYINPUT80), .A3(new_n558), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n564));
  AND2_X1   g0364(.A1(G97), .A2(G107), .ZN(new_n565));
  NOR2_X1   g0365(.A1(G97), .A2(G107), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g0367(.A(G97), .B(G107), .ZN(new_n568));
  NAND2_X1  g0368(.A1(KEYINPUT6), .A2(G107), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(KEYINPUT79), .B2(KEYINPUT6), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n567), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n445), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n292), .A2(G77), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n225), .B1(new_n331), .B2(new_n332), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n298), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n563), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n553), .A2(new_n556), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT83), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT83), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n553), .A2(new_n580), .A3(new_n556), .A4(new_n577), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n281), .A2(G45), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n275), .A2(G250), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n228), .A2(new_n262), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n390), .A2(G1698), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n268), .A2(new_n586), .A3(new_n270), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G116), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n585), .B1(new_n590), .B2(new_n279), .ZN(new_n591));
  INV_X1    g0391(.A(G274), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n583), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(G169), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n374), .A2(new_n299), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n236), .A2(G33), .A3(G97), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT19), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n236), .A2(new_n257), .A3(G68), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n566), .A2(KEYINPUT84), .A3(new_n220), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT84), .B1(new_n566), .B2(new_n220), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n414), .A2(new_n598), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n601), .A2(new_n602), .B1(new_n445), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n599), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n596), .B1(new_n605), .B2(new_n298), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n464), .A2(new_n374), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n595), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n591), .A2(new_n594), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n426), .ZN(new_n611));
  INV_X1    g0411(.A(G200), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n591), .B2(new_n594), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n588), .A2(new_n589), .B1(new_n277), .B2(new_n278), .ZN(new_n614));
  NOR4_X1   g0414(.A1(new_n614), .A2(new_n310), .A3(new_n593), .A4(new_n585), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n463), .A2(new_n220), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n596), .B(new_n617), .C1(new_n605), .C2(new_n298), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n608), .A2(new_n611), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n542), .A2(new_n551), .A3(new_n552), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n554), .A2(new_n555), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n620), .A2(G200), .B1(new_n621), .B2(G190), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n331), .A2(new_n332), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G107), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n572), .A3(new_n573), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n625), .A2(new_n298), .B1(new_n561), .B2(new_n562), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n582), .A2(new_n619), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n537), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n442), .A2(new_n629), .ZN(G372));
  INV_X1    g0430(.A(new_n552), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT81), .B1(new_n548), .B2(new_n279), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n631), .A2(new_n555), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n626), .B1(new_n633), .B2(new_n426), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n634), .A2(new_n619), .A3(new_n635), .A4(new_n556), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n608), .A2(new_n611), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n579), .A2(new_n619), .A3(new_n581), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(KEYINPUT26), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n500), .A2(new_n506), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n499), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n529), .A2(new_n534), .A3(new_n535), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n579), .A2(new_n581), .B1(new_n626), .B2(new_n622), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(new_n619), .A4(new_n492), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n442), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT18), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n358), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n434), .A2(G179), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n422), .A3(new_n424), .ZN(new_n653));
  INV_X1    g0453(.A(new_n440), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n411), .A2(new_n653), .B1(new_n438), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n651), .B1(new_n655), .B2(new_n370), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n315), .A2(new_n317), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n309), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n649), .A2(new_n658), .ZN(G369));
  NOR2_X1   g0459(.A1(new_n445), .A2(new_n213), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n281), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n530), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT88), .B1(new_n644), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n536), .A2(new_n669), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT88), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n643), .A2(new_n672), .A3(new_n668), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n499), .A2(new_n666), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n492), .A2(new_n510), .A3(new_n677), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n500), .A2(new_n506), .A3(KEYINPUT87), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n507), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n499), .A3(new_n666), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n666), .B(KEYINPUT89), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n499), .A2(new_n684), .A3(new_n641), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n534), .A2(new_n535), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n666), .B1(new_n687), .B2(new_n529), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(new_n492), .A3(new_n510), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n683), .A2(new_n685), .A3(new_n689), .ZN(G399));
  NOR3_X1   g0490(.A1(new_n601), .A2(new_n602), .A3(G116), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT90), .Z(new_n692));
  INV_X1    g0492(.A(new_n215), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n286), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n692), .A2(new_n281), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n240), .B2(new_n694), .ZN(new_n696));
  XNOR2_X1  g0496(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n684), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n640), .B2(new_n647), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n510), .A2(new_n644), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n703), .A2(new_n619), .A3(new_n646), .A4(new_n492), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n579), .A2(new_n635), .A3(new_n619), .A4(new_n581), .ZN(new_n705));
  INV_X1    g0505(.A(new_n619), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT26), .B1(new_n706), .B2(new_n578), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n705), .A2(new_n707), .A3(new_n637), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n666), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n702), .B1(new_n701), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n526), .A2(new_n426), .A3(new_n609), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n503), .A2(new_n504), .B1(new_n279), .B2(new_n475), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n621), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT93), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n713), .A2(KEYINPUT30), .A3(new_n621), .A4(new_n714), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n620), .A2(new_n426), .A3(new_n488), .A4(new_n526), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n718), .B(new_n719), .C1(new_n610), .C2(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n715), .A2(new_n717), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n716), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n666), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n629), .A2(new_n684), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n719), .B1(new_n720), .B2(new_n610), .ZN(new_n727));
  OAI211_X1 g0527(.A(KEYINPUT31), .B(new_n699), .C1(new_n727), .C2(new_n722), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT92), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n712), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n711), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n698), .B1(new_n732), .B2(G1), .ZN(G364));
  AOI21_X1  g0533(.A(new_n281), .B1(new_n660), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n694), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n676), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G330), .B2(new_n674), .ZN(new_n738));
  INV_X1    g0538(.A(new_n736), .ZN(new_n739));
  INV_X1    g0539(.A(G45), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n240), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n693), .A2(new_n257), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n741), .B(new_n742), .C1(new_n255), .C2(new_n740), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n215), .A2(G355), .A3(new_n257), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n743), .B(new_n744), .C1(G116), .C2(new_n215), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n237), .B1(G20), .B2(new_n289), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n739), .B1(new_n745), .B2(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT94), .Z(new_n752));
  NOR2_X1   g0552(.A1(new_n236), .A2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n612), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G283), .ZN(new_n756));
  INV_X1    g0556(.A(G329), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n271), .B1(new_n755), .B2(new_n756), .C1(new_n757), .C2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n236), .B1(G190), .B2(new_n758), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT97), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(KEYINPUT97), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G294), .ZN(new_n766));
  INV_X1    g0566(.A(G326), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n426), .A2(new_n310), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n445), .A2(G200), .A3(new_n768), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(KEYINPUT98), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n753), .A2(G179), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n612), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n760), .B(new_n771), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n754), .A2(G20), .A3(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G303), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n772), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G311), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n445), .A2(new_n612), .A3(new_n768), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n770), .A2(KEYINPUT98), .B1(G322), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n779), .A2(new_n782), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n759), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G159), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(KEYINPUT32), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n777), .A2(G68), .B1(KEYINPUT32), .B2(new_n790), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n781), .A2(G87), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n257), .B(new_n793), .C1(new_n755), .C2(new_n225), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT95), .Z(new_n795));
  INV_X1    g0595(.A(new_n769), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G50), .A2(new_n796), .B1(new_n786), .B2(G58), .ZN(new_n797));
  INV_X1    g0597(.A(new_n783), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n798), .B2(new_n377), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G97), .B2(new_n764), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n792), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n788), .B1(new_n791), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n752), .B1(new_n802), .B2(new_n749), .ZN(new_n803));
  INV_X1    g0603(.A(new_n748), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n674), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n738), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  AOI22_X1  g0607(.A1(new_n783), .A2(G159), .B1(G143), .B2(new_n786), .ZN(new_n808));
  INV_X1    g0608(.A(G137), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n809), .B2(new_n769), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n777), .B2(G150), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT34), .Z(new_n812));
  INV_X1    g0612(.A(new_n755), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G68), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n789), .A2(G132), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n271), .B1(new_n781), .B2(G50), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n812), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G58), .B2(new_n764), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n755), .A2(new_n220), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n777), .B2(G283), .ZN(new_n820));
  INV_X1    g0620(.A(G303), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n512), .B2(new_n798), .C1(new_n821), .C2(new_n769), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n780), .A2(new_n225), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n271), .B1(new_n765), .B2(new_n516), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n759), .A2(new_n825), .B1(new_n766), .B2(new_n785), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n749), .B1(new_n818), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n749), .A2(new_n746), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT99), .Z(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n377), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n393), .A2(new_n289), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n832), .A2(new_n384), .A3(new_n439), .A4(new_n667), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n384), .A2(new_n666), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n394), .B2(new_n397), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n833), .B1(new_n835), .B2(new_n654), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n739), .B1(new_n836), .B2(new_n746), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n828), .A2(new_n831), .A3(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT100), .Z(new_n839));
  INV_X1    g0639(.A(new_n730), .ZN(new_n840));
  INV_X1    g0640(.A(new_n836), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n700), .A2(new_n841), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n699), .B(new_n836), .C1(new_n640), .C2(new_n647), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n840), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n739), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n839), .A2(new_n846), .ZN(G384));
  AND3_X1   g0647(.A1(new_n492), .A2(new_n510), .A3(new_n536), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n848), .A2(new_n619), .A3(new_n646), .A4(new_n684), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n724), .A2(new_n725), .ZN(new_n850));
  OAI211_X1 g0650(.A(KEYINPUT31), .B(new_n666), .C1(new_n721), .C2(new_n723), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n411), .A2(new_n666), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n433), .A2(new_n438), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT101), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n433), .A2(new_n438), .A3(KEYINPUT101), .A4(new_n853), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n653), .A2(new_n411), .A3(new_n666), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n852), .A2(new_n860), .A3(new_n841), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT16), .B1(new_n340), .B2(new_n336), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n324), .B1(new_n342), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n357), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n664), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n368), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT102), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n343), .B1(new_n357), .B2(new_n865), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(new_n368), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT102), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n867), .A2(new_n873), .A3(KEYINPUT37), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n869), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n866), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n359), .B2(new_n370), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(KEYINPUT38), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n343), .A2(new_n865), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n368), .B(KEYINPUT17), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(new_n651), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n872), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n871), .B1(new_n870), .B2(new_n368), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n879), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT40), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n861), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT40), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n867), .A2(new_n873), .A3(KEYINPUT37), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n873), .B1(new_n867), .B2(KEYINPUT37), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n891), .A2(new_n892), .A3(new_n883), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n866), .B1(new_n651), .B2(new_n881), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n879), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n878), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n890), .B1(new_n861), .B2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n889), .A2(new_n898), .A3(new_n442), .A4(new_n852), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n889), .A2(G330), .A3(new_n898), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n442), .A2(G330), .A3(new_n852), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n711), .A2(new_n442), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n658), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n903), .B(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n887), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n653), .A2(new_n411), .A3(new_n667), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n878), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n833), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n896), .B(new_n860), .C1(new_n843), .C2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n651), .A2(new_n865), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n912), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT103), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT103), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n912), .A2(new_n914), .A3(new_n919), .A4(new_n916), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n906), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n281), .B2(new_n660), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n512), .B1(new_n571), .B2(KEYINPUT35), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n924), .B(new_n238), .C1(KEYINPUT35), .C2(new_n571), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT36), .ZN(new_n926));
  INV_X1    g0726(.A(new_n240), .ZN(new_n927));
  OAI21_X1  g0727(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n927), .A2(new_n928), .B1(G50), .B2(new_n203), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(G1), .A3(new_n213), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n923), .A2(new_n926), .A3(new_n930), .ZN(G367));
  INV_X1    g0731(.A(G317), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n271), .B1(new_n755), .B2(new_n516), .C1(new_n932), .C2(new_n759), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n933), .A2(KEYINPUT110), .B1(new_n756), .B2(new_n798), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n776), .A2(new_n766), .B1(new_n225), .B2(new_n765), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n934), .B(new_n935), .C1(G303), .C2(new_n786), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n781), .A2(KEYINPUT46), .A3(G116), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n796), .A2(G311), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT46), .B1(new_n781), .B2(G116), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n933), .B2(KEYINPUT110), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n936), .A2(new_n937), .A3(new_n938), .A4(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n765), .A2(new_n203), .ZN(new_n942));
  INV_X1    g0742(.A(G159), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n257), .B1(new_n809), .B2(new_n759), .C1(new_n776), .C2(new_n943), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n942), .B(new_n944), .C1(G143), .C2(new_n796), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n786), .A2(G150), .B1(G58), .B2(new_n781), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n945), .B(new_n946), .C1(new_n239), .C2(new_n798), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n755), .A2(new_n377), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n941), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT47), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n950), .A2(new_n749), .ZN(new_n951));
  INV_X1    g0751(.A(new_n742), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n750), .B1(new_n215), .B2(new_n375), .C1(new_n952), .C2(new_n248), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n637), .A2(new_n618), .A3(new_n667), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n619), .B1(new_n618), .B2(new_n667), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n736), .B(new_n953), .C1(new_n956), .C2(new_n804), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n951), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n683), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n684), .A2(new_n578), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n699), .A2(new_n577), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(new_n646), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n964), .A2(KEYINPUT45), .A3(new_n685), .A4(new_n689), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n689), .A2(new_n685), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n966), .B1(new_n967), .B2(new_n963), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n963), .ZN(new_n970));
  XNOR2_X1  g0770(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT107), .Z(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n967), .A2(new_n963), .A3(new_n972), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n960), .B1(new_n969), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n965), .A2(new_n968), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n978), .A2(new_n683), .A3(new_n975), .A4(new_n974), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n678), .B(new_n681), .C1(new_n644), .C2(new_n666), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n689), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n676), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n675), .A2(new_n981), .A3(new_n689), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n710), .A2(new_n701), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n840), .A2(new_n985), .A3(new_n986), .A4(new_n702), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT108), .B1(new_n980), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n984), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n675), .B1(new_n689), .B2(new_n981), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n991), .A2(new_n711), .A3(new_n730), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT108), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n992), .A2(new_n993), .A3(new_n977), .A4(new_n979), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n731), .B1(new_n988), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n694), .B(KEYINPUT41), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n734), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n582), .B1(new_n963), .B2(new_n510), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n684), .ZN(new_n1000));
  OAI21_X1  g0800(.A(KEYINPUT42), .B1(new_n963), .B2(new_n689), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT104), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1000), .A2(KEYINPUT104), .A3(new_n1001), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT43), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n956), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n963), .A2(new_n689), .A3(KEYINPUT42), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT105), .Z(new_n1010));
  NAND4_X1  g0810(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1008), .A2(new_n1007), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n683), .A2(new_n963), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n1011), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1016), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n998), .A2(new_n1019), .A3(KEYINPUT109), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT109), .B1(new_n998), .B2(new_n1019), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n959), .B1(new_n1020), .B2(new_n1021), .ZN(G387));
  NOR2_X1   g0822(.A1(new_n776), .A2(new_n295), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G77), .B2(new_n781), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n239), .B2(new_n785), .C1(new_n203), .C2(new_n798), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G159), .B2(new_n796), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n789), .A2(G150), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n765), .A2(new_n375), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G97), .B2(new_n813), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n257), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n796), .A2(G322), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n932), .B2(new_n785), .C1(new_n798), .C2(new_n821), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n777), .B2(G311), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT48), .Z(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n756), .B2(new_n765), .C1(new_n766), .C2(new_n780), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT49), .Z(new_n1036));
  OAI221_X1 g0836(.A(new_n271), .B1(new_n755), .B2(new_n512), .C1(new_n767), .C2(new_n759), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1030), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n749), .ZN(new_n1039));
  AOI211_X1 g0839(.A(G45), .B(new_n692), .C1(G68), .C2(G77), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n372), .A2(G50), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT50), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n692), .A2(new_n215), .A3(new_n257), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n742), .B1(new_n245), .B2(new_n740), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1040), .A2(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n215), .A2(G107), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n750), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n678), .A2(new_n681), .A3(new_n748), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1039), .A2(new_n736), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n731), .A2(new_n991), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(new_n694), .A3(new_n987), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n985), .A2(new_n735), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT111), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1049), .A2(new_n1051), .A3(new_n1053), .ZN(G393));
  AOI22_X1  g0854(.A1(new_n988), .A2(new_n994), .B1(new_n980), .B2(new_n987), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1055), .A2(new_n694), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n963), .A2(new_n748), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n750), .B1(new_n516), .B2(new_n215), .C1(new_n952), .C2(new_n252), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n777), .A2(G303), .B1(G322), .B2(new_n789), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n764), .A2(G116), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n825), .A2(new_n785), .B1(new_n769), .B2(new_n932), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT52), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n755), .A2(new_n225), .B1(new_n756), .B2(new_n780), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n257), .B(new_n1063), .C1(G294), .C2(new_n783), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n798), .A2(new_n372), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n777), .B2(G50), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n764), .A2(G77), .ZN(new_n1068));
  INV_X1    g0868(.A(G150), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1069), .A2(new_n769), .B1(new_n785), .B2(new_n943), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT51), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n780), .A2(new_n203), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1072), .B(new_n819), .C1(G143), .C2(new_n789), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1067), .A2(new_n1068), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1065), .B1(new_n1074), .B2(new_n271), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n749), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1057), .A2(new_n736), .A3(new_n1058), .A4(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n980), .B(KEYINPUT112), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n734), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1056), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(G390));
  AOI21_X1  g0881(.A(new_n913), .B1(new_n700), .B2(new_n841), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n860), .B1(new_n730), .B2(new_n841), .ZN(new_n1084));
  AND4_X1   g0884(.A1(G330), .A2(new_n852), .A3(new_n860), .A4(new_n841), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n726), .A2(new_n729), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1087), .A2(G330), .A3(new_n841), .A4(new_n860), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n835), .A2(new_n654), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n913), .B1(new_n710), .B2(new_n1089), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n852), .A2(G330), .A3(new_n841), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1088), .B(new_n1090), .C1(new_n1091), .C2(new_n860), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n901), .A2(new_n904), .A3(new_n658), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT113), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n859), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n856), .B2(new_n857), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n643), .B1(new_n680), .B2(new_n499), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n491), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n499), .A2(new_n489), .A3(new_n1101), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n628), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n667), .B(new_n1089), .C1(new_n1103), .C2(new_n708), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1099), .B1(new_n1104), .B2(new_n833), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n910), .B1(new_n878), .B2(new_n886), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1097), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(KEYINPUT113), .B(new_n1106), .C1(new_n1090), .C2(new_n1099), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n909), .B1(new_n1082), .B2(new_n1099), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n908), .A2(new_n911), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1088), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1096), .B(new_n1115), .C1(new_n1116), .C2(new_n1085), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1094), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1118));
  AOI221_X4 g0918(.A(new_n1088), .B1(new_n1111), .B2(new_n1112), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1085), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n694), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n747), .B1(new_n908), .B2(new_n911), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n830), .A2(new_n295), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n736), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT114), .Z(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT54), .B(G143), .Z(new_n1127));
  NAND2_X1  g0927(.A1(new_n783), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n776), .B2(new_n809), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n271), .B1(new_n1129), .B2(KEYINPUT115), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n789), .A2(G125), .ZN(new_n1131));
  INV_X1    g0931(.A(G132), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1130), .B(new_n1131), .C1(new_n1132), .C2(new_n785), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n781), .A2(G150), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1129), .A2(KEYINPUT115), .ZN(new_n1136));
  INV_X1    g0936(.A(G128), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n769), .A2(new_n1137), .ZN(new_n1138));
  NOR4_X1   g0938(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n239), .B2(new_n755), .C1(new_n943), .C2(new_n765), .ZN(new_n1140));
  OR2_X1    g0940(.A1(new_n1140), .A2(KEYINPUT116), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(KEYINPUT116), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n777), .A2(G107), .B1(G283), .B2(new_n796), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1143), .B(new_n814), .C1(new_n516), .C2(new_n798), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G294), .B2(new_n789), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1068), .B1(new_n512), .B2(new_n785), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT117), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1145), .A2(new_n271), .A3(new_n793), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1141), .A2(new_n1142), .A3(new_n1148), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1123), .B(new_n1126), .C1(new_n1149), .C2(new_n749), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1115), .B1(new_n1116), .B2(new_n1085), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n735), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1122), .A2(new_n1152), .ZN(G378));
  NAND2_X1  g0953(.A1(new_n1121), .A2(new_n1095), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n307), .A2(new_n865), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n318), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n318), .A2(new_n1155), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OR3_X1    g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n921), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n918), .A2(new_n1162), .A3(new_n920), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n900), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n900), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n918), .A2(new_n920), .A3(new_n1162), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1162), .B1(new_n918), .B2(new_n920), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1154), .A2(KEYINPUT57), .A3(new_n1166), .A4(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(new_n694), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1154), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1168), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n900), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1170), .A2(new_n1166), .A3(KEYINPUT120), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1173), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1172), .B1(new_n1179), .B2(KEYINPUT57), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1163), .A2(new_n746), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n829), .A2(new_n239), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n777), .A2(G132), .B1(G125), .B2(new_n796), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n765), .A2(new_n1069), .B1(new_n809), .B2(new_n798), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G128), .B2(new_n786), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n781), .A2(new_n1127), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT119), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1183), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT59), .Z(new_n1189));
  AOI211_X1 g0989(.A(G33), .B(G41), .C1(new_n789), .C2(G124), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n943), .C2(new_n755), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n786), .A2(G107), .B1(G77), .B2(new_n781), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n798), .B2(new_n375), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1193), .B(new_n942), .C1(G283), .C2(new_n789), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n755), .A2(new_n202), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT118), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G116), .B2(new_n796), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n257), .A2(new_n286), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n516), .C2(new_n776), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT58), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n239), .B1(G33), .B2(G41), .C1(new_n257), .C2(new_n286), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1191), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n749), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1181), .A2(new_n736), .A3(new_n1182), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n1209), .B2(new_n735), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1180), .A2(new_n1210), .ZN(G375));
  NAND3_X1  g1011(.A1(new_n1086), .A2(new_n1094), .A3(new_n1092), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1096), .A2(new_n996), .A3(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n257), .B1(new_n943), .B2(new_n780), .C1(new_n765), .C2(new_n239), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1132), .A2(new_n769), .B1(new_n785), .B2(new_n809), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n777), .B2(new_n1127), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT121), .Z(new_n1217));
  NAND2_X1  g1017(.A1(new_n783), .A2(G150), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1196), .A3(new_n1218), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1214), .B(new_n1219), .C1(G128), .C2(new_n789), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n776), .A2(new_n512), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n271), .B1(new_n377), .B2(new_n755), .C1(new_n798), .C2(new_n225), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n786), .A2(G283), .B1(G97), .B2(new_n781), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n766), .B2(new_n769), .C1(new_n821), .C2(new_n759), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1221), .A2(new_n1028), .A3(new_n1222), .A4(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n749), .B1(new_n1220), .B2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n736), .C1(new_n747), .C2(new_n860), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n203), .B2(new_n830), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1093), .B2(new_n735), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1213), .A2(new_n1229), .ZN(G381));
  NAND2_X1  g1030(.A1(new_n1171), .A2(new_n694), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1170), .A2(new_n1166), .A3(KEYINPUT120), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT120), .B1(new_n1170), .B2(new_n1166), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1154), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1231), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n735), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1207), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1236), .A2(new_n1238), .A3(G378), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n998), .A2(new_n1019), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT109), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n998), .A2(KEYINPUT109), .A3(new_n1019), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n958), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(G381), .A2(G384), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(G393), .A2(G396), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1244), .A2(new_n1080), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT122), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1239), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(G378), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1180), .A2(new_n1251), .A3(new_n1210), .ZN(new_n1252));
  OAI21_X1  g1052(.A(KEYINPUT122), .B1(new_n1252), .B2(new_n1247), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(G407));
  NAND2_X1  g1054(.A1(new_n665), .A2(G213), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT123), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1239), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(G407), .A2(G213), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT124), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(G407), .A2(KEYINPUT124), .A3(G213), .A4(new_n1257), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(G409));
  NOR3_X1   g1062(.A1(new_n1175), .A2(new_n1176), .A3(new_n734), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1179), .B2(new_n996), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(G378), .A2(new_n1208), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1256), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(G378), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT60), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1096), .B(new_n694), .C1(new_n1268), .C2(new_n1212), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1212), .A2(new_n1268), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1229), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(G384), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1266), .A2(new_n1267), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT62), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT125), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1256), .A2(G2897), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1271), .A2(new_n839), .A3(new_n846), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G384), .B(new_n1229), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1281), .A2(new_n1276), .A3(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1276), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1278), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1251), .B1(new_n1180), .B2(new_n1210), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n996), .B(new_n1154), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1263), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1265), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1256), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1280), .B(new_n1285), .C1(new_n1286), .C2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1266), .A2(new_n1267), .A3(new_n1293), .A4(new_n1272), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1274), .A2(new_n1275), .A3(new_n1292), .A4(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G387), .A2(G390), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n959), .B(new_n1080), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(G393), .B(G396), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1296), .A2(new_n1297), .A3(new_n1299), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1301), .A2(KEYINPUT126), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT126), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1295), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1292), .A2(KEYINPUT63), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1273), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1296), .A2(new_n1297), .A3(new_n1299), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1299), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1266), .A2(new_n1267), .A3(KEYINPUT63), .A4(new_n1272), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1311), .A2(new_n1312), .A3(new_n1275), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1308), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1306), .A2(new_n1314), .ZN(G405));
  NAND2_X1  g1115(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1316), .A2(KEYINPUT127), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1267), .A2(new_n1252), .A3(new_n1272), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1272), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n1239), .B2(new_n1286), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1316), .A2(KEYINPUT127), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1317), .A2(new_n1318), .A3(new_n1320), .A4(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1318), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(KEYINPUT127), .A3(new_n1316), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(G402));
endmodule


