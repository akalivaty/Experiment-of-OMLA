//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G257), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n210), .B(new_n211), .C1(new_n202), .C2(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n209), .B(new_n219), .C1(G87), .C2(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G1), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(KEYINPUT1), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OR3_X1    g0024(.A1(new_n220), .A2(KEYINPUT1), .A3(new_n223), .ZN(new_n225));
  INV_X1    g0025(.A(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(G20), .ZN(new_n231));
  INV_X1    g0031(.A(G68), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n217), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND4_X1  g0035(.A1(new_n231), .A2(G50), .A3(new_n233), .A4(new_n235), .ZN(new_n236));
  AND4_X1   g0036(.A1(new_n224), .A2(new_n225), .A3(new_n230), .A4(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n218), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(new_n221), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n202), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  AND3_X1   g0056(.A1(new_n253), .A2(new_n234), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT68), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n221), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n256), .A2(new_n234), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT65), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  OR2_X1    g0068(.A1(KEYINPUT8), .A2(G58), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT8), .A2(G58), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G150), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n222), .A2(new_n273), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n268), .A2(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(G20), .B2(new_n203), .ZN(new_n276));
  INV_X1    g0076(.A(new_n261), .ZN(new_n277));
  OAI221_X1 g0077(.A(new_n255), .B1(new_n202), .B2(new_n263), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n273), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G222), .A2(G1698), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(G223), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n234), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n286), .B(new_n288), .C1(G77), .C2(new_n282), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT67), .B(G45), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n221), .B(G274), .C1(new_n290), .C2(G41), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  OAI211_X1 g0092(.A(G1), .B(G13), .C1(new_n273), .C2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n221), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n289), .B(new_n291), .C1(new_n212), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n278), .B(new_n298), .C1(G179), .C2(new_n296), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT9), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n278), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n296), .A2(G200), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n278), .A2(new_n301), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n296), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n300), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NOR2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  OAI211_X1 g0112(.A(G232), .B(new_n284), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT69), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT69), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n282), .A2(new_n315), .A3(G232), .A4(new_n284), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n311), .A2(new_n312), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G107), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n282), .A2(G238), .A3(G1698), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n314), .A2(new_n316), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n288), .ZN(new_n321));
  INV_X1    g0121(.A(G244), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n291), .B1(new_n322), .B2(new_n295), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n297), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n327));
  NOR2_X1   g0127(.A1(G20), .A2(G33), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT70), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n269), .A2(new_n329), .A3(new_n270), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n231), .A2(G77), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n273), .B1(new_n264), .B2(new_n266), .ZN(new_n333));
  XOR2_X1   g0133(.A(KEYINPUT15), .B(G87), .Z(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n261), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n277), .A2(G77), .A3(new_n259), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n253), .A2(G77), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n323), .B1(new_n320), .B2(new_n288), .ZN(new_n342));
  INV_X1    g0142(.A(G179), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n326), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(G190), .ZN(new_n346));
  INV_X1    g0146(.A(G200), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n342), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n345), .B1(new_n348), .B2(new_n341), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n310), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n218), .A2(G1698), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n352), .B1(G226), .B2(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n353));
  AND2_X1   g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n293), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n221), .A2(G274), .ZN(new_n357));
  INV_X1    g0157(.A(new_n290), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n357), .B1(new_n358), .B2(new_n292), .ZN(new_n359));
  INV_X1    g0159(.A(G238), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n295), .A2(new_n360), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n356), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT13), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR4_X1   g0164(.A1(new_n356), .A2(new_n359), .A3(new_n361), .A4(KEYINPUT13), .ZN(new_n365));
  OAI21_X1  g0165(.A(G169), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT14), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n364), .A2(new_n365), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G179), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(G169), .C1(new_n364), .C2(new_n365), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n333), .A2(G77), .B1(G50), .B2(new_n328), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n232), .A2(G20), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n277), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT11), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n254), .A2(new_n232), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT12), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n277), .A2(G68), .A3(new_n259), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n372), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n368), .A2(G190), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n384), .B(new_n381), .C1(new_n347), .C2(new_n368), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT71), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G58), .A2(G68), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n222), .B1(new_n233), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G159), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n274), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n388), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n389), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n394), .B2(new_n201), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n328), .A2(G159), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(KEYINPUT71), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n267), .A2(new_n317), .A3(KEYINPUT7), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n280), .A2(new_n222), .A3(new_n281), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n232), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n387), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n267), .A2(new_n317), .A3(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n400), .A2(KEYINPUT7), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(G68), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(KEYINPUT16), .A3(new_n393), .A4(new_n397), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n408), .A3(new_n261), .ZN(new_n409));
  MUX2_X1   g0209(.A(new_n263), .B(new_n253), .S(new_n271), .Z(new_n410));
  NOR2_X1   g0210(.A1(new_n295), .A2(new_n218), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(G223), .A2(G1698), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n317), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n212), .A2(G1698), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n414), .A2(new_n415), .B1(G33), .B2(G87), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n291), .B(new_n412), .C1(new_n416), .C2(new_n293), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G200), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n282), .B(new_n415), .C1(G223), .C2(G1698), .ZN(new_n419));
  INV_X1    g0219(.A(G87), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(new_n273), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n288), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n422), .A2(G190), .A3(new_n291), .A4(new_n412), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n409), .A2(new_n410), .A3(new_n418), .A4(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT17), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT72), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT18), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n409), .A2(new_n410), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n422), .A2(G179), .A3(new_n291), .A4(new_n412), .ZN(new_n429));
  INV_X1    g0229(.A(new_n417), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n429), .B1(new_n430), .B2(new_n297), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n427), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT72), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n428), .A2(new_n431), .A3(new_n427), .A4(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n425), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  XOR2_X1   g0237(.A(new_n437), .B(KEYINPUT73), .Z(new_n438));
  AND3_X1   g0238(.A1(new_n351), .A2(new_n386), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n334), .A2(new_n253), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT19), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT76), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT19), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n445), .A3(new_n354), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n267), .ZN(new_n447));
  NOR3_X1   g0247(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n267), .A2(G33), .A3(G97), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n443), .A2(new_n445), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n267), .A2(new_n282), .A3(G68), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n441), .B1(new_n455), .B2(new_n261), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n221), .A2(G33), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n277), .A2(KEYINPUT74), .A3(new_n253), .A4(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n253), .A2(new_n457), .A3(new_n234), .A4(new_n256), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT74), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n334), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n360), .A2(new_n284), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n322), .A2(G1698), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n464), .B(new_n465), .C1(new_n311), .C2(new_n312), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G116), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n293), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n221), .A2(G45), .A3(G274), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n221), .A2(G45), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(G250), .C1(new_n287), .C2(new_n234), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n468), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n456), .A2(new_n463), .B1(new_n474), .B2(new_n297), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n343), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n420), .B1(new_n458), .B2(new_n461), .ZN(new_n477));
  AOI211_X1 g0277(.A(new_n441), .B(new_n477), .C1(new_n261), .C2(new_n455), .ZN(new_n478));
  NOR4_X1   g0278(.A1(new_n468), .A2(new_n305), .A3(new_n472), .A4(new_n469), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(G200), .B2(new_n474), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n475), .A2(new_n476), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n207), .B1(new_n458), .B2(new_n461), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n399), .A2(new_n402), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G107), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n328), .A2(G77), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT6), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n207), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(G97), .A2(G107), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(KEYINPUT6), .A3(G97), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n267), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n484), .A2(new_n485), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n482), .B1(new_n494), .B2(new_n261), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n253), .A2(G97), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(G244), .B(new_n284), .C1(new_n311), .C2(new_n312), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n282), .A2(KEYINPUT4), .A3(G244), .A4(new_n284), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n282), .A2(G250), .A3(G1698), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n288), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT75), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(G41), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n292), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n292), .A2(KEYINPUT5), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n470), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n288), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n221), .B(G45), .C1(new_n292), .C2(KEYINPUT5), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n508), .B2(new_n509), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n513), .A2(G257), .B1(G274), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n505), .A2(new_n305), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(G200), .B1(new_n505), .B2(new_n516), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n495), .B(new_n497), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n482), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n487), .B1(new_n399), .B2(new_n402), .ZN(new_n521));
  INV_X1    g0321(.A(new_n485), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n521), .A2(new_n522), .A3(new_n492), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n520), .B(new_n497), .C1(new_n523), .C2(new_n277), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n505), .A2(new_n516), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n297), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n505), .A2(new_n343), .A3(new_n516), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n481), .A2(KEYINPUT77), .A3(new_n519), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n267), .A2(new_n282), .A3(G87), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT22), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(KEYINPUT81), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT23), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n264), .A2(new_n266), .A3(new_n535), .A4(new_n487), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n222), .A2(G33), .A3(G116), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT23), .B1(new_n222), .B2(G107), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n267), .A2(new_n282), .A3(G87), .A4(new_n532), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n534), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n534), .A2(new_n539), .A3(KEYINPUT24), .A4(new_n540), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n261), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n462), .A2(G107), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n253), .A2(G107), .ZN(new_n547));
  XNOR2_X1  g0347(.A(KEYINPUT82), .B(KEYINPUT25), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n513), .A2(G264), .ZN(new_n551));
  OR2_X1    g0351(.A1(G250), .A2(G1698), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n208), .A2(G1698), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n552), .B(new_n553), .C1(new_n311), .C2(new_n312), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT83), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G294), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n551), .B1(new_n559), .B2(new_n288), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n515), .A2(G274), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n343), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n554), .A2(new_n556), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT83), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n288), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n513), .A2(G264), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n297), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n550), .A2(new_n562), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n566), .A2(new_n305), .A3(new_n561), .A4(new_n567), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(KEYINPUT84), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n550), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n347), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(KEYINPUT84), .A3(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n529), .A2(new_n570), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n513), .A2(G270), .ZN(new_n578));
  OAI211_X1 g0378(.A(G264), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n579));
  OAI211_X1 g0379(.A(G257), .B(new_n284), .C1(new_n311), .C2(new_n312), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n280), .A2(G303), .A3(new_n281), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n288), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n578), .A2(new_n583), .A3(new_n561), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(new_n343), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n273), .A2(G97), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n265), .A2(G20), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n502), .B(new_n586), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(G116), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n256), .A2(new_n234), .B1(G20), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT20), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n589), .A2(KEYINPUT20), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT78), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n257), .A2(new_n597), .A3(G116), .A4(new_n457), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT78), .B1(new_n459), .B2(new_n590), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n254), .A2(new_n590), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n585), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT80), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n513), .A2(G270), .B1(G274), .B2(new_n515), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n297), .B1(new_n605), .B2(new_n583), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI211_X1 g0409(.A(KEYINPUT80), .B(KEYINPUT21), .C1(new_n602), .C2(new_n606), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n603), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n602), .A2(KEYINPUT21), .A3(new_n606), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT79), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT79), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n602), .A2(new_n614), .A3(new_n606), .A4(KEYINPUT21), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT77), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n519), .A2(new_n528), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n478), .A2(new_n480), .ZN(new_n620));
  INV_X1    g0420(.A(new_n441), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n333), .A2(G97), .B1(new_n443), .B2(new_n445), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n317), .A2(new_n231), .A3(new_n232), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n448), .B1(new_n446), .B2(new_n267), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n621), .B(new_n463), .C1(new_n625), .C2(new_n277), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n474), .A2(new_n297), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(new_n476), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n620), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n618), .B1(new_n619), .B2(new_n629), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n589), .A2(KEYINPUT20), .A3(new_n591), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT20), .B1(new_n589), .B2(new_n591), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n601), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n598), .A2(new_n599), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n584), .A2(G200), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n635), .B(new_n636), .C1(new_n305), .C2(new_n584), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n617), .A2(new_n630), .A3(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n440), .A2(new_n577), .A3(new_n638), .ZN(G372));
  INV_X1    g0439(.A(new_n383), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n345), .A2(KEYINPUT87), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT87), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n326), .A2(new_n642), .A3(new_n341), .A4(new_n344), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n385), .B(new_n425), .C1(new_n640), .C2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n428), .A2(new_n431), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT86), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT86), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n428), .A2(new_n431), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n647), .A2(KEYINPUT18), .A3(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n428), .A2(new_n431), .A3(new_n648), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n648), .B1(new_n428), .B2(new_n431), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n434), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n645), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n308), .A2(new_n309), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n300), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n584), .A2(G169), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n608), .B1(new_n635), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT80), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n607), .A2(new_n604), .A3(new_n608), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n613), .A2(new_n615), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n661), .A2(new_n570), .A3(new_n603), .A4(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n619), .B1(new_n573), .B2(new_n575), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT85), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n473), .B2(new_n347), .ZN(new_n666));
  INV_X1    g0466(.A(new_n479), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n462), .A2(G87), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n666), .A2(new_n456), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n473), .A2(new_n665), .A3(new_n347), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n628), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n663), .A2(new_n664), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT26), .B1(new_n629), .B2(new_n528), .ZN(new_n674));
  INV_X1    g0474(.A(new_n628), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n671), .A2(new_n528), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n673), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n656), .B1(new_n440), .B2(new_n680), .ZN(G369));
  INV_X1    g0481(.A(G330), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n659), .A2(new_n660), .B1(new_n585), .B2(new_n602), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n231), .A2(new_n226), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n221), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n635), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n683), .A2(new_n662), .A3(new_n637), .A4(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n692), .B1(new_n611), .B2(new_n616), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n682), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n570), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n550), .A2(new_n690), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n576), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n570), .A2(new_n690), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n699), .A2(new_n700), .B1(new_n617), .B2(new_n690), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT88), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n696), .A2(new_n701), .A3(KEYINPUT88), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n690), .B1(new_n683), .B2(new_n662), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT84), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n560), .A2(new_n707), .A3(new_n305), .A4(new_n561), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n546), .A3(new_n545), .A4(new_n549), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n574), .A2(KEYINPUT84), .A3(new_n571), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n698), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n570), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n700), .B1(new_n706), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n705), .A2(new_n713), .ZN(G399));
  NOR2_X1   g0514(.A1(new_n227), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G1), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n448), .A2(new_n590), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n233), .A2(G50), .ZN(new_n719));
  OAI22_X1  g0519(.A1(new_n717), .A2(new_n718), .B1(new_n719), .B2(new_n716), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n529), .A2(new_n570), .A3(new_n576), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n683), .A2(new_n662), .A3(new_n637), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n722), .A2(new_n723), .A3(new_n630), .A4(new_n691), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n566), .A2(new_n567), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n725), .A2(new_n343), .A3(new_n584), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n525), .A2(new_n474), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT89), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n568), .A2(new_n584), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n343), .A3(new_n525), .A4(new_n474), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n726), .B(new_n727), .C1(new_n729), .C2(KEYINPUT30), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n690), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT31), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n738), .A3(new_n690), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n682), .B1(new_n724), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT26), .B1(new_n671), .B2(new_n528), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n524), .A2(new_n527), .A3(new_n526), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n481), .A2(new_n677), .A3(new_n743), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n742), .A2(new_n744), .A3(new_n628), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n673), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT90), .B1(new_n746), .B2(new_n691), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT90), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n748), .B(new_n690), .C1(new_n673), .C2(new_n745), .ZN(new_n749));
  OAI21_X1  g0549(.A(KEYINPUT29), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n679), .A2(new_n691), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT29), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n741), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n721), .B1(new_n754), .B2(G1), .ZN(G364));
  AOI21_X1  g0555(.A(new_n234), .B1(G20), .B2(new_n297), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n267), .A2(G190), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G179), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n347), .ZN(new_n759));
  XNOR2_X1  g0559(.A(KEYINPUT33), .B(G317), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n759), .A2(new_n760), .B1(new_n763), .B2(G329), .ZN(new_n764));
  INV_X1    g0564(.A(G294), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n305), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n267), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G303), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n347), .A2(G179), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(G20), .A3(G190), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n764), .B1(new_n765), .B2(new_n767), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n267), .A2(new_n343), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G190), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n282), .B1(new_n774), .B2(G322), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n757), .A2(G179), .A3(new_n347), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n772), .A2(G190), .A3(G200), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT92), .ZN(new_n779));
  INV_X1    g0579(.A(G326), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n775), .B1(new_n776), .B2(new_n777), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n757), .A2(new_n769), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n771), .B(new_n781), .C1(G283), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n762), .A2(new_n391), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT32), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n787), .B1(new_n207), .B2(new_n767), .C1(new_n487), .C2(new_n782), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n786), .A2(KEYINPUT32), .B1(new_n202), .B2(new_n778), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n770), .A2(new_n420), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n317), .ZN(new_n791));
  INV_X1    g0591(.A(G77), .ZN(new_n792));
  INV_X1    g0592(.A(new_n774), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n791), .B1(new_n792), .B2(new_n777), .C1(new_n793), .C2(new_n217), .ZN(new_n794));
  INV_X1    g0594(.A(new_n759), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n232), .ZN(new_n796));
  NOR4_X1   g0596(.A1(new_n788), .A2(new_n789), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n756), .B1(new_n784), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n226), .A2(new_n273), .A3(KEYINPUT91), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT91), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G13), .B2(G33), .ZN(new_n801));
  AOI21_X1  g0601(.A(G20), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n756), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n227), .A2(new_n282), .ZN(new_n805));
  INV_X1    g0605(.A(G45), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n805), .B1(new_n719), .B2(new_n290), .C1(new_n251), .C2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(G116), .B2(new_n228), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n227), .A2(new_n317), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(G355), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n694), .A2(new_n695), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n802), .B(KEYINPUT93), .Z(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n798), .B1(new_n804), .B2(new_n810), .C1(new_n811), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n717), .B1(G45), .B2(new_n684), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n811), .A2(G330), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n696), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT94), .Z(G396));
  INV_X1    g0621(.A(new_n777), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G150), .A2(new_n759), .B1(new_n822), .B2(G159), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n778), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G143), .B2(new_n774), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT34), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n282), .B1(new_n762), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n782), .A2(new_n232), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n217), .B2(new_n767), .ZN(new_n832));
  INV_X1    g0632(.A(new_n770), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(G50), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G283), .A2(new_n759), .B1(new_n822), .B2(G116), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n420), .B2(new_n782), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n317), .B1(new_n207), .B2(new_n767), .C1(new_n793), .C2(new_n765), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n762), .A2(new_n776), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n778), .A2(new_n768), .B1(new_n487), .B2(new_n770), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n756), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n690), .A2(new_n341), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n644), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT95), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n350), .A2(new_n842), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT95), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n644), .A2(new_n847), .A3(new_n843), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n799), .A2(new_n801), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n756), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n792), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n841), .A2(new_n815), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT96), .Z(new_n856));
  NAND2_X1  g0656(.A1(new_n751), .A2(new_n850), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n679), .A2(new_n691), .A3(new_n849), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(new_n741), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n817), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n856), .A2(new_n861), .ZN(G384));
  INV_X1    g0662(.A(new_n688), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n428), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n424), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n647), .A3(new_n649), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n646), .A2(new_n864), .A3(new_n868), .A4(new_n424), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT98), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT37), .B1(new_n428), .B2(new_n431), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n872), .A2(KEYINPUT98), .A3(new_n424), .A4(new_n864), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n653), .A2(new_n650), .A3(new_n425), .ZN(new_n876));
  INV_X1    g0676(.A(new_n864), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(KEYINPUT97), .A2(KEYINPUT16), .ZN(new_n882));
  INV_X1    g0682(.A(new_n407), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n883), .B2(new_n398), .ZN(new_n884));
  OR2_X1    g0684(.A1(KEYINPUT97), .A2(KEYINPUT16), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n407), .A2(new_n393), .A3(new_n397), .A4(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n261), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n410), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n431), .B2(new_n863), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n868), .B1(new_n889), .B2(new_n424), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT98), .B1(new_n865), .B2(new_n872), .ZN(new_n892));
  INV_X1    g0692(.A(new_n873), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n888), .A2(new_n863), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n437), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(new_n897), .A3(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n881), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n382), .A2(new_n690), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n383), .A2(new_n385), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n372), .A2(new_n382), .A3(new_n690), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n849), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n724), .B2(new_n740), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT40), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT17), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n424), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n424), .A2(new_n908), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n909), .A2(new_n910), .A3(new_n432), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n895), .B1(new_n911), .B2(new_n436), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n890), .B1(new_n871), .B2(new_n873), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n912), .A2(new_n913), .A3(new_n880), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n894), .B2(new_n897), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n847), .B1(new_n644), .B2(new_n843), .ZN(new_n917));
  AOI211_X1 g0717(.A(KEYINPUT95), .B(new_n842), .C1(new_n641), .C2(new_n643), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n919), .A2(new_n846), .B1(new_n901), .B2(new_n902), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n638), .A2(new_n577), .A3(new_n690), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n737), .A2(new_n739), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n907), .B1(new_n916), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT99), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n724), .A2(new_n740), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(new_n920), .C1(new_n914), .C2(new_n915), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT99), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n928), .A3(new_n907), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n906), .B1(new_n925), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(new_n439), .A3(new_n926), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n905), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n880), .B1(new_n912), .B2(new_n913), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n898), .ZN(new_n934));
  AOI211_X1 g0734(.A(KEYINPUT99), .B(KEYINPUT40), .C1(new_n905), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n928), .B1(new_n927), .B2(new_n907), .ZN(new_n936));
  OAI211_X1 g0736(.A(G330), .B(new_n932), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n439), .A2(new_n741), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n931), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n439), .A2(new_n750), .A3(new_n753), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n941), .A2(new_n656), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n940), .B(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT39), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT38), .B1(new_n875), .B2(new_n878), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n944), .B1(new_n945), .B2(new_n914), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n383), .A2(new_n690), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n933), .A2(new_n898), .A3(KEYINPUT39), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n903), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n345), .A2(new_n690), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n950), .B1(new_n858), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n934), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n653), .A2(new_n650), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n688), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n943), .B(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n221), .B2(new_n684), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n490), .A2(new_n491), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n235), .B(new_n231), .C1(new_n960), .C2(KEYINPUT35), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n590), .B(new_n961), .C1(KEYINPUT35), .C2(new_n960), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT36), .Z(new_n963));
  NAND2_X1  g0763(.A1(new_n389), .A2(G77), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n719), .A2(new_n964), .B1(G50), .B2(new_n232), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(G1), .A3(new_n226), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n959), .A2(new_n963), .A3(new_n966), .ZN(G367));
  OAI211_X1 g0767(.A(new_n662), .B(new_n603), .C1(new_n609), .C2(new_n610), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n573), .A2(new_n575), .B1(new_n550), .B2(new_n690), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n570), .A4(new_n691), .ZN(new_n970));
  INV_X1    g0770(.A(new_n700), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n619), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n690), .A2(new_n524), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(KEYINPUT42), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n972), .A2(new_n973), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n974), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT42), .B1(new_n970), .B2(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n976), .B(new_n978), .C1(new_n528), .C2(new_n690), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n691), .A2(new_n478), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n675), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n671), .B2(new_n980), .ZN(new_n982));
  OR3_X1    g0782(.A1(new_n979), .A2(KEYINPUT43), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n743), .A2(new_n690), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n977), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n705), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n979), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n983), .A2(new_n987), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n987), .B1(new_n983), .B2(new_n991), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n715), .B(KEYINPUT41), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT102), .ZN(new_n997));
  INV_X1    g0797(.A(new_n970), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n712), .A2(new_n971), .B1(new_n968), .B2(new_n691), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n701), .A2(KEYINPUT102), .A3(new_n970), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n696), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT103), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n696), .A2(new_n701), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT103), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1000), .A2(new_n1001), .A3(new_n1006), .A4(new_n1002), .ZN(new_n1007));
  AND3_X1   g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT44), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n713), .B2(new_n985), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n972), .A2(KEYINPUT44), .A3(new_n986), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n970), .A2(new_n971), .A3(new_n985), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n713), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1012), .A2(new_n1017), .A3(KEYINPUT100), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n705), .B1(new_n1018), .B2(KEYINPUT101), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n696), .A2(new_n701), .A3(KEYINPUT88), .ZN(new_n1020));
  OAI21_X1  g0820(.A(KEYINPUT101), .B1(new_n1020), .B2(new_n702), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1021), .A2(KEYINPUT100), .B1(new_n1017), .B2(new_n1012), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1008), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n996), .B1(new_n1023), .B2(new_n754), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n221), .B1(new_n684), .B2(G45), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n994), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n282), .B1(new_n777), .B2(new_n202), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n778), .B(KEYINPUT92), .Z(new_n1029));
  AOI22_X1  g0829(.A1(new_n1029), .A2(G143), .B1(G150), .B2(new_n774), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n762), .A2(new_n824), .B1(new_n217), .B2(new_n770), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT105), .Z(new_n1032));
  NAND2_X1  g0832(.A1(new_n783), .A2(G77), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n767), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(G68), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1028), .B(new_n1036), .C1(G159), .C2(new_n759), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT106), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n795), .A2(new_n765), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n779), .A2(new_n776), .B1(new_n768), .B2(new_n793), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT104), .Z(new_n1041));
  AOI22_X1  g0841(.A1(new_n783), .A2(G97), .B1(G107), .B2(new_n1034), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n282), .B1(new_n763), .B2(G317), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n822), .A2(G283), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n833), .A2(G116), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT46), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1038), .B1(new_n1039), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT47), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n756), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n244), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n804), .B1(new_n1054), .B2(new_n805), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n334), .A2(new_n227), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n817), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT107), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1053), .A2(KEYINPUT107), .A3(new_n1057), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n813), .C2(new_n982), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1027), .A2(new_n1062), .ZN(G387));
  NAND2_X1  g0863(.A1(new_n926), .A2(G330), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n746), .A2(new_n691), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n748), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n746), .A2(KEYINPUT90), .A3(new_n691), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n752), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n753), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1008), .A2(new_n1070), .A3(new_n716), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G311), .A2(new_n759), .B1(new_n774), .B2(G317), .ZN(new_n1073));
  INV_X1    g0873(.A(G322), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1073), .B1(new_n768), .B2(new_n777), .C1(new_n779), .C2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT48), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1034), .A2(G283), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n833), .A2(G294), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1079), .A2(KEYINPUT49), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1079), .A2(KEYINPUT49), .B1(G116), .B2(new_n783), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n763), .A2(G326), .ZN(new_n1082));
  AND4_X1   g0882(.A1(new_n317), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n822), .A2(G68), .B1(new_n763), .B2(G150), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n391), .B2(new_n778), .C1(new_n202), .C2(new_n793), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1034), .A2(new_n334), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n792), .B2(new_n770), .C1(new_n207), .C2(new_n782), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n795), .A2(new_n271), .ZN(new_n1088));
  NOR4_X1   g0888(.A1(new_n1085), .A2(new_n317), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n756), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n327), .A2(new_n330), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(G50), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT108), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT50), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n806), .B1(new_n232), .B2(new_n792), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1094), .A2(new_n718), .A3(new_n1095), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n241), .A2(new_n358), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1097), .A2(new_n805), .B1(new_n718), .B2(new_n809), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1096), .A2(new_n1098), .B1(G107), .B2(new_n228), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n803), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n812), .B1(new_n699), .B2(new_n700), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1090), .A2(new_n815), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1008), .A2(new_n754), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1026), .B1(new_n1103), .B2(new_n715), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1072), .B(new_n1102), .C1(new_n1104), .C2(new_n1105), .ZN(G393));
  OAI21_X1  g0906(.A(new_n715), .B1(new_n1070), .B2(new_n1105), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1025), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n705), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1112), .A2(KEYINPUT109), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(KEYINPUT109), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1108), .A2(new_n1111), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n817), .B1(new_n986), .B2(new_n802), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n805), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n248), .A2(new_n1117), .B1(new_n207), .B2(new_n228), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n804), .B2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n793), .A2(new_n391), .B1(new_n272), .B2(new_n778), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT51), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n759), .A2(G50), .B1(new_n763), .B2(G143), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1034), .A2(G77), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n782), .B2(new_n420), .C1(new_n1091), .C2(new_n777), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n317), .B(new_n1124), .C1(G68), .C2(new_n833), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1121), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n778), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G311), .A2(new_n774), .B1(new_n1127), .B2(G317), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT52), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G303), .B2(new_n759), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n783), .A2(G107), .B1(G283), .B2(new_n833), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1131), .B(new_n317), .C1(new_n1074), .C2(new_n762), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT110), .Z(new_n1133));
  OAI211_X1 g0933(.A(new_n1130), .B(new_n1133), .C1(new_n765), .C2(new_n777), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n767), .A2(new_n590), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1126), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1119), .B1(new_n756), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1103), .A2(new_n716), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1115), .A2(new_n1140), .ZN(G390));
  NAND2_X1  g0941(.A1(new_n741), .A2(new_n920), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n947), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n899), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n849), .B1(new_n747), .B2(new_n749), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n952), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n1147), .B2(new_n903), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n858), .A2(new_n952), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n903), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1150), .A2(new_n1144), .B1(new_n946), .B2(new_n948), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1143), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n946), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n948), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1153), .A2(new_n1154), .B1(new_n953), .B2(new_n947), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n950), .B1(new_n1146), .B2(new_n952), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1142), .C1(new_n1156), .C2(new_n1145), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n941), .A2(new_n656), .A3(new_n938), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n903), .B1(new_n741), .B2(new_n849), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1149), .B1(new_n1143), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1142), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1163), .B2(new_n1147), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1159), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1158), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1152), .A2(new_n1157), .A3(new_n1159), .A4(new_n1164), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n715), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1152), .A2(new_n1157), .A3(new_n1026), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n851), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n793), .A2(new_n590), .B1(new_n207), .B2(new_n777), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n830), .B(new_n1171), .C1(G294), .C2(new_n763), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n759), .A2(G107), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n282), .B(new_n790), .C1(new_n1127), .C2(G283), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1172), .A2(new_n1123), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  XOR2_X1   g0975(.A(KEYINPUT54), .B(G143), .Z(new_n1176));
  NAND2_X1  g0976(.A1(new_n822), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n795), .B2(new_n824), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n317), .B(new_n1178), .C1(G125), .C2(new_n763), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1034), .A2(G159), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n774), .A2(G132), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1127), .A2(G128), .B1(new_n783), .B2(G50), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n770), .A2(new_n272), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n1185));
  XNOR2_X1  g0985(.A(new_n1184), .B(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1175), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n756), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n853), .A2(new_n271), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1170), .A2(new_n815), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1169), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1168), .A2(new_n1191), .ZN(G378));
  NAND2_X1  g0992(.A1(new_n278), .A2(new_n863), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n310), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n310), .A2(new_n1193), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1196), .B(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n937), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n925), .A2(new_n929), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1196), .B(new_n1197), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1201), .A2(G330), .A3(new_n932), .A4(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n957), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1200), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1204), .B1(new_n1200), .B2(new_n1203), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1026), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n817), .B1(new_n1199), .B2(new_n851), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n202), .B1(new_n311), .B2(G41), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n777), .A2(new_n824), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n774), .A2(G128), .B1(new_n833), .B2(new_n1176), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT112), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(G150), .C2(new_n1034), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1127), .A2(G125), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n828), .C2(new_n795), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n783), .A2(G159), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G41), .B1(new_n763), .B2(G124), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1216), .A2(new_n273), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1209), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n782), .A2(new_n217), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n774), .A2(G107), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n822), .A2(new_n334), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1034), .A2(G68), .B1(G77), .B2(new_n833), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n763), .A2(G283), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1222), .B(new_n1227), .C1(G116), .C2(new_n1127), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n759), .A2(G97), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n292), .A3(new_n317), .A4(new_n1229), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT58), .Z(new_n1231));
  OAI21_X1  g1031(.A(new_n756), .B1(new_n1221), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n853), .A2(new_n202), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1208), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT113), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1207), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1167), .A2(new_n1159), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT57), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n716), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1202), .B1(new_n930), .B2(G330), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n937), .A2(new_n1199), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n957), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1200), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(KEYINPUT114), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT114), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1205), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1239), .B1(new_n1167), .B2(new_n1159), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1236), .B1(new_n1240), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(G375));
  INV_X1    g1051(.A(new_n1159), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1164), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n995), .A3(new_n1165), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n817), .B1(new_n232), .B2(new_n853), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G116), .A2(new_n759), .B1(new_n822), .B2(G107), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(new_n1033), .A3(new_n1086), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n282), .B1(new_n763), .B2(G303), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n207), .B2(new_n770), .C1(new_n765), .C2(new_n778), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1258), .B(new_n1260), .C1(G283), .C2(new_n774), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT115), .Z(new_n1262));
  NOR2_X1   g1062(.A1(new_n778), .A2(new_n828), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n759), .A2(new_n1176), .B1(new_n822), .B2(G150), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1264), .B1(new_n202), .B2(new_n767), .C1(new_n824), .C2(new_n793), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1263), .B(new_n1265), .C1(G128), .C2(new_n763), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1266), .B(new_n282), .C1(new_n391), .C2(new_n770), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1262), .B1(new_n1222), .B2(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(KEYINPUT116), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n756), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1256), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT117), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n950), .A2(new_n851), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1272), .A2(new_n1273), .B1(new_n1026), .B2(new_n1164), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1255), .A2(new_n1274), .ZN(G381));
  NAND4_X1  g1075(.A1(new_n1027), .A2(new_n1062), .A3(new_n1115), .A4(new_n1140), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1102), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1108), .B2(new_n1008), .ZN(new_n1278));
  INV_X1    g1078(.A(G396), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n1072), .ZN(new_n1280));
  NOR4_X1   g1080(.A1(new_n1276), .A2(G381), .A3(new_n1280), .A4(G384), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT118), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G378), .A2(KEYINPUT119), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT119), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1168), .A2(new_n1284), .A3(new_n1191), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1250), .A2(new_n1286), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1282), .A2(new_n1287), .ZN(G407));
  OAI211_X1 g1088(.A(G407), .B(G213), .C1(G343), .C2(new_n1287), .ZN(G409));
  INV_X1    g1089(.A(KEYINPUT121), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1279), .B1(new_n1278), .B2(new_n1072), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1105), .B1(new_n1107), .B2(new_n1025), .ZN(new_n1292));
  NOR4_X1   g1092(.A1(new_n1292), .A2(G396), .A3(new_n1071), .A4(new_n1277), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1290), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G393), .A2(G396), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(KEYINPUT121), .A3(new_n1280), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(G390), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1276), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT123), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1299), .A2(KEYINPUT123), .A3(new_n1296), .A4(new_n1294), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1303));
  AND4_X1   g1103(.A1(new_n1027), .A2(new_n1062), .A3(new_n1115), .A4(new_n1140), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n1027), .A2(new_n1062), .B1(new_n1115), .B2(new_n1140), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT122), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1303), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1303), .B2(new_n1306), .ZN(new_n1309));
  OAI22_X1  g1109(.A1(new_n1300), .A2(new_n1302), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1310), .B(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(G213), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1313), .A2(G343), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1236), .ZN(new_n1315));
  AOI22_X1  g1115(.A1(new_n1243), .A2(new_n1244), .B1(new_n1159), .B2(new_n1167), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n715), .B1(new_n1316), .B2(KEYINPUT57), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1245), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G378), .B(new_n1315), .C1(new_n1317), .C2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1245), .A2(new_n1026), .A3(new_n1247), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1237), .B(new_n995), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1235), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1286), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1314), .B1(new_n1319), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT60), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n715), .B(new_n1165), .C1(new_n1254), .C2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT60), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1274), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(G384), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT62), .B1(new_n1324), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT125), .ZN(new_n1334));
  AOI22_X1  g1134(.A1(new_n1250), .A2(G378), .B1(new_n1286), .B2(new_n1322), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1334), .B1(new_n1335), .B2(new_n1314), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1314), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1337), .A2(KEYINPUT125), .A3(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1336), .A2(new_n1339), .ZN(new_n1340));
  AND2_X1   g1140(.A1(new_n1332), .A2(KEYINPUT62), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1333), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1332), .A2(G2897), .A3(new_n1314), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1314), .A2(G2897), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1344), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1336), .A2(new_n1339), .A3(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT61), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1312), .B1(new_n1342), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT124), .ZN(new_n1351));
  OAI21_X1  g1151(.A(KEYINPUT122), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1303), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT123), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1355), .B1(new_n1303), .B2(new_n1306), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1301), .ZN(new_n1357));
  AOI211_X1 g1157(.A(new_n1351), .B(KEYINPUT61), .C1(new_n1354), .C2(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(KEYINPUT124), .B1(new_n1310), .B2(new_n1348), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  XOR2_X1   g1160(.A(KEYINPUT120), .B(KEYINPUT63), .Z(new_n1361));
  AOI21_X1  g1161(.A(new_n1361), .B1(new_n1324), .B2(new_n1332), .ZN(new_n1362));
  AND2_X1   g1162(.A1(new_n1332), .A2(KEYINPUT63), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1362), .B1(new_n1340), .B2(new_n1363), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1346), .B1(new_n1314), .B2(new_n1335), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1360), .A2(new_n1364), .A3(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1350), .A2(new_n1366), .ZN(G405));
  AOI21_X1  g1167(.A(new_n1250), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1319), .ZN(new_n1369));
  OR3_X1    g1169(.A1(new_n1368), .A2(new_n1369), .A3(new_n1332), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n1332), .B1(new_n1368), .B2(new_n1369), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1372));
  OR2_X1    g1172(.A1(new_n1310), .A2(KEYINPUT127), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1310), .A2(KEYINPUT127), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1372), .A2(new_n1373), .A3(new_n1374), .ZN(new_n1375));
  NAND4_X1  g1175(.A1(new_n1370), .A2(KEYINPUT127), .A3(new_n1310), .A4(new_n1371), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1375), .A2(new_n1376), .ZN(G402));
endmodule


