//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT66), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(G116), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT2), .B(G113), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  AND3_X1   g010(.A1(new_n191), .A2(KEYINPUT67), .A3(new_n193), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT67), .B1(new_n191), .B2(new_n193), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n196), .B1(new_n199), .B2(new_n195), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT0), .B(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(G137), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n209), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n211), .A2(G137), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n213), .A2(G134), .ZN(new_n222));
  OAI21_X1  g036(.A(G131), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n202), .A3(new_n204), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT64), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n207), .A2(new_n229), .A3(new_n226), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n202), .A2(new_n204), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n232), .B1(new_n234), .B2(new_n225), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n224), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n220), .B1(new_n236), .B2(KEYINPUT65), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n233), .A2(G128), .B1(new_n202), .B2(new_n204), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n228), .B2(new_n230), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n238), .B1(new_n240), .B2(new_n224), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n200), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n229), .B1(new_n207), .B2(new_n226), .ZN(new_n243));
  AND4_X1   g057(.A1(new_n229), .A2(new_n226), .A3(new_n202), .A4(new_n204), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n235), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n224), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n196), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n194), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n191), .A2(KEYINPUT67), .A3(new_n193), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n195), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n219), .A2(new_n217), .ZN(new_n253));
  INV_X1    g067(.A(new_n209), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n247), .A2(new_n248), .A3(new_n252), .A4(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI211_X1 g071(.A(KEYINPUT69), .B(KEYINPUT28), .C1(new_n242), .C2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n245), .A2(KEYINPUT65), .A3(new_n246), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n241), .A2(new_n260), .A3(new_n255), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n252), .A2(new_n248), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n259), .B1(new_n263), .B2(new_n256), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n256), .B2(new_n259), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n258), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(G237), .A2(G953), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G210), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT27), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G101), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n241), .A2(new_n260), .A3(new_n255), .A4(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n219), .A2(new_n217), .ZN(new_n278));
  OAI22_X1  g092(.A1(new_n278), .A2(new_n209), .B1(new_n240), .B2(new_n224), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT30), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n200), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT68), .A2(KEYINPUT31), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n256), .A2(new_n272), .A3(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n274), .B(new_n275), .C1(new_n281), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(new_n280), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n262), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n274), .A2(new_n275), .ZN(new_n287));
  INV_X1    g101(.A(new_n283), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n267), .A2(new_n273), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(G472), .A2(G902), .ZN(new_n291));
  XOR2_X1   g105(.A(new_n291), .B(KEYINPUT70), .Z(new_n292));
  OAI21_X1  g106(.A(KEYINPUT32), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n294));
  INV_X1    g108(.A(new_n292), .ZN(new_n295));
  INV_X1    g109(.A(new_n266), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n242), .A2(new_n257), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n296), .B1(new_n297), .B2(new_n259), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n272), .B1(new_n298), .B2(new_n258), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n289), .A2(new_n284), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n294), .B(new_n295), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n263), .A2(new_n256), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n266), .B1(new_n303), .B2(KEYINPUT28), .ZN(new_n304));
  AOI211_X1 g118(.A(new_n265), .B(new_n259), .C1(new_n263), .C2(new_n256), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n272), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n281), .A2(new_n257), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n273), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT29), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n256), .A2(new_n259), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n279), .A2(new_n262), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT71), .A3(new_n256), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n279), .A2(new_n314), .A3(new_n262), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n311), .B1(new_n316), .B2(new_n259), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n272), .A2(KEYINPUT29), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G472), .B1(new_n309), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n302), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT9), .B(G234), .ZN(new_n322));
  OAI21_X1  g136(.A(G221), .B1(new_n322), .B2(G902), .ZN(new_n323));
  XOR2_X1   g137(.A(new_n323), .B(KEYINPUT76), .Z(new_n324));
  INV_X1    g138(.A(G469), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(new_n310), .ZN(new_n326));
  XNOR2_X1  g140(.A(G110), .B(G140), .ZN(new_n327));
  INV_X1    g141(.A(G227), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(G953), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n327), .B(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n331));
  INV_X1    g145(.A(G104), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(G107), .ZN(new_n333));
  INV_X1    g147(.A(G107), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT3), .A3(G104), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G101), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n334), .B2(G104), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n332), .A2(KEYINPUT77), .A3(G107), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n336), .A2(new_n337), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT78), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n339), .A2(new_n340), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n337), .A4(new_n336), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n336), .A2(new_n339), .A3(new_n340), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G101), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n342), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n337), .B1(new_n343), .B2(new_n336), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(new_n350), .B2(KEYINPUT79), .ZN(new_n351));
  AND4_X1   g165(.A1(KEYINPUT79), .A2(new_n346), .A3(new_n349), .A4(G101), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n254), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n334), .A2(G104), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n332), .A2(G107), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n337), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n342), .B2(new_n345), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n233), .A2(KEYINPUT80), .ZN(new_n359));
  OAI21_X1  g173(.A(G128), .B1(new_n233), .B2(KEYINPUT80), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n232), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n231), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n240), .A2(new_n364), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n354), .A2(new_n365), .A3(new_n278), .A4(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n353), .A2(new_n254), .B1(new_n358), .B2(new_n366), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n278), .B1(new_n370), .B2(new_n365), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n330), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n342), .A2(new_n345), .ZN(new_n373));
  INV_X1    g187(.A(new_n357), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n373), .A2(new_n374), .A3(new_n362), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n245), .B1(new_n373), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n253), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT12), .ZN(new_n378));
  INV_X1    g192(.A(new_n330), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT12), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n380), .B(new_n253), .C1(new_n375), .C2(new_n376), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n378), .A2(new_n368), .A3(new_n379), .A4(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(G902), .B1(new_n372), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n326), .B1(new_n383), .B2(new_n325), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n378), .A2(new_n368), .A3(new_n381), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n330), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n354), .A2(new_n365), .A3(new_n367), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n253), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n368), .A3(new_n379), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(G469), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n324), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G234), .ZN(new_n392));
  OAI21_X1  g206(.A(G217), .B1(new_n392), .B2(G902), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT72), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G125), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT16), .ZN(new_n398));
  XNOR2_X1  g212(.A(G125), .B(G140), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(KEYINPUT16), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G146), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n201), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT23), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT74), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT23), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT66), .B(G119), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n408), .B1(new_n409), .B2(G128), .ZN(new_n410));
  NAND2_X1  g224(.A1(KEYINPUT23), .A2(G119), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT73), .B1(new_n411), .B2(G128), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT73), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n413), .A2(new_n225), .A3(KEYINPUT23), .A4(G119), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G110), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n188), .A2(new_n190), .A3(G128), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n410), .A2(new_n415), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n418), .A2(KEYINPUT75), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n417), .B1(new_n187), .B2(G128), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT24), .B(G110), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n418), .B2(KEYINPUT75), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n403), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G125), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G140), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n397), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT16), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n201), .B1(new_n429), .B2(new_n398), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n401), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n410), .A2(new_n415), .A3(new_n417), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G110), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n431), .B(new_n433), .C1(new_n420), .C2(new_n421), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT22), .B(G137), .ZN(new_n435));
  INV_X1    g249(.A(G953), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(G221), .A3(G234), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n435), .B(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n424), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n424), .B2(new_n434), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT25), .B1(new_n441), .B2(new_n310), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT25), .ZN(new_n443));
  NOR4_X1   g257(.A1(new_n439), .A2(new_n440), .A3(new_n443), .A4(G902), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n395), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n393), .A2(new_n310), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n321), .A2(new_n391), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G110), .B(G122), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n353), .A2(new_n262), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT5), .B1(new_n197), .B2(new_n198), .ZN(new_n457));
  OAI21_X1  g271(.A(G113), .B1(new_n191), .B2(KEYINPUT5), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n196), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT81), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(new_n358), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n461), .B1(new_n460), .B2(new_n358), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n455), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT5), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n466), .B1(new_n250), .B2(new_n251), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n248), .B1(new_n467), .B2(new_n458), .ZN(new_n468));
  INV_X1    g282(.A(new_n358), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT81), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n470), .A2(new_n456), .A3(new_n454), .A4(new_n462), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n465), .A2(KEYINPUT6), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n240), .A2(new_n425), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n209), .A2(G125), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n436), .A2(G224), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n475), .B(new_n476), .Z(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n455), .C1(new_n463), .C2(new_n464), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n472), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT83), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n473), .A2(new_n474), .B1(new_n481), .B2(new_n476), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n476), .A2(KEYINPUT7), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n471), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT82), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n460), .B2(new_n358), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT82), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n459), .B1(new_n466), .B2(new_n194), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n358), .A2(new_n248), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n454), .B(KEYINPUT8), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n485), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n480), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G210), .B1(G237), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n480), .A2(new_n496), .A3(new_n494), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n453), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(G475), .A2(G902), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n268), .A2(G143), .A3(G214), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(G143), .B1(new_n268), .B2(G214), .ZN(new_n504));
  OAI211_X1 g318(.A(KEYINPUT18), .B(G131), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n427), .A2(G146), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n402), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n268), .A2(G214), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n203), .ZN(new_n509));
  NAND2_X1  g323(.A1(KEYINPUT18), .A2(G131), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n502), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n505), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT84), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT84), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n505), .A2(new_n507), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n509), .A2(new_n502), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G131), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n509), .A2(new_n215), .A3(new_n502), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(KEYINPUT17), .A3(G131), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n521), .A2(new_n430), .A3(new_n401), .A4(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(G113), .B(G122), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(new_n332), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n516), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n518), .A2(new_n520), .B1(new_n400), .B2(G146), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n399), .A2(KEYINPUT19), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n399), .A2(KEYINPUT19), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT85), .B1(new_n530), .B2(new_n201), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT85), .ZN(new_n532));
  AOI211_X1 g346(.A(new_n532), .B(G146), .C1(new_n528), .C2(new_n529), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n527), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n525), .B1(new_n534), .B2(new_n516), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n501), .B1(new_n526), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT20), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT20), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n538), .B(new_n501), .C1(new_n526), .C2(new_n535), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n225), .A2(G143), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT87), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n203), .A2(G128), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n211), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT88), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT88), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n542), .A2(new_n546), .A3(new_n211), .A4(new_n543), .ZN(new_n547));
  INV_X1    g361(.A(G122), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(G116), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n192), .A2(G122), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(new_n334), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT87), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n541), .B(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT13), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n543), .B(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G134), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n545), .A2(new_n547), .A3(new_n552), .A4(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n549), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT89), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n559), .B(new_n560), .C1(KEYINPUT14), .C2(new_n550), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n550), .A2(KEYINPUT14), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(new_n549), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT89), .B1(new_n559), .B2(KEYINPUT14), .ZN(new_n564));
  OAI211_X1 g378(.A(G107), .B(new_n561), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n551), .A2(new_n334), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n542), .A2(new_n211), .A3(new_n543), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n211), .B1(new_n542), .B2(new_n543), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n565), .B(new_n566), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n558), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G217), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n322), .A2(new_n571), .A3(G953), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT90), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n558), .A2(new_n569), .A3(new_n572), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n570), .A2(KEYINPUT90), .A3(new_n573), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n310), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G478), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT15), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n525), .B1(new_n516), .B2(new_n523), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n310), .B1(new_n526), .B2(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT86), .B(G475), .Z(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n581), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n577), .A2(new_n310), .A3(new_n578), .A4(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n540), .A2(new_n582), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G237), .ZN(new_n590));
  OAI211_X1 g404(.A(G902), .B(G953), .C1(new_n392), .C2(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(KEYINPUT91), .Z(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT21), .B(G898), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n436), .A2(G952), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n392), .B2(new_n590), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT92), .B1(new_n589), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n582), .A2(new_n588), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT92), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n537), .A2(new_n539), .B1(new_n584), .B2(new_n585), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n600), .A2(new_n601), .A3(new_n597), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n500), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n451), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n337), .ZN(G3));
  OAI21_X1  g421(.A(new_n273), .B1(new_n304), .B2(new_n305), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n289), .A2(new_n284), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n310), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n611), .A2(G472), .B1(new_n295), .B2(new_n610), .ZN(new_n612));
  INV_X1    g426(.A(new_n382), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n379), .B1(new_n388), .B2(new_n368), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n325), .B(new_n310), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n326), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n390), .ZN(new_n617));
  INV_X1    g431(.A(new_n324), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n612), .A2(new_n617), .A3(new_n618), .A4(new_n450), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT93), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n579), .A2(new_n580), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n577), .A2(new_n622), .A3(new_n578), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n574), .A2(KEYINPUT33), .A3(new_n576), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n623), .A2(G478), .A3(new_n310), .A4(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n602), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n480), .A2(new_n496), .A3(new_n494), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n496), .B1(new_n480), .B2(new_n494), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n452), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n620), .A2(new_n597), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND2_X1  g447(.A1(new_n582), .A2(new_n588), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n597), .B(KEYINPUT94), .Z(new_n635));
  AND3_X1   g449(.A1(new_n634), .A2(new_n602), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n620), .A2(new_n500), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  INV_X1    g453(.A(KEYINPUT95), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n441), .A2(KEYINPUT25), .A3(new_n310), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n424), .A2(new_n434), .ZN(new_n642));
  INV_X1    g456(.A(new_n438), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n424), .A2(new_n434), .A3(new_n438), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n310), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n443), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n394), .B1(new_n641), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n643), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n642), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n447), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n640), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n445), .A2(KEYINPUT95), .A3(new_n651), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n391), .A2(new_n612), .A3(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(new_n605), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  NAND2_X1  g473(.A1(new_n500), .A2(new_n321), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n634), .A2(new_n602), .ZN(new_n662));
  INV_X1    g476(.A(new_n596), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n592), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n661), .A2(new_n391), .A3(new_n655), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  NAND2_X1  g482(.A1(new_n498), .A2(new_n499), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT38), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n391), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n665), .B(KEYINPUT39), .Z(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  OR3_X1    g489(.A1(new_n673), .A2(KEYINPUT40), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT40), .B1(new_n673), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n316), .A2(new_n273), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n272), .B1(new_n281), .B2(new_n257), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n310), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n293), .A2(new_n301), .B1(G472), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n600), .A2(new_n602), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n452), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n681), .A2(new_n655), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n672), .A2(new_n676), .A3(new_n677), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  INV_X1    g500(.A(new_n626), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n665), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n391), .A3(new_n655), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n660), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n201), .ZN(G48));
  AOI21_X1  g505(.A(new_n449), .B1(new_n302), .B2(new_n320), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n372), .A2(new_n382), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n310), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n615), .A3(new_n323), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n630), .A2(new_n597), .A3(new_n692), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT96), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n698), .B(new_n700), .ZN(G15));
  NAND4_X1  g515(.A1(new_n692), .A2(new_n697), .A3(new_n500), .A4(new_n636), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  AOI22_X1  g517(.A1(new_n302), .A2(new_n320), .B1(new_n599), .B2(new_n603), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(new_n500), .A3(new_n655), .A4(new_n697), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  OAI211_X1 g520(.A(new_n682), .B(new_n452), .C1(new_n627), .C2(new_n628), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n615), .A2(new_n695), .A3(new_n323), .A4(new_n635), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n317), .A2(new_n273), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n292), .B1(new_n710), .B2(new_n609), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT97), .ZN(new_n712));
  AOI21_X1  g526(.A(G902), .B1(new_n608), .B2(new_n609), .ZN(new_n713));
  INV_X1    g527(.A(G472), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI211_X1 g529(.A(KEYINPUT97), .B(G472), .C1(new_n290), .C2(G902), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n711), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n708), .A2(new_n709), .A3(new_n450), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  AND2_X1   g533(.A1(new_n697), .A2(new_n500), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n715), .A2(new_n716), .ZN(new_n721));
  INV_X1    g535(.A(new_n711), .ZN(new_n722));
  AND4_X1   g536(.A1(KEYINPUT98), .A2(new_n721), .A3(new_n655), .A4(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT98), .B1(new_n717), .B2(new_n655), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n688), .B(new_n720), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  INV_X1    g540(.A(new_n323), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n386), .A2(new_n389), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT99), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT99), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n389), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(G469), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n727), .B1(new_n732), .B2(new_n384), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n627), .A2(new_n628), .A3(new_n453), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n692), .A2(new_n688), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT100), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n735), .A2(KEYINPUT100), .A3(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n215), .ZN(G33));
  NAND4_X1  g555(.A1(new_n692), .A2(new_n666), .A3(new_n733), .A4(new_n734), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  INV_X1    g557(.A(KEYINPUT102), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n729), .A2(KEYINPUT45), .A3(new_n731), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n325), .B1(new_n728), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n326), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  OR3_X1    g562(.A1(new_n748), .A2(KEYINPUT101), .A3(KEYINPUT46), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT101), .B1(new_n748), .B2(KEYINPUT46), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(KEYINPUT46), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n749), .A2(new_n615), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n323), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n744), .B1(new_n753), .B2(new_n675), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n752), .A2(KEYINPUT102), .A3(new_n323), .A4(new_n674), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n655), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n625), .A2(new_n621), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n759), .B2(new_n602), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n759), .A2(new_n758), .A3(new_n602), .ZN(new_n761));
  OR4_X1    g575(.A1(new_n612), .A2(new_n757), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n734), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n756), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  INV_X1    g583(.A(new_n321), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n770), .A2(new_n449), .A3(new_n688), .A4(new_n734), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n753), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n752), .A2(KEYINPUT47), .A3(new_n323), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n396), .ZN(G42));
  XNOR2_X1  g590(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n696), .A2(new_n452), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT114), .B1(new_n671), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n669), .A2(new_n670), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT38), .B1(new_n498), .B2(new_n499), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n778), .B(KEYINPUT114), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n761), .A2(new_n760), .A3(new_n596), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n783), .A2(new_n450), .A3(new_n717), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n779), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT116), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n786), .B1(new_n779), .B2(new_n785), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT115), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n696), .A2(new_n669), .A3(new_n453), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n663), .A3(new_n450), .A4(new_n681), .ZN(new_n794));
  INV_X1    g608(.A(new_n602), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n794), .A2(new_n795), .A3(new_n759), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n723), .A2(new_n724), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n793), .A2(new_n783), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT118), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT118), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n774), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT47), .B1(new_n752), .B2(new_n323), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n695), .A2(new_n615), .A3(new_n324), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT113), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n784), .A2(new_n734), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n802), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n777), .B1(new_n792), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n595), .B1(new_n794), .B2(new_n687), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n798), .A2(new_n692), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT48), .Z(new_n813));
  AOI211_X1 g627(.A(new_n811), .B(new_n813), .C1(new_n720), .C2(new_n784), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n773), .A2(new_n816), .A3(new_n774), .A4(new_n805), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n734), .A3(new_n784), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n803), .A2(new_n804), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n816), .B1(new_n819), .B2(new_n805), .ZN(new_n820));
  OAI211_X1 g634(.A(KEYINPUT51), .B(new_n802), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n777), .A2(KEYINPUT117), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n821), .A2(new_n822), .B1(new_n791), .B2(new_n788), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n815), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n665), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n445), .A2(new_n651), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT106), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n445), .A2(KEYINPUT106), .A3(new_n651), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n680), .A2(G472), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n302), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n733), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT107), .B1(new_n833), .B2(new_n707), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n730), .B1(new_n386), .B2(new_n389), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n389), .A2(new_n730), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n835), .A2(new_n836), .A3(new_n325), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n615), .A2(new_n616), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n323), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n681), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT107), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n841), .A3(new_n708), .A4(new_n830), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n834), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n690), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n667), .A3(new_n844), .A4(new_n725), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n690), .B1(new_n834), .B2(new_n842), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(KEYINPUT52), .A3(new_n667), .A4(new_n725), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n733), .A2(new_n734), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n688), .B(new_n851), .C1(new_n723), .C2(new_n724), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n600), .A2(new_n602), .A3(new_n825), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n302), .B2(new_n320), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n391), .A3(new_n655), .A4(new_n734), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n742), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT105), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT105), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n852), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n705), .A2(new_n718), .A3(new_n698), .A4(new_n702), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n740), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n669), .A2(new_n452), .A3(new_n626), .A4(new_n635), .ZN(new_n864));
  OAI22_X1  g678(.A1(new_n451), .A2(new_n605), .B1(new_n864), .B2(new_n619), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n669), .A2(new_n452), .A3(new_n636), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n656), .A2(new_n605), .B1(new_n619), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(KEYINPUT104), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT104), .ZN(new_n869));
  OAI221_X1 g683(.A(new_n869), .B1(new_n619), .B2(new_n866), .C1(new_n605), .C2(new_n656), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n861), .A2(new_n863), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT53), .B1(new_n850), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n852), .A2(new_n856), .A3(new_n859), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n859), .B1(new_n852), .B2(new_n856), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n735), .A2(KEYINPUT100), .A3(KEYINPUT42), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT42), .B1(new_n735), .B2(KEYINPUT100), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n698), .A2(new_n705), .A3(new_n718), .A4(new_n702), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n868), .A3(new_n880), .A4(new_n870), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n847), .A2(KEYINPUT108), .A3(new_n849), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT108), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n845), .A2(new_n884), .A3(new_n846), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n882), .A2(new_n883), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n873), .A2(new_n887), .A3(KEYINPUT54), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT109), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n873), .A2(new_n887), .A3(KEYINPUT109), .A4(KEYINPUT54), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n886), .B1(new_n850), .B2(new_n872), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT110), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n847), .A2(new_n849), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n882), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT110), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT111), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n863), .A2(new_n898), .B1(new_n858), .B2(new_n860), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n868), .A2(KEYINPUT53), .A3(new_n870), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n879), .A2(new_n880), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(KEYINPUT111), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n883), .A2(new_n899), .A3(new_n902), .A4(new_n885), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n894), .A2(new_n897), .A3(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n890), .B(new_n891), .C1(new_n904), .C2(KEYINPUT54), .ZN(new_n905));
  OAI22_X1  g719(.A1(new_n824), .A2(new_n905), .B1(G952), .B2(G953), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n695), .A2(new_n615), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT49), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n602), .A3(new_n759), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(KEYINPUT49), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n832), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n450), .A2(new_n452), .A3(new_n618), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT103), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n671), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n906), .A2(new_n914), .ZN(G75));
  NAND3_X1  g729(.A1(new_n904), .A2(G210), .A3(G902), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n472), .A2(new_n479), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n477), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT55), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n920), .B1(new_n916), .B2(new_n917), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n436), .A2(G952), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G51));
  XNOR2_X1  g738(.A(new_n326), .B(KEYINPUT57), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n883), .A2(new_n885), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n871), .B(KEYINPUT53), .C1(new_n863), .C2(new_n898), .ZN(new_n928));
  OAI22_X1  g742(.A1(new_n901), .A2(KEYINPUT111), .B1(new_n874), .B2(new_n875), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n892), .A2(new_n893), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n926), .B1(new_n931), .B2(new_n897), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n903), .B1(new_n896), .B2(KEYINPUT110), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n893), .B(KEYINPUT53), .C1(new_n882), .C2(new_n895), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT54), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n925), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n693), .B(KEYINPUT120), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n904), .A2(G902), .A3(new_n745), .A4(new_n747), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n923), .B1(new_n938), .B2(new_n939), .ZN(G54));
  NAND4_X1  g754(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n526), .A2(new_n535), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n943), .A2(new_n944), .A3(new_n923), .ZN(G60));
  AND2_X1   g759(.A1(new_n623), .A2(new_n624), .ZN(new_n946));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT59), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n905), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n949), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n931), .A2(new_n926), .A3(new_n897), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n950), .A2(new_n923), .A3(new_n954), .ZN(G63));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT60), .Z(new_n957));
  OAI211_X1 g771(.A(new_n650), .B(new_n957), .C1(new_n933), .C2(new_n934), .ZN(new_n958));
  INV_X1    g772(.A(new_n923), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n441), .B1(new_n904), .B2(new_n957), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT121), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n962), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n965), .B(new_n964), .C1(new_n960), .C2(new_n961), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(G66));
  INV_X1    g783(.A(new_n593), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n436), .B1(new_n970), .B2(G224), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n871), .A2(new_n880), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n436), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n918), .B1(G898), .B2(new_n436), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n973), .B(new_n974), .Z(G69));
  INV_X1    g789(.A(new_n692), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n734), .A2(new_n391), .A3(new_n674), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n976), .B(new_n977), .C1(new_n687), .C2(new_n662), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n775), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n725), .A2(new_n667), .A3(new_n844), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n685), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n979), .A2(new_n983), .A3(new_n768), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n436), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n285), .B(new_n530), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n976), .A2(new_n707), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n756), .B1(new_n767), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n879), .A2(new_n742), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n775), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n991), .A2(new_n993), .A3(new_n981), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n994), .A2(G953), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n988), .B1(G900), .B2(G953), .ZN(new_n996));
  AOI22_X1  g810(.A1(new_n989), .A2(KEYINPUT122), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT124), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n328), .B2(new_n664), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT123), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n987), .B1(new_n985), .B2(new_n436), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT122), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1000), .A2(new_n998), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n1000), .A2(new_n998), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1003), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n996), .B1(new_n994), .B2(G953), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n1005), .B(new_n1006), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n1004), .A2(new_n1010), .ZN(G72));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  AND3_X1   g827(.A1(new_n308), .A2(new_n679), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n873), .A2(new_n887), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT125), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1013), .B1(new_n985), .B2(new_n972), .ZN(new_n1018));
  INV_X1    g832(.A(new_n679), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1013), .B1(new_n994), .B2(new_n972), .ZN(new_n1021));
  INV_X1    g835(.A(new_n308), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n923), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1017), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(KEYINPUT126), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT126), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n1017), .A2(new_n1026), .A3(new_n1023), .A4(new_n1020), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1025), .A2(new_n1027), .ZN(G57));
endmodule


