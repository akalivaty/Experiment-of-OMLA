//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n188), .B(new_n190), .Z(new_n191));
  INV_X1    g005(.A(G131), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G134), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT65), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n193), .B(new_n194), .C1(new_n196), .C2(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n193), .B1(G134), .B2(new_n194), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n197), .A2(KEYINPUT65), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n195), .A2(G134), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G137), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n192), .B1(new_n202), .B2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(G137), .B1(new_n203), .B2(new_n204), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n200), .B1(new_n207), .B2(new_n193), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n192), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT68), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n205), .ZN(new_n212));
  OAI21_X1  g026(.A(G131), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT65), .B(G134), .ZN(new_n215));
  AOI21_X1  g029(.A(G131), .B1(new_n215), .B2(G137), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n202), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT3), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT77), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G107), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(G104), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT3), .ZN(new_n227));
  AOI21_X1  g041(.A(G101), .B1(new_n219), .B2(G107), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n226), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n222), .A2(new_n224), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n219), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n229), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT64), .B(G143), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(G146), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(KEYINPUT64), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  AOI21_X1  g056(.A(G146), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n244));
  OAI21_X1  g058(.A(G128), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n242), .A3(G146), .ZN(new_n247));
  INV_X1    g061(.A(new_n236), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n234), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT77), .B(G107), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n226), .B1(new_n253), .B2(G104), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT3), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(G104), .B2(new_n221), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n253), .B2(new_n220), .ZN(new_n257));
  AOI22_X1  g071(.A1(G101), .A2(new_n254), .B1(new_n257), .B2(new_n228), .ZN(new_n258));
  OAI21_X1  g072(.A(G128), .B1(new_n236), .B2(new_n244), .ZN(new_n259));
  INV_X1    g073(.A(G146), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n259), .B1(new_n243), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n251), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n211), .B(new_n218), .C1(new_n252), .C2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n234), .A2(new_n262), .A3(new_n251), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n247), .A2(new_n248), .A3(new_n250), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n239), .B2(new_n245), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n269), .B2(new_n234), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n206), .A2(new_n210), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(new_n266), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n265), .A2(new_n266), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT10), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n269), .B2(new_n234), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT78), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n234), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n229), .B(KEYINPUT78), .C1(new_n232), .C2(new_n233), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n274), .B1(new_n262), .B2(new_n251), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n261), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n281), .B1(new_n237), .B2(G146), .ZN(new_n282));
  AND2_X1   g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT0), .A2(G128), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n282), .A2(new_n285), .B1(new_n238), .B2(new_n283), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n219), .A2(G107), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n225), .A2(new_n227), .A3(new_n287), .ZN(new_n288));
  AOI22_X1  g102(.A1(KEYINPUT4), .A2(new_n229), .B1(new_n288), .B2(G101), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n288), .A2(KEYINPUT4), .A3(G101), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n275), .A2(new_n280), .A3(new_n291), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n206), .A2(new_n210), .A3(KEYINPUT68), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n214), .B1(new_n213), .B2(new_n217), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n191), .B1(new_n273), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n191), .ZN(new_n298));
  OAI211_X1 g112(.A(KEYINPUT79), .B(new_n298), .C1(new_n292), .C2(new_n295), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n292), .A2(new_n295), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n211), .A2(new_n218), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n302), .A2(new_n280), .A3(new_n275), .A4(new_n291), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT79), .B1(new_n303), .B2(new_n298), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n297), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT80), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT80), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n297), .B(new_n307), .C1(new_n301), .C2(new_n304), .ZN(new_n308));
  AOI21_X1  g122(.A(G902), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G469), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n187), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n308), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n298), .B1(new_n292), .B2(new_n295), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT79), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n300), .A3(new_n299), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n307), .B1(new_n317), .B2(new_n297), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n312), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT81), .A3(G469), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n273), .A2(new_n314), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n298), .B1(new_n300), .B2(new_n303), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n310), .B(new_n312), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n311), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT88), .ZN(new_n325));
  OAI21_X1  g139(.A(G210), .B1(G237), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G116), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT66), .B1(new_n328), .B2(G119), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT66), .ZN(new_n330));
  INV_X1    g144(.A(G119), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(G116), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(G119), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G113), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT2), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT2), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G113), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(new_n338), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n341), .A2(new_n329), .A3(new_n332), .A4(new_n333), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n342), .A3(KEYINPUT67), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n342), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT67), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n343), .B(new_n346), .C1(new_n289), .C2(new_n290), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n328), .A2(G119), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n335), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n334), .B2(new_n349), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n351), .A2(new_n342), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n277), .A2(new_n352), .A3(new_n278), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G110), .B(G122), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n347), .A2(new_n353), .A3(new_n355), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(KEYINPUT6), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G125), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n262), .A2(new_n360), .A3(new_n251), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n285), .B1(new_n243), .B2(new_n261), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n247), .A2(new_n283), .A3(new_n248), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT82), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n262), .A2(new_n360), .A3(new_n251), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n366), .B(new_n367), .C1(new_n286), .C2(new_n360), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT83), .B(G224), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n189), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n365), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n371), .B1(new_n365), .B2(new_n368), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n354), .A2(new_n375), .A3(new_n356), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n359), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(KEYINPUT86), .B(new_n367), .C1(new_n286), .C2(new_n360), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT86), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n262), .A2(new_n251), .A3(new_n379), .A4(new_n360), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n370), .A2(KEYINPUT7), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT87), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OR3_X1    g199(.A1(new_n361), .A2(new_n364), .A3(new_n381), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n378), .A2(new_n382), .A3(KEYINPUT87), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(new_n358), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n389), .B1(new_n352), .B2(new_n258), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n351), .A2(KEYINPUT84), .A3(new_n342), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n351), .A2(new_n342), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n234), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n390), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(KEYINPUT85), .A3(new_n391), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n355), .B(KEYINPUT8), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n312), .B1(new_n388), .B2(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n325), .B(new_n327), .C1(new_n377), .C2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n359), .A2(new_n374), .A3(new_n376), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n378), .A2(new_n382), .A3(KEYINPUT87), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT87), .B1(new_n378), .B2(new_n382), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n394), .A2(new_n391), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n396), .B(new_n397), .C1(new_n407), .C2(new_n390), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n406), .A2(new_n408), .A3(new_n358), .A4(new_n386), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n403), .A2(new_n312), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n325), .B1(new_n410), .B2(new_n327), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n403), .A2(new_n409), .A3(new_n312), .A4(new_n326), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n402), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G214), .B1(G237), .B2(G902), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT9), .B(G234), .ZN(new_n417));
  INV_X1    g231(.A(G217), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n417), .A2(new_n418), .A3(G953), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n240), .A2(new_n242), .A3(G128), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n249), .A2(G143), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G134), .B1(new_n420), .B2(new_n421), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT94), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n421), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(G128), .A3(new_n237), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT94), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .A4(G134), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n420), .A2(new_n215), .A3(new_n422), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G122), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G116), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n328), .A2(G122), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n231), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n222), .A2(new_n224), .B1(new_n435), .B2(new_n436), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT92), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n253), .A2(new_n435), .A3(new_n436), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n231), .A2(new_n437), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT92), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n433), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n431), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT95), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n431), .A2(new_n445), .A3(KEYINPUT95), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n436), .A2(KEYINPUT14), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n435), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n436), .A2(KEYINPUT14), .ZN(new_n453));
  OAI21_X1  g267(.A(G107), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT96), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n441), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n437), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT96), .B1(new_n457), .B2(new_n253), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n454), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n215), .B1(new_n420), .B2(new_n422), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n433), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT97), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n441), .B(new_n455), .ZN(new_n463));
  INV_X1    g277(.A(new_n460), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n432), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT97), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n463), .A2(new_n465), .A3(new_n466), .A4(new_n454), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n419), .B1(new_n450), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n431), .A2(KEYINPUT95), .A3(new_n445), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT95), .B1(new_n431), .B2(new_n445), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n468), .B(new_n419), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n312), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT98), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT99), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(KEYINPUT15), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(KEYINPUT15), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n482));
  INV_X1    g296(.A(new_n419), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n472), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT98), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n312), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT18), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(KEYINPUT90), .ZN(new_n490));
  INV_X1    g304(.A(G237), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n189), .A3(G214), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(KEYINPUT89), .A3(new_n240), .A4(new_n242), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n491), .A2(new_n189), .A3(G143), .A4(G214), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT89), .B1(new_n237), .B2(new_n492), .ZN(new_n496));
  OAI211_X1 g310(.A(G131), .B(new_n490), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G140), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G125), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n360), .A2(G140), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT75), .ZN(new_n501));
  OR3_X1    g315(.A1(new_n360), .A2(KEYINPUT75), .A3(G140), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(G146), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n499), .A2(new_n500), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n260), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n240), .A2(new_n242), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n491), .A2(new_n189), .A3(G214), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n494), .A3(new_n493), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n489), .A2(new_n192), .A3(KEYINPUT90), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n497), .B(new_n506), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(G113), .B(G122), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n219), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT91), .ZN(new_n516));
  OAI21_X1  g330(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n510), .A2(new_n192), .A3(new_n494), .A4(new_n493), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT16), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT16), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n499), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G146), .ZN(new_n526));
  OAI211_X1 g340(.A(KEYINPUT17), .B(G131), .C1(new_n495), .C2(new_n496), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n260), .A3(new_n524), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n513), .B(new_n516), .C1(new_n521), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n520), .A2(new_n528), .A3(new_n526), .A4(new_n527), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n515), .B1(new_n532), .B2(new_n513), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n312), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G475), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n189), .A2(G952), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(G234), .B2(G237), .ZN(new_n537));
  INV_X1    g351(.A(G898), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n189), .B1(KEYINPUT21), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(KEYINPUT21), .B2(new_n538), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n312), .B1(G234), .B2(G237), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT20), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n504), .A2(KEYINPUT19), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n501), .A2(new_n502), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n546), .B1(new_n547), .B2(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n526), .B1(new_n548), .B2(G146), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n517), .A2(new_n519), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n513), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n515), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n530), .ZN(new_n554));
  NOR2_X1   g368(.A1(G475), .A2(G902), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n545), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n555), .ZN(new_n557));
  AOI211_X1 g371(.A(KEYINPUT20), .B(new_n557), .C1(new_n553), .C2(new_n530), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n535), .B(new_n544), .C1(new_n556), .C2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n474), .A2(new_n481), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n488), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n414), .A2(new_n416), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G221), .ZN(new_n564));
  INV_X1    g378(.A(new_n417), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n564), .B1(new_n565), .B2(new_n312), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n324), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT22), .B(G137), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n569), .B(new_n570), .Z(new_n571));
  NAND2_X1  g385(.A1(new_n526), .A2(new_n528), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n331), .A2(G128), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT73), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n249), .A2(G119), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT73), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n331), .A2(G128), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n574), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT24), .B(G110), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT74), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT23), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n573), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n575), .B1(new_n582), .B2(new_n583), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n578), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n581), .B1(G110), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n572), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n579), .A2(new_n580), .ZN(new_n591));
  INV_X1    g405(.A(G110), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n586), .A2(new_n592), .A3(new_n578), .A4(new_n587), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n591), .A2(new_n593), .B1(new_n260), .B2(new_n504), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n526), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(KEYINPUT76), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n572), .A2(new_n589), .B1(new_n594), .B2(new_n526), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT76), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n571), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n571), .B1(new_n598), .B2(new_n599), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n312), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT25), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n596), .A2(KEYINPUT76), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n598), .A2(new_n599), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n602), .B1(new_n609), .B2(new_n571), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(KEYINPUT25), .A3(new_n312), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n418), .B1(G234), .B2(new_n312), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(G902), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n612), .A2(new_n613), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n286), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n293), .A2(new_n294), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n197), .A2(G137), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n215), .B2(G137), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G131), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n217), .A2(new_n263), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT69), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n202), .A2(new_n216), .B1(G131), .B2(new_n620), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT69), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n263), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n618), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n346), .A2(new_n343), .ZN(new_n629));
  AND4_X1   g443(.A1(new_n625), .A2(new_n217), .A3(new_n263), .A4(new_n621), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n625), .B1(new_n624), .B2(new_n263), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n211), .A2(new_n286), .A3(new_n218), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(KEYINPUT30), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n622), .B1(new_n271), .B2(new_n617), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT30), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n629), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n628), .A2(new_n629), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n491), .A2(new_n189), .A3(G210), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT27), .Z(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT26), .B(G101), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT70), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n633), .A2(new_n623), .A3(new_n626), .A4(new_n629), .ZN(new_n645));
  INV_X1    g459(.A(new_n629), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n635), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT28), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n629), .A2(new_n622), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT28), .B1(new_n633), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n642), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT29), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n634), .A2(new_n637), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n645), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT70), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n642), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n644), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT71), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n633), .A2(new_n623), .A3(new_n626), .A4(new_n629), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT28), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT29), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n651), .A2(new_n663), .A3(new_n642), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT72), .B1(new_n665), .B2(new_n312), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT72), .ZN(new_n667));
  AOI211_X1 g481(.A(new_n667), .B(G902), .C1(new_n662), .C2(new_n664), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT71), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n644), .A2(new_n653), .A3(new_n657), .A4(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n659), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G472), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n623), .A2(KEYINPUT30), .A3(new_n626), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n618), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n213), .A2(new_n217), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n676), .A2(new_n286), .B1(new_n263), .B2(new_n624), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n646), .B1(new_n677), .B2(KEYINPUT30), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n645), .B(new_n643), .C1(new_n675), .C2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT31), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n654), .A2(KEYINPUT31), .A3(new_n645), .A4(new_n643), .ZN(new_n682));
  INV_X1    g496(.A(new_n651), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n649), .A2(new_n683), .ZN(new_n684));
  AOI22_X1  g498(.A1(new_n681), .A2(new_n682), .B1(new_n684), .B2(new_n642), .ZN(new_n685));
  NOR2_X1   g499(.A1(G472), .A2(G902), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT32), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n681), .A2(new_n682), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n684), .A2(new_n642), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT32), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n692), .A3(new_n686), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n616), .B1(new_n673), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n568), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G101), .ZN(G3));
  AND2_X1   g511(.A1(new_n324), .A2(new_n567), .ZN(new_n698));
  AOI21_X1  g512(.A(G902), .B1(new_n689), .B2(new_n690), .ZN(new_n699));
  INV_X1    g513(.A(G472), .ZN(new_n700));
  OAI22_X1  g514(.A1(new_n699), .A2(new_n700), .B1(new_n685), .B2(new_n687), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n616), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n703), .B(KEYINPUT100), .Z(new_n704));
  OAI21_X1  g518(.A(KEYINPUT33), .B1(new_n419), .B2(KEYINPUT101), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n485), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n705), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n484), .A2(new_n472), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n476), .A2(G902), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n475), .A2(new_n476), .A3(new_n487), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n706), .A2(KEYINPUT102), .A3(new_n708), .A4(new_n709), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n535), .B1(new_n556), .B2(new_n558), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n410), .A2(new_n327), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n416), .B1(new_n718), .B2(new_n412), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n544), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n704), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT34), .B(G104), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G6));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n488), .A2(new_n561), .ZN(new_n726));
  INV_X1    g540(.A(new_n716), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n725), .B1(new_n728), .B2(new_n720), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n716), .B1(new_n488), .B2(new_n561), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(KEYINPUT103), .A3(new_n544), .A4(new_n719), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n704), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT35), .B(G107), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G9));
  INV_X1    g549(.A(new_n571), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(KEYINPUT36), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n596), .B(new_n737), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n612), .A2(new_n613), .B1(new_n614), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT104), .B1(new_n701), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n739), .ZN(new_n741));
  OAI21_X1  g555(.A(G472), .B1(new_n685), .B2(G902), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n691), .A2(new_n686), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n741), .A2(new_n742), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n568), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g561(.A(KEYINPUT37), .B(G110), .Z(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G12));
  AOI22_X1  g563(.A1(new_n672), .A2(G472), .B1(new_n688), .B2(new_n693), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n741), .A2(new_n719), .ZN(new_n751));
  INV_X1    g565(.A(new_n542), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n189), .A2(G900), .ZN(new_n753));
  OR3_X1    g567(.A1(new_n752), .A2(KEYINPUT105), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n537), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT105), .B1(new_n752), .B2(new_n753), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n730), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n750), .A2(new_n751), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n698), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G128), .ZN(G30));
  XNOR2_X1  g575(.A(new_n757), .B(KEYINPUT39), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n324), .A2(new_n567), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT40), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n638), .A2(new_n642), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n660), .A2(new_n661), .A3(new_n643), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n766), .A2(G902), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n700), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n769), .B1(new_n688), .B2(new_n693), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n739), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n414), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n726), .A2(new_n716), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n772), .A2(new_n774), .A3(new_n416), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n763), .A2(new_n764), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n765), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n508), .ZN(G45));
  NAND3_X1  g593(.A1(new_n715), .A2(new_n716), .A3(new_n757), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n750), .A2(new_n751), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n698), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT107), .B(G146), .Z(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G48));
  OAI21_X1  g598(.A(new_n312), .B1(new_n321), .B2(new_n322), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(G469), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n323), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n566), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n695), .A2(new_n721), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(KEYINPUT41), .B(G113), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G15));
  NAND3_X1  g605(.A1(new_n695), .A2(new_n732), .A3(new_n788), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G116), .ZN(G18));
  AOI21_X1  g607(.A(new_n739), .B1(new_n673), .B2(new_n694), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n788), .A2(new_n719), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n562), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT108), .B(G119), .Z(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(G21));
  INV_X1    g613(.A(new_n742), .ZN(new_n800));
  INV_X1    g614(.A(new_n662), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n642), .B1(new_n801), .B2(new_n651), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(new_n689), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n687), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n800), .A2(new_n804), .A3(new_n616), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n726), .A2(new_n716), .A3(new_n719), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n544), .A3(new_n806), .A4(new_n788), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G122), .ZN(G24));
  OAI211_X1 g622(.A(new_n741), .B(new_n742), .C1(new_n687), .C2(new_n803), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n809), .A2(new_n780), .A3(new_n795), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(new_n360), .ZN(G27));
  NOR2_X1   g625(.A1(new_n310), .A2(new_n312), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n323), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n317), .A2(G469), .A3(new_n297), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n566), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n402), .A2(new_n411), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n413), .A2(new_n416), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n615), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n673), .B2(new_n694), .ZN(new_n820));
  INV_X1    g634(.A(new_n780), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT42), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT42), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n750), .A2(new_n819), .A3(new_n823), .A4(new_n780), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G131), .ZN(G33));
  AND3_X1   g640(.A1(new_n730), .A2(KEYINPUT109), .A3(new_n757), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT109), .B1(new_n730), .B2(new_n757), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n820), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G134), .ZN(G36));
  NAND2_X1  g645(.A1(new_n715), .A2(new_n727), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT43), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n739), .B1(new_n742), .B2(new_n744), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n836), .A2(KEYINPUT44), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n762), .A2(new_n567), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT45), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n313), .B2(new_n318), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(G469), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT110), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n843), .A3(G469), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n317), .A2(KEYINPUT45), .A3(new_n297), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT46), .B1(new_n846), .B2(new_n813), .ZN(new_n847));
  INV_X1    g661(.A(new_n323), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(KEYINPUT46), .A3(new_n813), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n838), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n834), .A2(KEYINPUT44), .A3(new_n835), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n402), .A2(new_n411), .A3(new_n413), .A4(new_n416), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n852), .A2(KEYINPUT111), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT111), .B1(new_n852), .B2(new_n853), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n837), .B(new_n851), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(KEYINPUT112), .B(G137), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n856), .B(new_n857), .ZN(G39));
  NAND3_X1  g672(.A1(new_n821), .A2(new_n616), .A3(new_n853), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n673), .A2(new_n694), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT47), .ZN(new_n863));
  INV_X1    g677(.A(new_n850), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n864), .A2(new_n847), .A3(new_n848), .ZN(new_n865));
  OAI211_X1 g679(.A(KEYINPUT113), .B(new_n863), .C1(new_n865), .C2(new_n566), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n849), .A2(new_n850), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT113), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n566), .B1(new_n868), .B2(KEYINPUT47), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n863), .A2(KEYINPUT113), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n862), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(new_n498), .ZN(G42));
  NAND3_X1  g687(.A1(new_n786), .A2(new_n566), .A3(new_n323), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n866), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n834), .A2(new_n537), .A3(new_n805), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n817), .A2(new_n818), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n788), .A2(new_n817), .A3(new_n818), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n834), .A2(new_n537), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT116), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n800), .A2(new_n804), .A3(new_n739), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT50), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n774), .A2(new_n416), .A3(new_n788), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n876), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n876), .B2(new_n886), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n880), .A2(new_n615), .A3(new_n770), .A4(new_n537), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT117), .Z(new_n891));
  INV_X1    g705(.A(new_n715), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n727), .A3(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n884), .A2(new_n889), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT51), .B1(new_n879), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n876), .A2(new_n795), .ZN(new_n896));
  INV_X1    g710(.A(new_n717), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n536), .B(new_n896), .C1(new_n891), .C2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT48), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n882), .A2(new_n899), .A3(new_n695), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n882), .B2(new_n695), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n879), .A2(new_n894), .A3(KEYINPUT51), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n908), .A2(new_n780), .ZN(new_n909));
  AOI22_X1  g723(.A1(new_n820), .A2(new_n829), .B1(new_n883), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT115), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n488), .A2(new_n561), .A3(new_n727), .A4(new_n757), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n877), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n912), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n853), .A2(new_n914), .A3(KEYINPUT115), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n698), .A2(new_n916), .A3(new_n794), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n910), .B(new_n917), .C1(new_n822), .C2(new_n824), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n568), .B1(new_n746), .B2(new_n695), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT114), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n717), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n715), .A2(KEYINPUT114), .A3(new_n716), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n728), .A3(new_n922), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n414), .A2(new_n416), .A3(new_n543), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n698), .A2(new_n923), .A3(new_n702), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n789), .A2(new_n792), .A3(new_n797), .A4(new_n807), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n918), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT52), .ZN(new_n929));
  INV_X1    g743(.A(new_n795), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n883), .A2(new_n821), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n751), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n860), .A2(new_n730), .A3(new_n932), .A4(new_n757), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n324), .A2(new_n567), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n815), .A2(new_n323), .A3(new_n813), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n936), .A2(new_n567), .A3(new_n757), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n771), .A2(new_n739), .A3(new_n806), .A4(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n860), .A2(new_n932), .A3(new_n821), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(new_n934), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n929), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n810), .B1(new_n759), .B2(new_n698), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n937), .A2(new_n726), .A3(new_n716), .A4(new_n719), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n943), .A2(new_n770), .A3(new_n741), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n781), .B2(new_n698), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n942), .A2(new_n945), .A3(KEYINPUT52), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n928), .A2(new_n947), .A3(KEYINPUT53), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT53), .B1(new_n928), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n907), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT53), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n942), .A2(new_n945), .A3(KEYINPUT52), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT52), .B1(new_n942), .B2(new_n945), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n919), .A2(new_n925), .ZN(new_n955));
  AND4_X1   g769(.A1(new_n789), .A2(new_n792), .A3(new_n797), .A4(new_n807), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n910), .A2(new_n917), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n955), .A2(new_n956), .A3(new_n825), .A4(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n951), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n928), .A2(new_n947), .A3(KEYINPUT53), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(KEYINPUT54), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n950), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n879), .A2(new_n894), .A3(KEYINPUT118), .A4(KEYINPUT51), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n903), .A2(new_n906), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(G952), .A2(G953), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT119), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n787), .B(KEYINPUT49), .ZN(new_n968));
  NOR4_X1   g782(.A1(new_n968), .A2(new_n616), .A3(new_n566), .A4(new_n416), .ZN(new_n969));
  INV_X1    g783(.A(new_n832), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n969), .A2(new_n770), .A3(new_n774), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(G75));
  NAND2_X1  g786(.A1(new_n959), .A2(new_n960), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(G210), .A3(G902), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT56), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n359), .A2(new_n376), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(new_n374), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n977), .A2(new_n377), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT55), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n974), .A2(new_n975), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n979), .B1(new_n974), .B2(new_n975), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n189), .A2(G952), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(G51));
  XOR2_X1   g797(.A(new_n812), .B(KEYINPUT57), .Z(new_n984));
  OAI22_X1  g798(.A1(new_n962), .A2(new_n984), .B1(new_n322), .B2(new_n321), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n846), .B(KEYINPUT120), .Z(new_n986));
  NAND3_X1  g800(.A1(new_n973), .A2(G902), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n982), .B1(new_n985), .B2(new_n987), .ZN(G54));
  NAND4_X1  g802(.A1(new_n973), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n989));
  INV_X1    g803(.A(new_n554), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n991), .A2(new_n992), .A3(new_n982), .ZN(G60));
  NAND2_X1  g807(.A1(G478), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT59), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n950), .A2(new_n961), .A3(new_n995), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n706), .A2(new_n708), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n982), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n950), .A2(new_n961), .A3(new_n997), .A4(new_n995), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(KEYINPUT121), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n1002), .A2(KEYINPUT121), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(G63));
  NAND2_X1  g819(.A1(G217), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT60), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n738), .B(new_n1008), .C1(new_n948), .C2(new_n949), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1007), .B1(new_n959), .B2(new_n960), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n1009), .B(new_n1000), .C1(new_n1010), .C2(new_n610), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT122), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n1011), .A2(new_n1012), .A3(KEYINPUT61), .ZN(new_n1013));
  AOI21_X1  g827(.A(KEYINPUT61), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1013), .A2(new_n1014), .ZN(G66));
  OAI21_X1  g829(.A(new_n540), .B1(new_n189), .B2(new_n369), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT123), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n955), .A2(new_n956), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1017), .B1(new_n1018), .B2(new_n189), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n976), .B1(new_n538), .B2(G953), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(G69));
  OAI21_X1  g835(.A(new_n634), .B1(KEYINPUT30), .B2(new_n677), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(new_n548), .Z(new_n1023));
  AND4_X1   g837(.A1(new_n782), .A2(new_n825), .A3(new_n830), .A4(new_n942), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n851), .A2(new_n695), .A3(new_n806), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1024), .A2(new_n856), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n189), .B1(new_n1026), .B2(new_n872), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1023), .B1(new_n1027), .B2(new_n753), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1029), .B(KEYINPUT126), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n765), .A2(new_n776), .A3(new_n777), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n942), .A2(new_n782), .ZN(new_n1033));
  OAI21_X1  g847(.A(KEYINPUT62), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT62), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n778), .A2(new_n1035), .A3(new_n782), .A4(new_n942), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n763), .A2(new_n695), .A3(new_n853), .A4(new_n923), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1037), .B(KEYINPUT124), .ZN(new_n1038));
  NAND4_X1  g852(.A1(new_n1034), .A2(new_n856), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1039), .A2(new_n872), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1023), .B1(new_n1040), .B2(G953), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(KEYINPUT125), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT125), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n1043), .B(new_n1023), .C1(new_n1040), .C2(G953), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1031), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1041), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1029), .B1(new_n1046), .B2(new_n1028), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1045), .A2(new_n1047), .ZN(G72));
  NOR3_X1   g862(.A1(new_n1026), .A2(new_n872), .A3(new_n1018), .ZN(new_n1049));
  NAND2_X1  g863(.A1(G472), .A2(G902), .ZN(new_n1050));
  XOR2_X1   g864(.A(new_n1050), .B(KEYINPUT63), .Z(new_n1051));
  INV_X1    g865(.A(new_n1051), .ZN(new_n1052));
  OAI211_X1 g866(.A(new_n642), .B(new_n638), .C1(new_n1049), .C2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n644), .A2(new_n679), .A3(new_n657), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1054), .A2(new_n1051), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1055), .B(KEYINPUT127), .Z(new_n1056));
  AOI21_X1  g870(.A(new_n982), .B1(new_n973), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1040), .ZN(new_n1059));
  OAI21_X1  g873(.A(new_n1051), .B1(new_n1059), .B2(new_n1018), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n1058), .B1(new_n766), .B2(new_n1060), .ZN(G57));
endmodule


